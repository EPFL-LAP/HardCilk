module ram_2x17 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [16:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [16:0] W0_data;
	reg [16:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 17'bxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_AddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_prot,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_prot
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [13:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_prot;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [13:0] io_deq_bits_addr;
	output wire [2:0] io_deq_bits_prot;
	wire [16:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x17 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_prot, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[13:0];
	assign io_deq_bits_prot = _ram_ext_R0_data[16:14];
endmodule
module ram_2x66 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [65:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [65:0] W0_data;
	reg [65:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 66'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	wire [65:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x66 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_resp, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[63:0];
	assign io_deq_bits_resp = _ram_ext_R0_data[65:64];
endmodule
module ram_2x72 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [71:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [71:0] W0_data;
	reg [71:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 72'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [7:0] io_enq_bits_strb;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [7:0] io_deq_bits_strb;
	wire [71:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x72 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_strb, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[63:0];
	assign io_deq_bits_strb = _ram_ext_R0_data[71:64];
endmodule
module ram_2x2 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [1:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [1:0] W0_data;
	reg [1:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 2'bxx);
endmodule
module Queue2_WriteResponseChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_resp;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x2 ram_resp_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_resp),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_resp)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module ram_8x3 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [2:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [2:0] R0_data;
	input [2:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [2:0] W0_data;
	reg [2:0] Memory [0:7];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 3'bxxx);
endmodule
module Queue8_UInt3 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits;
	wire io_enq_ready_0;
	wire [2:0] _ram_ext_R0_data;
	reg [2:0] enq_ptr_value;
	reg [2:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire io_deq_valid_0 = io_enq_valid | ~empty;
	wire do_deq = (~empty & io_deq_ready) & io_deq_valid_0;
	wire do_enq = (~(empty & io_deq_ready) & io_enq_ready_0) & io_enq_valid;
	assign io_enq_ready_0 = io_deq_ready | ~(ptr_match & maybe_full);
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 3'h0;
			deq_ptr_value <= 3'h0;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 3'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 3'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_8x3 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = io_enq_ready_0;
	assign io_deq_valid = io_deq_valid_0;
	assign io_deq_bits = (empty ? io_enq_bits : _ram_ext_R0_data);
endmodule
module elasticDemux (
	io_source_ready,
	io_source_valid,
	io_source_bits_addr,
	io_source_bits_prot,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_addr,
	io_sinks_0_bits_prot,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_addr,
	io_sinks_1_bits_prot,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_2_bits_addr,
	io_sinks_2_bits_prot,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_3_bits_addr,
	io_sinks_3_bits_prot,
	io_sinks_4_ready,
	io_sinks_4_valid,
	io_sinks_4_bits_addr,
	io_sinks_4_bits_prot,
	io_sinks_5_ready,
	io_sinks_5_valid,
	io_sinks_5_bits_addr,
	io_sinks_5_bits_prot,
	io_sinks_6_ready,
	io_sinks_6_valid,
	io_sinks_6_bits_addr,
	io_sinks_6_bits_prot,
	io_sinks_7_ready,
	io_sinks_7_valid,
	io_sinks_7_bits_addr,
	io_sinks_7_bits_prot,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [13:0] io_source_bits_addr;
	input [2:0] io_source_bits_prot;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [13:0] io_sinks_0_bits_addr;
	output wire [2:0] io_sinks_0_bits_prot;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [13:0] io_sinks_1_bits_addr;
	output wire [2:0] io_sinks_1_bits_prot;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	output wire [13:0] io_sinks_2_bits_addr;
	output wire [2:0] io_sinks_2_bits_prot;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire [13:0] io_sinks_3_bits_addr;
	output wire [2:0] io_sinks_3_bits_prot;
	input io_sinks_4_ready;
	output wire io_sinks_4_valid;
	output wire [13:0] io_sinks_4_bits_addr;
	output wire [2:0] io_sinks_4_bits_prot;
	input io_sinks_5_ready;
	output wire io_sinks_5_valid;
	output wire [13:0] io_sinks_5_bits_addr;
	output wire [2:0] io_sinks_5_bits_prot;
	input io_sinks_6_ready;
	output wire io_sinks_6_valid;
	output wire [13:0] io_sinks_6_bits_addr;
	output wire [2:0] io_sinks_6_bits_prot;
	input io_sinks_7_ready;
	output wire io_sinks_7_valid;
	output wire [13:0] io_sinks_7_bits_addr;
	output wire [2:0] io_sinks_7_bits_prot;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [7:0] _GEN = {io_sinks_7_ready, io_sinks_6_ready, io_sinks_5_ready, io_sinks_4_ready, io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 3'h0);
	assign io_sinks_0_bits_addr = io_source_bits_addr;
	assign io_sinks_0_bits_prot = io_source_bits_prot;
	assign io_sinks_1_valid = valid & (io_select_bits == 3'h1);
	assign io_sinks_1_bits_addr = io_source_bits_addr;
	assign io_sinks_1_bits_prot = io_source_bits_prot;
	assign io_sinks_2_valid = valid & (io_select_bits == 3'h2);
	assign io_sinks_2_bits_addr = io_source_bits_addr;
	assign io_sinks_2_bits_prot = io_source_bits_prot;
	assign io_sinks_3_valid = valid & (io_select_bits == 3'h3);
	assign io_sinks_3_bits_addr = io_source_bits_addr;
	assign io_sinks_3_bits_prot = io_source_bits_prot;
	assign io_sinks_4_valid = valid & (io_select_bits == 3'h4);
	assign io_sinks_4_bits_addr = io_source_bits_addr;
	assign io_sinks_4_bits_prot = io_source_bits_prot;
	assign io_sinks_5_valid = valid & (io_select_bits == 3'h5);
	assign io_sinks_5_bits_addr = io_source_bits_addr;
	assign io_sinks_5_bits_prot = io_source_bits_prot;
	assign io_sinks_6_valid = valid & (io_select_bits == 3'h6);
	assign io_sinks_6_bits_addr = io_source_bits_addr;
	assign io_sinks_6_bits_prot = io_source_bits_prot;
	assign io_sinks_7_valid = valid & (&io_select_bits);
	assign io_sinks_7_bits_addr = io_source_bits_addr;
	assign io_sinks_7_bits_prot = io_source_bits_prot;
	assign io_select_ready = fire;
endmodule
module elasticMux (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_data,
	io_sources_0_bits_resp,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_data,
	io_sources_1_bits_resp,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_data,
	io_sources_2_bits_resp,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_data,
	io_sources_3_bits_resp,
	io_sources_4_ready,
	io_sources_4_valid,
	io_sources_4_bits_data,
	io_sources_4_bits_resp,
	io_sources_5_ready,
	io_sources_5_valid,
	io_sources_5_bits_data,
	io_sources_5_bits_resp,
	io_sources_6_ready,
	io_sources_6_valid,
	io_sources_6_bits_data,
	io_sources_6_bits_resp,
	io_sources_7_ready,
	io_sources_7_valid,
	io_sources_7_bits_data,
	io_sources_7_bits_resp,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_data,
	io_sink_bits_resp,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [63:0] io_sources_0_bits_data;
	input [1:0] io_sources_0_bits_resp;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [63:0] io_sources_1_bits_data;
	input [1:0] io_sources_1_bits_resp;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [63:0] io_sources_2_bits_data;
	input [1:0] io_sources_2_bits_resp;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [63:0] io_sources_3_bits_data;
	input [1:0] io_sources_3_bits_resp;
	output wire io_sources_4_ready;
	input io_sources_4_valid;
	input [63:0] io_sources_4_bits_data;
	input [1:0] io_sources_4_bits_resp;
	output wire io_sources_5_ready;
	input io_sources_5_valid;
	input [63:0] io_sources_5_bits_data;
	input [1:0] io_sources_5_bits_resp;
	output wire io_sources_6_ready;
	input io_sources_6_valid;
	input [63:0] io_sources_6_bits_data;
	input [1:0] io_sources_6_bits_resp;
	output wire io_sources_7_ready;
	input io_sources_7_valid;
	input [63:0] io_sources_7_bits_data;
	input [1:0] io_sources_7_bits_resp;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [63:0] io_sink_bits_data;
	output wire [1:0] io_sink_bits_resp;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire [7:0] _GEN = {io_sources_7_valid, io_sources_6_valid, io_sources_5_valid, io_sources_4_valid, io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [511:0] _GEN_0 = {io_sources_7_bits_data, io_sources_6_bits_data, io_sources_5_bits_data, io_sources_4_bits_data, io_sources_3_bits_data, io_sources_2_bits_data, io_sources_1_bits_data, io_sources_0_bits_data};
	wire [15:0] _GEN_1 = {io_sources_7_bits_resp, io_sources_6_bits_resp, io_sources_5_bits_resp, io_sources_4_bits_resp, io_sources_3_bits_resp, io_sources_2_bits_resp, io_sources_1_bits_resp, io_sources_0_bits_resp};
	wire valid = io_select_valid & _GEN[io_select_bits];
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & (io_select_bits == 3'h0);
	assign io_sources_1_ready = fire & (io_select_bits == 3'h1);
	assign io_sources_2_ready = fire & (io_select_bits == 3'h2);
	assign io_sources_3_ready = fire & (io_select_bits == 3'h3);
	assign io_sources_4_ready = fire & (io_select_bits == 3'h4);
	assign io_sources_5_ready = fire & (io_select_bits == 3'h5);
	assign io_sources_6_ready = fire & (io_select_bits == 3'h6);
	assign io_sources_7_ready = fire & (&io_select_bits);
	assign io_sink_valid = valid;
	assign io_sink_bits_data = _GEN_0[io_select_bits * 64+:64];
	assign io_sink_bits_resp = _GEN_1[io_select_bits * 2+:2];
	assign io_select_ready = fire;
endmodule
module elasticDemux_2 (
	io_source_ready,
	io_source_valid,
	io_source_bits_data,
	io_source_bits_strb,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_data,
	io_sinks_0_bits_strb,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_data,
	io_sinks_1_bits_strb,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_2_bits_data,
	io_sinks_2_bits_strb,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_3_bits_data,
	io_sinks_3_bits_strb,
	io_sinks_4_ready,
	io_sinks_4_valid,
	io_sinks_4_bits_data,
	io_sinks_4_bits_strb,
	io_sinks_5_ready,
	io_sinks_5_valid,
	io_sinks_5_bits_data,
	io_sinks_5_bits_strb,
	io_sinks_6_ready,
	io_sinks_6_valid,
	io_sinks_6_bits_data,
	io_sinks_6_bits_strb,
	io_sinks_7_ready,
	io_sinks_7_valid,
	io_sinks_7_bits_data,
	io_sinks_7_bits_strb,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [63:0] io_source_bits_data;
	input [7:0] io_source_bits_strb;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [63:0] io_sinks_0_bits_data;
	output wire [7:0] io_sinks_0_bits_strb;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [63:0] io_sinks_1_bits_data;
	output wire [7:0] io_sinks_1_bits_strb;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	output wire [63:0] io_sinks_2_bits_data;
	output wire [7:0] io_sinks_2_bits_strb;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire [63:0] io_sinks_3_bits_data;
	output wire [7:0] io_sinks_3_bits_strb;
	input io_sinks_4_ready;
	output wire io_sinks_4_valid;
	output wire [63:0] io_sinks_4_bits_data;
	output wire [7:0] io_sinks_4_bits_strb;
	input io_sinks_5_ready;
	output wire io_sinks_5_valid;
	output wire [63:0] io_sinks_5_bits_data;
	output wire [7:0] io_sinks_5_bits_strb;
	input io_sinks_6_ready;
	output wire io_sinks_6_valid;
	output wire [63:0] io_sinks_6_bits_data;
	output wire [7:0] io_sinks_6_bits_strb;
	input io_sinks_7_ready;
	output wire io_sinks_7_valid;
	output wire [63:0] io_sinks_7_bits_data;
	output wire [7:0] io_sinks_7_bits_strb;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [7:0] _GEN = {io_sinks_7_ready, io_sinks_6_ready, io_sinks_5_ready, io_sinks_4_ready, io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 3'h0);
	assign io_sinks_0_bits_data = io_source_bits_data;
	assign io_sinks_0_bits_strb = io_source_bits_strb;
	assign io_sinks_1_valid = valid & (io_select_bits == 3'h1);
	assign io_sinks_1_bits_data = io_source_bits_data;
	assign io_sinks_1_bits_strb = io_source_bits_strb;
	assign io_sinks_2_valid = valid & (io_select_bits == 3'h2);
	assign io_sinks_2_bits_data = io_source_bits_data;
	assign io_sinks_2_bits_strb = io_source_bits_strb;
	assign io_sinks_3_valid = valid & (io_select_bits == 3'h3);
	assign io_sinks_3_bits_data = io_source_bits_data;
	assign io_sinks_3_bits_strb = io_source_bits_strb;
	assign io_sinks_4_valid = valid & (io_select_bits == 3'h4);
	assign io_sinks_4_bits_data = io_source_bits_data;
	assign io_sinks_4_bits_strb = io_source_bits_strb;
	assign io_sinks_5_valid = valid & (io_select_bits == 3'h5);
	assign io_sinks_5_bits_data = io_source_bits_data;
	assign io_sinks_5_bits_strb = io_source_bits_strb;
	assign io_sinks_6_valid = valid & (io_select_bits == 3'h6);
	assign io_sinks_6_bits_data = io_source_bits_data;
	assign io_sinks_6_bits_strb = io_source_bits_strb;
	assign io_sinks_7_valid = valid & (&io_select_bits);
	assign io_sinks_7_bits_data = io_source_bits_data;
	assign io_sinks_7_bits_strb = io_source_bits_strb;
	assign io_select_ready = fire;
endmodule
module elasticMux_1 (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_resp,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_resp,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_resp,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_resp,
	io_sources_4_ready,
	io_sources_4_valid,
	io_sources_4_bits_resp,
	io_sources_5_ready,
	io_sources_5_valid,
	io_sources_5_bits_resp,
	io_sources_6_ready,
	io_sources_6_valid,
	io_sources_6_bits_resp,
	io_sources_7_ready,
	io_sources_7_valid,
	io_sources_7_bits_resp,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_resp,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [1:0] io_sources_0_bits_resp;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [1:0] io_sources_1_bits_resp;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [1:0] io_sources_2_bits_resp;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [1:0] io_sources_3_bits_resp;
	output wire io_sources_4_ready;
	input io_sources_4_valid;
	input [1:0] io_sources_4_bits_resp;
	output wire io_sources_5_ready;
	input io_sources_5_valid;
	input [1:0] io_sources_5_bits_resp;
	output wire io_sources_6_ready;
	input io_sources_6_valid;
	input [1:0] io_sources_6_bits_resp;
	output wire io_sources_7_ready;
	input io_sources_7_valid;
	input [1:0] io_sources_7_bits_resp;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [1:0] io_sink_bits_resp;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire [7:0] _GEN = {io_sources_7_valid, io_sources_6_valid, io_sources_5_valid, io_sources_4_valid, io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [15:0] _GEN_0 = {io_sources_7_bits_resp, io_sources_6_bits_resp, io_sources_5_bits_resp, io_sources_4_bits_resp, io_sources_3_bits_resp, io_sources_2_bits_resp, io_sources_1_bits_resp, io_sources_0_bits_resp};
	wire valid = io_select_valid & _GEN[io_select_bits];
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & (io_select_bits == 3'h0);
	assign io_sources_1_ready = fire & (io_select_bits == 3'h1);
	assign io_sources_2_ready = fire & (io_select_bits == 3'h2);
	assign io_sources_3_ready = fire & (io_select_bits == 3'h3);
	assign io_sources_4_ready = fire & (io_select_bits == 3'h4);
	assign io_sources_5_ready = fire & (io_select_bits == 3'h5);
	assign io_sources_6_ready = fire & (io_select_bits == 3'h6);
	assign io_sources_7_ready = fire & (&io_select_bits);
	assign io_sink_valid = valid;
	assign io_sink_bits_resp = _GEN_0[io_select_bits * 2+:2];
	assign io_select_ready = fire;
endmodule
module axi4LiteDemux (
	clock,
	reset,
	s_axil_ar_ready,
	s_axil_ar_valid,
	s_axil_ar_bits_addr,
	s_axil_ar_bits_prot,
	s_axil_r_ready,
	s_axil_r_valid,
	s_axil_r_bits_data,
	s_axil_r_bits_resp,
	s_axil_aw_ready,
	s_axil_aw_valid,
	s_axil_aw_bits_addr,
	s_axil_aw_bits_prot,
	s_axil_w_ready,
	s_axil_w_valid,
	s_axil_w_bits_data,
	s_axil_w_bits_strb,
	s_axil_b_ready,
	s_axil_b_valid,
	s_axil_b_bits_resp,
	m_axil_0_ar_ready,
	m_axil_0_ar_valid,
	m_axil_0_ar_bits_addr,
	m_axil_0_ar_bits_prot,
	m_axil_0_r_ready,
	m_axil_0_r_valid,
	m_axil_0_r_bits_data,
	m_axil_0_r_bits_resp,
	m_axil_0_aw_ready,
	m_axil_0_aw_valid,
	m_axil_0_aw_bits_addr,
	m_axil_0_aw_bits_prot,
	m_axil_0_w_ready,
	m_axil_0_w_valid,
	m_axil_0_w_bits_data,
	m_axil_0_w_bits_strb,
	m_axil_0_b_ready,
	m_axil_0_b_valid,
	m_axil_0_b_bits_resp,
	m_axil_1_ar_ready,
	m_axil_1_ar_valid,
	m_axil_1_ar_bits_addr,
	m_axil_1_ar_bits_prot,
	m_axil_1_r_ready,
	m_axil_1_r_valid,
	m_axil_1_r_bits_data,
	m_axil_1_r_bits_resp,
	m_axil_1_aw_ready,
	m_axil_1_aw_valid,
	m_axil_1_aw_bits_addr,
	m_axil_1_aw_bits_prot,
	m_axil_1_w_ready,
	m_axil_1_w_valid,
	m_axil_1_w_bits_data,
	m_axil_1_w_bits_strb,
	m_axil_1_b_ready,
	m_axil_1_b_valid,
	m_axil_1_b_bits_resp,
	m_axil_2_ar_ready,
	m_axil_2_ar_valid,
	m_axil_2_ar_bits_addr,
	m_axil_2_ar_bits_prot,
	m_axil_2_r_ready,
	m_axil_2_r_valid,
	m_axil_2_r_bits_data,
	m_axil_2_r_bits_resp,
	m_axil_2_aw_ready,
	m_axil_2_aw_valid,
	m_axil_2_aw_bits_addr,
	m_axil_2_aw_bits_prot,
	m_axil_2_w_ready,
	m_axil_2_w_valid,
	m_axil_2_w_bits_data,
	m_axil_2_w_bits_strb,
	m_axil_2_b_ready,
	m_axil_2_b_valid,
	m_axil_2_b_bits_resp,
	m_axil_3_ar_ready,
	m_axil_3_ar_valid,
	m_axil_3_ar_bits_addr,
	m_axil_3_ar_bits_prot,
	m_axil_3_r_ready,
	m_axil_3_r_valid,
	m_axil_3_r_bits_data,
	m_axil_3_r_bits_resp,
	m_axil_3_aw_ready,
	m_axil_3_aw_valid,
	m_axil_3_aw_bits_addr,
	m_axil_3_aw_bits_prot,
	m_axil_3_w_ready,
	m_axil_3_w_valid,
	m_axil_3_w_bits_data,
	m_axil_3_w_bits_strb,
	m_axil_3_b_ready,
	m_axil_3_b_valid,
	m_axil_3_b_bits_resp,
	m_axil_4_ar_ready,
	m_axil_4_ar_valid,
	m_axil_4_ar_bits_addr,
	m_axil_4_ar_bits_prot,
	m_axil_4_r_ready,
	m_axil_4_r_valid,
	m_axil_4_r_bits_data,
	m_axil_4_r_bits_resp,
	m_axil_4_aw_ready,
	m_axil_4_aw_valid,
	m_axil_4_aw_bits_addr,
	m_axil_4_aw_bits_prot,
	m_axil_4_w_ready,
	m_axil_4_w_valid,
	m_axil_4_w_bits_data,
	m_axil_4_w_bits_strb,
	m_axil_4_b_ready,
	m_axil_4_b_valid,
	m_axil_4_b_bits_resp,
	m_axil_5_ar_ready,
	m_axil_5_ar_valid,
	m_axil_5_ar_bits_addr,
	m_axil_5_ar_bits_prot,
	m_axil_5_r_ready,
	m_axil_5_r_valid,
	m_axil_5_r_bits_data,
	m_axil_5_r_bits_resp,
	m_axil_5_aw_ready,
	m_axil_5_aw_valid,
	m_axil_5_aw_bits_addr,
	m_axil_5_aw_bits_prot,
	m_axil_5_w_ready,
	m_axil_5_w_valid,
	m_axil_5_w_bits_data,
	m_axil_5_w_bits_strb,
	m_axil_5_b_ready,
	m_axil_5_b_valid,
	m_axil_5_b_bits_resp,
	m_axil_6_ar_ready,
	m_axil_6_ar_valid,
	m_axil_6_ar_bits_addr,
	m_axil_6_ar_bits_prot,
	m_axil_6_r_ready,
	m_axil_6_r_valid,
	m_axil_6_r_bits_data,
	m_axil_6_r_bits_resp,
	m_axil_6_aw_ready,
	m_axil_6_aw_valid,
	m_axil_6_aw_bits_addr,
	m_axil_6_aw_bits_prot,
	m_axil_6_w_ready,
	m_axil_6_w_valid,
	m_axil_6_w_bits_data,
	m_axil_6_w_bits_strb,
	m_axil_6_b_ready,
	m_axil_6_b_valid,
	m_axil_6_b_bits_resp,
	m_axil_7_ar_ready,
	m_axil_7_ar_valid,
	m_axil_7_ar_bits_addr,
	m_axil_7_ar_bits_prot,
	m_axil_7_r_ready,
	m_axil_7_r_valid,
	m_axil_7_r_bits_data,
	m_axil_7_r_bits_resp,
	m_axil_7_aw_ready,
	m_axil_7_aw_valid,
	m_axil_7_aw_bits_addr,
	m_axil_7_aw_bits_prot,
	m_axil_7_w_ready,
	m_axil_7_w_valid,
	m_axil_7_w_bits_data,
	m_axil_7_w_bits_strb,
	m_axil_7_b_ready,
	m_axil_7_b_valid,
	m_axil_7_b_bits_resp
);
	input clock;
	input reset;
	output wire s_axil_ar_ready;
	input s_axil_ar_valid;
	input [13:0] s_axil_ar_bits_addr;
	input [2:0] s_axil_ar_bits_prot;
	input s_axil_r_ready;
	output wire s_axil_r_valid;
	output wire [63:0] s_axil_r_bits_data;
	output wire [1:0] s_axil_r_bits_resp;
	output wire s_axil_aw_ready;
	input s_axil_aw_valid;
	input [13:0] s_axil_aw_bits_addr;
	input [2:0] s_axil_aw_bits_prot;
	output wire s_axil_w_ready;
	input s_axil_w_valid;
	input [63:0] s_axil_w_bits_data;
	input [7:0] s_axil_w_bits_strb;
	input s_axil_b_ready;
	output wire s_axil_b_valid;
	output wire [1:0] s_axil_b_bits_resp;
	input m_axil_0_ar_ready;
	output wire m_axil_0_ar_valid;
	output wire [13:0] m_axil_0_ar_bits_addr;
	output wire [2:0] m_axil_0_ar_bits_prot;
	output wire m_axil_0_r_ready;
	input m_axil_0_r_valid;
	input [63:0] m_axil_0_r_bits_data;
	input [1:0] m_axil_0_r_bits_resp;
	input m_axil_0_aw_ready;
	output wire m_axil_0_aw_valid;
	output wire [13:0] m_axil_0_aw_bits_addr;
	output wire [2:0] m_axil_0_aw_bits_prot;
	input m_axil_0_w_ready;
	output wire m_axil_0_w_valid;
	output wire [63:0] m_axil_0_w_bits_data;
	output wire [7:0] m_axil_0_w_bits_strb;
	output wire m_axil_0_b_ready;
	input m_axil_0_b_valid;
	input [1:0] m_axil_0_b_bits_resp;
	input m_axil_1_ar_ready;
	output wire m_axil_1_ar_valid;
	output wire [13:0] m_axil_1_ar_bits_addr;
	output wire [2:0] m_axil_1_ar_bits_prot;
	output wire m_axil_1_r_ready;
	input m_axil_1_r_valid;
	input [63:0] m_axil_1_r_bits_data;
	input [1:0] m_axil_1_r_bits_resp;
	input m_axil_1_aw_ready;
	output wire m_axil_1_aw_valid;
	output wire [13:0] m_axil_1_aw_bits_addr;
	output wire [2:0] m_axil_1_aw_bits_prot;
	input m_axil_1_w_ready;
	output wire m_axil_1_w_valid;
	output wire [63:0] m_axil_1_w_bits_data;
	output wire [7:0] m_axil_1_w_bits_strb;
	output wire m_axil_1_b_ready;
	input m_axil_1_b_valid;
	input [1:0] m_axil_1_b_bits_resp;
	input m_axil_2_ar_ready;
	output wire m_axil_2_ar_valid;
	output wire [13:0] m_axil_2_ar_bits_addr;
	output wire [2:0] m_axil_2_ar_bits_prot;
	output wire m_axil_2_r_ready;
	input m_axil_2_r_valid;
	input [63:0] m_axil_2_r_bits_data;
	input [1:0] m_axil_2_r_bits_resp;
	input m_axil_2_aw_ready;
	output wire m_axil_2_aw_valid;
	output wire [13:0] m_axil_2_aw_bits_addr;
	output wire [2:0] m_axil_2_aw_bits_prot;
	input m_axil_2_w_ready;
	output wire m_axil_2_w_valid;
	output wire [63:0] m_axil_2_w_bits_data;
	output wire [7:0] m_axil_2_w_bits_strb;
	output wire m_axil_2_b_ready;
	input m_axil_2_b_valid;
	input [1:0] m_axil_2_b_bits_resp;
	input m_axil_3_ar_ready;
	output wire m_axil_3_ar_valid;
	output wire [13:0] m_axil_3_ar_bits_addr;
	output wire [2:0] m_axil_3_ar_bits_prot;
	output wire m_axil_3_r_ready;
	input m_axil_3_r_valid;
	input [63:0] m_axil_3_r_bits_data;
	input [1:0] m_axil_3_r_bits_resp;
	input m_axil_3_aw_ready;
	output wire m_axil_3_aw_valid;
	output wire [13:0] m_axil_3_aw_bits_addr;
	output wire [2:0] m_axil_3_aw_bits_prot;
	input m_axil_3_w_ready;
	output wire m_axil_3_w_valid;
	output wire [63:0] m_axil_3_w_bits_data;
	output wire [7:0] m_axil_3_w_bits_strb;
	output wire m_axil_3_b_ready;
	input m_axil_3_b_valid;
	input [1:0] m_axil_3_b_bits_resp;
	input m_axil_4_ar_ready;
	output wire m_axil_4_ar_valid;
	output wire [13:0] m_axil_4_ar_bits_addr;
	output wire [2:0] m_axil_4_ar_bits_prot;
	output wire m_axil_4_r_ready;
	input m_axil_4_r_valid;
	input [63:0] m_axil_4_r_bits_data;
	input [1:0] m_axil_4_r_bits_resp;
	input m_axil_4_aw_ready;
	output wire m_axil_4_aw_valid;
	output wire [13:0] m_axil_4_aw_bits_addr;
	output wire [2:0] m_axil_4_aw_bits_prot;
	input m_axil_4_w_ready;
	output wire m_axil_4_w_valid;
	output wire [63:0] m_axil_4_w_bits_data;
	output wire [7:0] m_axil_4_w_bits_strb;
	output wire m_axil_4_b_ready;
	input m_axil_4_b_valid;
	input [1:0] m_axil_4_b_bits_resp;
	input m_axil_5_ar_ready;
	output wire m_axil_5_ar_valid;
	output wire [13:0] m_axil_5_ar_bits_addr;
	output wire [2:0] m_axil_5_ar_bits_prot;
	output wire m_axil_5_r_ready;
	input m_axil_5_r_valid;
	input [63:0] m_axil_5_r_bits_data;
	input [1:0] m_axil_5_r_bits_resp;
	input m_axil_5_aw_ready;
	output wire m_axil_5_aw_valid;
	output wire [13:0] m_axil_5_aw_bits_addr;
	output wire [2:0] m_axil_5_aw_bits_prot;
	input m_axil_5_w_ready;
	output wire m_axil_5_w_valid;
	output wire [63:0] m_axil_5_w_bits_data;
	output wire [7:0] m_axil_5_w_bits_strb;
	output wire m_axil_5_b_ready;
	input m_axil_5_b_valid;
	input [1:0] m_axil_5_b_bits_resp;
	input m_axil_6_ar_ready;
	output wire m_axil_6_ar_valid;
	output wire [13:0] m_axil_6_ar_bits_addr;
	output wire [2:0] m_axil_6_ar_bits_prot;
	output wire m_axil_6_r_ready;
	input m_axil_6_r_valid;
	input [63:0] m_axil_6_r_bits_data;
	input [1:0] m_axil_6_r_bits_resp;
	input m_axil_6_aw_ready;
	output wire m_axil_6_aw_valid;
	output wire [13:0] m_axil_6_aw_bits_addr;
	output wire [2:0] m_axil_6_aw_bits_prot;
	input m_axil_6_w_ready;
	output wire m_axil_6_w_valid;
	output wire [63:0] m_axil_6_w_bits_data;
	output wire [7:0] m_axil_6_w_bits_strb;
	output wire m_axil_6_b_ready;
	input m_axil_6_b_valid;
	input [1:0] m_axil_6_b_bits_resp;
	input m_axil_7_ar_ready;
	output wire m_axil_7_ar_valid;
	output wire [13:0] m_axil_7_ar_bits_addr;
	output wire [2:0] m_axil_7_ar_bits_prot;
	output wire m_axil_7_r_ready;
	input m_axil_7_r_valid;
	input [63:0] m_axil_7_r_bits_data;
	input [1:0] m_axil_7_r_bits_resp;
	input m_axil_7_aw_ready;
	output wire m_axil_7_aw_valid;
	output wire [13:0] m_axil_7_aw_bits_addr;
	output wire [2:0] m_axil_7_aw_bits_prot;
	input m_axil_7_w_ready;
	output wire m_axil_7_w_valid;
	output wire [63:0] m_axil_7_w_bits_data;
	output wire [7:0] m_axil_7_w_bits_strb;
	output wire m_axil_7_b_ready;
	input m_axil_7_b_valid;
	input [1:0] m_axil_7_b_bits_resp;
	wire _write_mux_io_sink_valid;
	wire [1:0] _write_mux_io_sink_bits_resp;
	wire _write_mux_io_select_ready;
	wire _write_demux_1_io_source_ready;
	wire _write_demux_1_io_select_ready;
	wire _write_demux_io_source_ready;
	wire _write_demux_io_select_ready;
	wire _write_portQueueB_io_enq_ready;
	wire _write_portQueueB_io_deq_valid;
	wire [2:0] _write_portQueueB_io_deq_bits;
	wire _write_portQueueW_io_enq_ready;
	wire _write_portQueueW_io_deq_valid;
	wire [2:0] _write_portQueueW_io_deq_bits;
	wire _read_mux_io_sink_valid;
	wire [63:0] _read_mux_io_sink_bits_data;
	wire [1:0] _read_mux_io_sink_bits_resp;
	wire _read_mux_io_select_ready;
	wire _read_demux_io_source_ready;
	wire _read_demux_io_select_ready;
	wire _read_portQueue_io_enq_ready;
	wire _read_portQueue_io_deq_valid;
	wire [2:0] _read_portQueue_io_deq_bits;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [13:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [13:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	reg read_eagerFork_regs_0;
	reg read_eagerFork_regs_1;
	reg read_eagerFork_regs_2;
	wire read_eagerFork_arPort_ready_qual1_0 = _read_demux_io_source_ready | read_eagerFork_regs_0;
	wire read_eagerFork_arPort_ready_qual1_1 = _read_demux_io_select_ready | read_eagerFork_regs_1;
	wire read_eagerFork_arPort_ready_qual1_2 = _read_portQueue_io_enq_ready | read_eagerFork_regs_2;
	wire read_result_ready = (read_eagerFork_arPort_ready_qual1_0 & read_eagerFork_arPort_ready_qual1_1) & read_eagerFork_arPort_ready_qual1_2;
	reg write_eagerFork_regs_0;
	reg write_eagerFork_regs_1;
	reg write_eagerFork_regs_2;
	reg write_eagerFork_regs_3;
	wire write_eagerFork_awPort_ready_qual1_0 = _write_demux_io_source_ready | write_eagerFork_regs_0;
	wire write_eagerFork_awPort_ready_qual1_1 = _write_demux_io_select_ready | write_eagerFork_regs_1;
	wire write_eagerFork_awPort_ready_qual1_2 = _write_portQueueW_io_enq_ready | write_eagerFork_regs_2;
	wire write_eagerFork_awPort_ready_qual1_3 = _write_portQueueB_io_enq_ready | write_eagerFork_regs_3;
	wire write_result_ready = ((write_eagerFork_awPort_ready_qual1_0 & write_eagerFork_awPort_ready_qual1_1) & write_eagerFork_awPort_ready_qual1_2) & write_eagerFork_awPort_ready_qual1_3;
	always @(posedge clock)
		if (reset) begin
			read_eagerFork_regs_0 <= 1'h0;
			read_eagerFork_regs_1 <= 1'h0;
			read_eagerFork_regs_2 <= 1'h0;
			write_eagerFork_regs_0 <= 1'h0;
			write_eagerFork_regs_1 <= 1'h0;
			write_eagerFork_regs_2 <= 1'h0;
			write_eagerFork_regs_3 <= 1'h0;
		end
		else begin
			read_eagerFork_regs_0 <= (read_eagerFork_arPort_ready_qual1_0 & _s_axil__sourceBuffer_io_deq_valid) & ~read_result_ready;
			read_eagerFork_regs_1 <= (read_eagerFork_arPort_ready_qual1_1 & _s_axil__sourceBuffer_io_deq_valid) & ~read_result_ready;
			read_eagerFork_regs_2 <= (read_eagerFork_arPort_ready_qual1_2 & _s_axil__sourceBuffer_io_deq_valid) & ~read_result_ready;
			write_eagerFork_regs_0 <= (write_eagerFork_awPort_ready_qual1_0 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
			write_eagerFork_regs_1 <= (write_eagerFork_awPort_ready_qual1_1 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
			write_eagerFork_regs_2 <= (write_eagerFork_awPort_ready_qual1_2 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
			write_eagerFork_regs_3 <= (write_eagerFork_awPort_ready_qual1_3 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
		end
	Queue2_AddressChannel s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axil_ar_ready),
		.io_enq_valid(s_axil_ar_valid),
		.io_enq_bits_addr(s_axil_ar_bits_addr),
		.io_enq_bits_prot(s_axil_ar_bits_prot),
		.io_deq_ready(read_result_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_read_mux_io_sink_valid),
		.io_enq_bits_data(_read_mux_io_sink_bits_data),
		.io_enq_bits_resp(_read_mux_io_sink_bits_resp),
		.io_deq_ready(s_axil_r_ready),
		.io_deq_valid(s_axil_r_valid),
		.io_deq_bits_data(s_axil_r_bits_data),
		.io_deq_bits_resp(s_axil_r_bits_resp)
	);
	Queue2_AddressChannel s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axil_aw_ready),
		.io_enq_valid(s_axil_aw_valid),
		.io_enq_bits_addr(s_axil_aw_bits_addr),
		.io_enq_bits_prot(s_axil_aw_bits_prot),
		.io_deq_ready(write_result_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axil_w_ready),
		.io_enq_valid(s_axil_w_valid),
		.io_enq_bits_data(s_axil_w_bits_data),
		.io_enq_bits_strb(s_axil_w_bits_strb),
		.io_deq_ready(_write_demux_1_io_source_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_write_mux_io_sink_valid),
		.io_enq_bits_resp(_write_mux_io_sink_bits_resp),
		.io_deq_ready(s_axil_b_ready),
		.io_deq_valid(s_axil_b_valid),
		.io_deq_bits_resp(s_axil_b_bits_resp)
	);
	Queue8_UInt3 read_portQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_read_portQueue_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid & ~read_eagerFork_regs_2),
		.io_enq_bits(_s_axil__sourceBuffer_io_deq_bits_addr[8:6]),
		.io_deq_ready(_read_mux_io_select_ready),
		.io_deq_valid(_read_portQueue_io_deq_valid),
		.io_deq_bits(_read_portQueue_io_deq_bits)
	);
	elasticDemux read_demux(
		.io_source_ready(_read_demux_io_source_ready),
		.io_source_valid(_s_axil__sourceBuffer_io_deq_valid & ~read_eagerFork_regs_0),
		.io_source_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_source_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_sinks_0_ready(m_axil_0_ar_ready),
		.io_sinks_0_valid(m_axil_0_ar_valid),
		.io_sinks_0_bits_addr(m_axil_0_ar_bits_addr),
		.io_sinks_0_bits_prot(m_axil_0_ar_bits_prot),
		.io_sinks_1_ready(m_axil_1_ar_ready),
		.io_sinks_1_valid(m_axil_1_ar_valid),
		.io_sinks_1_bits_addr(m_axil_1_ar_bits_addr),
		.io_sinks_1_bits_prot(m_axil_1_ar_bits_prot),
		.io_sinks_2_ready(m_axil_2_ar_ready),
		.io_sinks_2_valid(m_axil_2_ar_valid),
		.io_sinks_2_bits_addr(m_axil_2_ar_bits_addr),
		.io_sinks_2_bits_prot(m_axil_2_ar_bits_prot),
		.io_sinks_3_ready(m_axil_3_ar_ready),
		.io_sinks_3_valid(m_axil_3_ar_valid),
		.io_sinks_3_bits_addr(m_axil_3_ar_bits_addr),
		.io_sinks_3_bits_prot(m_axil_3_ar_bits_prot),
		.io_sinks_4_ready(m_axil_4_ar_ready),
		.io_sinks_4_valid(m_axil_4_ar_valid),
		.io_sinks_4_bits_addr(m_axil_4_ar_bits_addr),
		.io_sinks_4_bits_prot(m_axil_4_ar_bits_prot),
		.io_sinks_5_ready(m_axil_5_ar_ready),
		.io_sinks_5_valid(m_axil_5_ar_valid),
		.io_sinks_5_bits_addr(m_axil_5_ar_bits_addr),
		.io_sinks_5_bits_prot(m_axil_5_ar_bits_prot),
		.io_sinks_6_ready(m_axil_6_ar_ready),
		.io_sinks_6_valid(m_axil_6_ar_valid),
		.io_sinks_6_bits_addr(m_axil_6_ar_bits_addr),
		.io_sinks_6_bits_prot(m_axil_6_ar_bits_prot),
		.io_sinks_7_ready(m_axil_7_ar_ready),
		.io_sinks_7_valid(m_axil_7_ar_valid),
		.io_sinks_7_bits_addr(m_axil_7_ar_bits_addr),
		.io_sinks_7_bits_prot(m_axil_7_ar_bits_prot),
		.io_select_ready(_read_demux_io_select_ready),
		.io_select_valid(_s_axil__sourceBuffer_io_deq_valid & ~read_eagerFork_regs_1),
		.io_select_bits(_s_axil__sourceBuffer_io_deq_bits_addr[8:6])
	);
	elasticMux read_mux(
		.io_sources_0_ready(m_axil_0_r_ready),
		.io_sources_0_valid(m_axil_0_r_valid),
		.io_sources_0_bits_data(m_axil_0_r_bits_data),
		.io_sources_0_bits_resp(m_axil_0_r_bits_resp),
		.io_sources_1_ready(m_axil_1_r_ready),
		.io_sources_1_valid(m_axil_1_r_valid),
		.io_sources_1_bits_data(m_axil_1_r_bits_data),
		.io_sources_1_bits_resp(m_axil_1_r_bits_resp),
		.io_sources_2_ready(m_axil_2_r_ready),
		.io_sources_2_valid(m_axil_2_r_valid),
		.io_sources_2_bits_data(m_axil_2_r_bits_data),
		.io_sources_2_bits_resp(m_axil_2_r_bits_resp),
		.io_sources_3_ready(m_axil_3_r_ready),
		.io_sources_3_valid(m_axil_3_r_valid),
		.io_sources_3_bits_data(m_axil_3_r_bits_data),
		.io_sources_3_bits_resp(m_axil_3_r_bits_resp),
		.io_sources_4_ready(m_axil_4_r_ready),
		.io_sources_4_valid(m_axil_4_r_valid),
		.io_sources_4_bits_data(m_axil_4_r_bits_data),
		.io_sources_4_bits_resp(m_axil_4_r_bits_resp),
		.io_sources_5_ready(m_axil_5_r_ready),
		.io_sources_5_valid(m_axil_5_r_valid),
		.io_sources_5_bits_data(m_axil_5_r_bits_data),
		.io_sources_5_bits_resp(m_axil_5_r_bits_resp),
		.io_sources_6_ready(m_axil_6_r_ready),
		.io_sources_6_valid(m_axil_6_r_valid),
		.io_sources_6_bits_data(m_axil_6_r_bits_data),
		.io_sources_6_bits_resp(m_axil_6_r_bits_resp),
		.io_sources_7_ready(m_axil_7_r_ready),
		.io_sources_7_valid(m_axil_7_r_valid),
		.io_sources_7_bits_data(m_axil_7_r_bits_data),
		.io_sources_7_bits_resp(m_axil_7_r_bits_resp),
		.io_sink_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_sink_valid(_read_mux_io_sink_valid),
		.io_sink_bits_data(_read_mux_io_sink_bits_data),
		.io_sink_bits_resp(_read_mux_io_sink_bits_resp),
		.io_select_ready(_read_mux_io_select_ready),
		.io_select_valid(_read_portQueue_io_deq_valid),
		.io_select_bits(_read_portQueue_io_deq_bits)
	);
	Queue8_UInt3 write_portQueueW(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueueW_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_2),
		.io_enq_bits(_s_axil__sourceBuffer_1_io_deq_bits_addr[8:6]),
		.io_deq_ready(_write_demux_1_io_select_ready),
		.io_deq_valid(_write_portQueueW_io_deq_valid),
		.io_deq_bits(_write_portQueueW_io_deq_bits)
	);
	Queue8_UInt3 write_portQueueB(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueueB_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_3),
		.io_enq_bits(_s_axil__sourceBuffer_1_io_deq_bits_addr[8:6]),
		.io_deq_ready(_write_mux_io_select_ready),
		.io_deq_valid(_write_portQueueB_io_deq_valid),
		.io_deq_bits(_write_portQueueB_io_deq_bits)
	);
	elasticDemux write_demux(
		.io_source_ready(_write_demux_io_source_ready),
		.io_source_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_0),
		.io_source_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_source_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_sinks_0_ready(m_axil_0_aw_ready),
		.io_sinks_0_valid(m_axil_0_aw_valid),
		.io_sinks_0_bits_addr(m_axil_0_aw_bits_addr),
		.io_sinks_0_bits_prot(m_axil_0_aw_bits_prot),
		.io_sinks_1_ready(m_axil_1_aw_ready),
		.io_sinks_1_valid(m_axil_1_aw_valid),
		.io_sinks_1_bits_addr(m_axil_1_aw_bits_addr),
		.io_sinks_1_bits_prot(m_axil_1_aw_bits_prot),
		.io_sinks_2_ready(m_axil_2_aw_ready),
		.io_sinks_2_valid(m_axil_2_aw_valid),
		.io_sinks_2_bits_addr(m_axil_2_aw_bits_addr),
		.io_sinks_2_bits_prot(m_axil_2_aw_bits_prot),
		.io_sinks_3_ready(m_axil_3_aw_ready),
		.io_sinks_3_valid(m_axil_3_aw_valid),
		.io_sinks_3_bits_addr(m_axil_3_aw_bits_addr),
		.io_sinks_3_bits_prot(m_axil_3_aw_bits_prot),
		.io_sinks_4_ready(m_axil_4_aw_ready),
		.io_sinks_4_valid(m_axil_4_aw_valid),
		.io_sinks_4_bits_addr(m_axil_4_aw_bits_addr),
		.io_sinks_4_bits_prot(m_axil_4_aw_bits_prot),
		.io_sinks_5_ready(m_axil_5_aw_ready),
		.io_sinks_5_valid(m_axil_5_aw_valid),
		.io_sinks_5_bits_addr(m_axil_5_aw_bits_addr),
		.io_sinks_5_bits_prot(m_axil_5_aw_bits_prot),
		.io_sinks_6_ready(m_axil_6_aw_ready),
		.io_sinks_6_valid(m_axil_6_aw_valid),
		.io_sinks_6_bits_addr(m_axil_6_aw_bits_addr),
		.io_sinks_6_bits_prot(m_axil_6_aw_bits_prot),
		.io_sinks_7_ready(m_axil_7_aw_ready),
		.io_sinks_7_valid(m_axil_7_aw_valid),
		.io_sinks_7_bits_addr(m_axil_7_aw_bits_addr),
		.io_sinks_7_bits_prot(m_axil_7_aw_bits_prot),
		.io_select_ready(_write_demux_io_select_ready),
		.io_select_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_1),
		.io_select_bits(_s_axil__sourceBuffer_1_io_deq_bits_addr[8:6])
	);
	elasticDemux_2 write_demux_1(
		.io_source_ready(_write_demux_1_io_source_ready),
		.io_source_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_source_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_source_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_sinks_0_ready(m_axil_0_w_ready),
		.io_sinks_0_valid(m_axil_0_w_valid),
		.io_sinks_0_bits_data(m_axil_0_w_bits_data),
		.io_sinks_0_bits_strb(m_axil_0_w_bits_strb),
		.io_sinks_1_ready(m_axil_1_w_ready),
		.io_sinks_1_valid(m_axil_1_w_valid),
		.io_sinks_1_bits_data(m_axil_1_w_bits_data),
		.io_sinks_1_bits_strb(m_axil_1_w_bits_strb),
		.io_sinks_2_ready(m_axil_2_w_ready),
		.io_sinks_2_valid(m_axil_2_w_valid),
		.io_sinks_2_bits_data(m_axil_2_w_bits_data),
		.io_sinks_2_bits_strb(m_axil_2_w_bits_strb),
		.io_sinks_3_ready(m_axil_3_w_ready),
		.io_sinks_3_valid(m_axil_3_w_valid),
		.io_sinks_3_bits_data(m_axil_3_w_bits_data),
		.io_sinks_3_bits_strb(m_axil_3_w_bits_strb),
		.io_sinks_4_ready(m_axil_4_w_ready),
		.io_sinks_4_valid(m_axil_4_w_valid),
		.io_sinks_4_bits_data(m_axil_4_w_bits_data),
		.io_sinks_4_bits_strb(m_axil_4_w_bits_strb),
		.io_sinks_5_ready(m_axil_5_w_ready),
		.io_sinks_5_valid(m_axil_5_w_valid),
		.io_sinks_5_bits_data(m_axil_5_w_bits_data),
		.io_sinks_5_bits_strb(m_axil_5_w_bits_strb),
		.io_sinks_6_ready(m_axil_6_w_ready),
		.io_sinks_6_valid(m_axil_6_w_valid),
		.io_sinks_6_bits_data(m_axil_6_w_bits_data),
		.io_sinks_6_bits_strb(m_axil_6_w_bits_strb),
		.io_sinks_7_ready(m_axil_7_w_ready),
		.io_sinks_7_valid(m_axil_7_w_valid),
		.io_sinks_7_bits_data(m_axil_7_w_bits_data),
		.io_sinks_7_bits_strb(m_axil_7_w_bits_strb),
		.io_select_ready(_write_demux_1_io_select_ready),
		.io_select_valid(_write_portQueueW_io_deq_valid),
		.io_select_bits(_write_portQueueW_io_deq_bits)
	);
	elasticMux_1 write_mux(
		.io_sources_0_ready(m_axil_0_b_ready),
		.io_sources_0_valid(m_axil_0_b_valid),
		.io_sources_0_bits_resp(m_axil_0_b_bits_resp),
		.io_sources_1_ready(m_axil_1_b_ready),
		.io_sources_1_valid(m_axil_1_b_valid),
		.io_sources_1_bits_resp(m_axil_1_b_bits_resp),
		.io_sources_2_ready(m_axil_2_b_ready),
		.io_sources_2_valid(m_axil_2_b_valid),
		.io_sources_2_bits_resp(m_axil_2_b_bits_resp),
		.io_sources_3_ready(m_axil_3_b_ready),
		.io_sources_3_valid(m_axil_3_b_valid),
		.io_sources_3_bits_resp(m_axil_3_b_bits_resp),
		.io_sources_4_ready(m_axil_4_b_ready),
		.io_sources_4_valid(m_axil_4_b_valid),
		.io_sources_4_bits_resp(m_axil_4_b_bits_resp),
		.io_sources_5_ready(m_axil_5_b_ready),
		.io_sources_5_valid(m_axil_5_b_valid),
		.io_sources_5_bits_resp(m_axil_5_b_bits_resp),
		.io_sources_6_ready(m_axil_6_b_ready),
		.io_sources_6_valid(m_axil_6_b_valid),
		.io_sources_6_bits_resp(m_axil_6_b_bits_resp),
		.io_sources_7_ready(m_axil_7_b_ready),
		.io_sources_7_valid(m_axil_7_b_valid),
		.io_sources_7_bits_resp(m_axil_7_b_bits_resp),
		.io_sink_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_sink_valid(_write_mux_io_sink_valid),
		.io_sink_bits_resp(_write_mux_io_sink_bits_resp),
		.io_select_ready(_write_mux_io_select_ready),
		.io_select_valid(_write_portQueueB_io_deq_valid),
		.io_select_bits(_write_portQueueB_io_deq_bits)
	);
endmodule
module SchedulerNetworkDataUnit (
	clock,
	reset,
	io_taskIn,
	io_taskOut,
	io_validIn,
	io_validOut,
	io_connSS_availableTask_ready,
	io_connSS_availableTask_valid,
	io_connSS_availableTask_bits,
	io_connSS_qOutTask_ready,
	io_connSS_qOutTask_valid,
	io_connSS_qOutTask_bits,
	io_occupied
);
	input clock;
	input reset;
	input [127:0] io_taskIn;
	output wire [127:0] io_taskOut;
	input io_validIn;
	output wire io_validOut;
	input io_connSS_availableTask_ready;
	output wire io_connSS_availableTask_valid;
	output wire [127:0] io_connSS_availableTask_bits;
	output wire io_connSS_qOutTask_ready;
	input io_connSS_qOutTask_valid;
	input [127:0] io_connSS_qOutTask_bits;
	output wire io_occupied;
	reg [127:0] taskReg;
	reg validReg;
	wire io_connSS_availableTask_valid_0 = io_connSS_availableTask_ready & io_validIn;
	wire _GEN = io_connSS_qOutTask_valid & ~io_validIn;
	always @(posedge clock)
		if (reset) begin
			taskReg <= 128'h00000000000000000000000000000000;
			validReg <= 1'h0;
		end
		else begin
			taskReg <= (io_connSS_availableTask_valid_0 ? 128'h00000000000000000000000000000000 : (_GEN ? io_connSS_qOutTask_bits : (io_validIn ? io_taskIn : 128'h00000000000000000000000000000000)));
			validReg <= ~io_connSS_availableTask_valid_0 & (_GEN | io_validIn);
		end
	assign io_taskOut = taskReg;
	assign io_validOut = validReg;
	assign io_connSS_availableTask_valid = io_connSS_availableTask_valid_0;
	assign io_connSS_availableTask_bits = (io_connSS_availableTask_valid_0 ? io_taskIn : 128'h00000000000000000000000000000000);
	assign io_connSS_qOutTask_ready = ~io_connSS_availableTask_valid_0 & _GEN;
	assign io_occupied = validReg;
endmodule
module SchedulerNetworkControlUnit (
	clock,
	reset,
	io_reqTaskIn,
	io_reqTaskOut,
	io_connSS_serveStealReq_valid,
	io_connSS_serveStealReq_ready,
	io_connSS_stealReq_valid,
	io_connSS_stealReq_ready
);
	input clock;
	input reset;
	input io_reqTaskIn;
	output wire io_reqTaskOut;
	input io_connSS_serveStealReq_valid;
	output wire io_connSS_serveStealReq_ready;
	input io_connSS_stealReq_valid;
	output wire io_connSS_stealReq_ready;
	reg stealReqReg;
	always @(posedge clock)
		if (reset)
			stealReqReg <= 1'h0;
		else
			stealReqReg <= io_reqTaskIn;
	assign io_reqTaskOut = io_connSS_stealReq_valid | (~io_connSS_serveStealReq_valid & stealReqReg);
	assign io_connSS_serveStealReq_ready = stealReqReg;
	assign io_connSS_stealReq_ready = ~stealReqReg;
endmodule
module SchedulerNetwork (
	clock,
	reset,
	io_connSS_0_ctrl_serveStealReq_valid,
	io_connSS_0_ctrl_serveStealReq_ready,
	io_connSS_0_data_availableTask_ready,
	io_connSS_0_data_availableTask_valid,
	io_connSS_0_data_availableTask_bits,
	io_connSS_0_data_qOutTask_ready,
	io_connSS_0_data_qOutTask_valid,
	io_connSS_0_data_qOutTask_bits,
	io_connSS_1_ctrl_serveStealReq_valid,
	io_connSS_1_ctrl_serveStealReq_ready,
	io_connSS_1_ctrl_stealReq_valid,
	io_connSS_1_ctrl_stealReq_ready,
	io_connSS_1_data_availableTask_ready,
	io_connSS_1_data_availableTask_valid,
	io_connSS_1_data_availableTask_bits,
	io_connSS_1_data_qOutTask_ready,
	io_connSS_1_data_qOutTask_valid,
	io_connSS_1_data_qOutTask_bits,
	io_connSS_2_ctrl_serveStealReq_valid,
	io_connSS_2_ctrl_serveStealReq_ready,
	io_connSS_2_ctrl_stealReq_valid,
	io_connSS_2_ctrl_stealReq_ready,
	io_connSS_2_data_availableTask_ready,
	io_connSS_2_data_availableTask_valid,
	io_connSS_2_data_availableTask_bits,
	io_connSS_2_data_qOutTask_ready,
	io_connSS_2_data_qOutTask_valid,
	io_connSS_2_data_qOutTask_bits,
	io_connSS_3_ctrl_serveStealReq_valid,
	io_connSS_3_ctrl_serveStealReq_ready,
	io_connSS_3_ctrl_stealReq_valid,
	io_connSS_3_ctrl_stealReq_ready,
	io_connSS_3_data_availableTask_ready,
	io_connSS_3_data_availableTask_valid,
	io_connSS_3_data_availableTask_bits,
	io_connSS_3_data_qOutTask_ready,
	io_connSS_3_data_qOutTask_valid,
	io_connSS_3_data_qOutTask_bits,
	io_connSS_4_ctrl_serveStealReq_valid,
	io_connSS_4_ctrl_serveStealReq_ready,
	io_connSS_4_ctrl_stealReq_valid,
	io_connSS_4_ctrl_stealReq_ready,
	io_connSS_4_data_availableTask_ready,
	io_connSS_4_data_availableTask_valid,
	io_connSS_4_data_availableTask_bits,
	io_connSS_4_data_qOutTask_ready,
	io_connSS_4_data_qOutTask_valid,
	io_connSS_4_data_qOutTask_bits,
	io_connSS_5_ctrl_serveStealReq_valid,
	io_connSS_5_ctrl_serveStealReq_ready,
	io_connSS_5_ctrl_stealReq_valid,
	io_connSS_5_ctrl_stealReq_ready,
	io_connSS_5_data_availableTask_ready,
	io_connSS_5_data_availableTask_valid,
	io_connSS_5_data_availableTask_bits,
	io_connSS_5_data_qOutTask_ready,
	io_connSS_5_data_qOutTask_valid,
	io_connSS_5_data_qOutTask_bits,
	io_connSS_6_ctrl_serveStealReq_valid,
	io_connSS_6_ctrl_serveStealReq_ready,
	io_connSS_6_ctrl_stealReq_valid,
	io_connSS_6_ctrl_stealReq_ready,
	io_connSS_6_data_availableTask_ready,
	io_connSS_6_data_availableTask_valid,
	io_connSS_6_data_availableTask_bits,
	io_connSS_6_data_qOutTask_ready,
	io_connSS_6_data_qOutTask_valid,
	io_connSS_6_data_qOutTask_bits,
	io_connSS_7_ctrl_serveStealReq_valid,
	io_connSS_7_ctrl_serveStealReq_ready,
	io_connSS_7_ctrl_stealReq_valid,
	io_connSS_7_ctrl_stealReq_ready,
	io_connSS_7_data_availableTask_ready,
	io_connSS_7_data_availableTask_valid,
	io_connSS_7_data_availableTask_bits,
	io_connSS_7_data_qOutTask_ready,
	io_connSS_7_data_qOutTask_valid,
	io_connSS_7_data_qOutTask_bits,
	io_connSS_8_ctrl_serveStealReq_valid,
	io_connSS_8_ctrl_serveStealReq_ready,
	io_connSS_8_ctrl_stealReq_valid,
	io_connSS_8_ctrl_stealReq_ready,
	io_connSS_8_data_availableTask_ready,
	io_connSS_8_data_availableTask_valid,
	io_connSS_8_data_availableTask_bits,
	io_connSS_8_data_qOutTask_ready,
	io_connSS_8_data_qOutTask_valid,
	io_connSS_8_data_qOutTask_bits,
	io_connSS_9_ctrl_serveStealReq_valid,
	io_connSS_9_ctrl_serveStealReq_ready,
	io_connSS_9_ctrl_stealReq_valid,
	io_connSS_9_ctrl_stealReq_ready,
	io_connSS_9_data_availableTask_ready,
	io_connSS_9_data_availableTask_valid,
	io_connSS_9_data_availableTask_bits,
	io_connSS_9_data_qOutTask_ready,
	io_connSS_9_data_qOutTask_valid,
	io_connSS_9_data_qOutTask_bits,
	io_connSS_10_ctrl_serveStealReq_valid,
	io_connSS_10_ctrl_serveStealReq_ready,
	io_connSS_10_ctrl_stealReq_valid,
	io_connSS_10_ctrl_stealReq_ready,
	io_connSS_10_data_availableTask_ready,
	io_connSS_10_data_availableTask_valid,
	io_connSS_10_data_availableTask_bits,
	io_connSS_10_data_qOutTask_ready,
	io_connSS_10_data_qOutTask_valid,
	io_connSS_10_data_qOutTask_bits,
	io_connSS_11_ctrl_serveStealReq_valid,
	io_connSS_11_ctrl_serveStealReq_ready,
	io_connSS_11_ctrl_stealReq_valid,
	io_connSS_11_ctrl_stealReq_ready,
	io_connSS_11_data_availableTask_ready,
	io_connSS_11_data_availableTask_valid,
	io_connSS_11_data_availableTask_bits,
	io_connSS_11_data_qOutTask_ready,
	io_connSS_11_data_qOutTask_valid,
	io_connSS_11_data_qOutTask_bits,
	io_connSS_12_ctrl_serveStealReq_valid,
	io_connSS_12_ctrl_serveStealReq_ready,
	io_connSS_12_ctrl_stealReq_valid,
	io_connSS_12_ctrl_stealReq_ready,
	io_connSS_12_data_availableTask_ready,
	io_connSS_12_data_availableTask_valid,
	io_connSS_12_data_availableTask_bits,
	io_connSS_12_data_qOutTask_ready,
	io_connSS_12_data_qOutTask_valid,
	io_connSS_12_data_qOutTask_bits,
	io_connSS_13_ctrl_serveStealReq_valid,
	io_connSS_13_ctrl_serveStealReq_ready,
	io_connSS_13_ctrl_stealReq_valid,
	io_connSS_13_ctrl_stealReq_ready,
	io_connSS_13_data_availableTask_ready,
	io_connSS_13_data_availableTask_valid,
	io_connSS_13_data_availableTask_bits,
	io_connSS_13_data_qOutTask_ready,
	io_connSS_13_data_qOutTask_valid,
	io_connSS_13_data_qOutTask_bits,
	io_connSS_14_ctrl_serveStealReq_valid,
	io_connSS_14_ctrl_serveStealReq_ready,
	io_connSS_14_ctrl_stealReq_valid,
	io_connSS_14_ctrl_stealReq_ready,
	io_connSS_14_data_availableTask_ready,
	io_connSS_14_data_availableTask_valid,
	io_connSS_14_data_availableTask_bits,
	io_connSS_14_data_qOutTask_ready,
	io_connSS_14_data_qOutTask_valid,
	io_connSS_14_data_qOutTask_bits,
	io_connSS_15_ctrl_serveStealReq_valid,
	io_connSS_15_ctrl_serveStealReq_ready,
	io_connSS_15_ctrl_stealReq_valid,
	io_connSS_15_ctrl_stealReq_ready,
	io_connSS_15_data_availableTask_ready,
	io_connSS_15_data_availableTask_valid,
	io_connSS_15_data_availableTask_bits,
	io_connSS_15_data_qOutTask_ready,
	io_connSS_15_data_qOutTask_valid,
	io_connSS_15_data_qOutTask_bits,
	io_connSS_16_ctrl_serveStealReq_valid,
	io_connSS_16_ctrl_serveStealReq_ready,
	io_connSS_16_ctrl_stealReq_valid,
	io_connSS_16_ctrl_stealReq_ready,
	io_connSS_16_data_availableTask_ready,
	io_connSS_16_data_availableTask_valid,
	io_connSS_16_data_availableTask_bits,
	io_connSS_16_data_qOutTask_ready,
	io_connSS_16_data_qOutTask_valid,
	io_connSS_16_data_qOutTask_bits,
	io_connSS_17_ctrl_serveStealReq_valid,
	io_connSS_17_ctrl_serveStealReq_ready,
	io_connSS_17_ctrl_stealReq_valid,
	io_connSS_17_ctrl_stealReq_ready,
	io_connSS_17_data_availableTask_ready,
	io_connSS_17_data_availableTask_valid,
	io_connSS_17_data_availableTask_bits,
	io_connSS_17_data_qOutTask_ready,
	io_connSS_17_data_qOutTask_valid,
	io_connSS_17_data_qOutTask_bits,
	io_connSS_18_ctrl_serveStealReq_valid,
	io_connSS_18_ctrl_serveStealReq_ready,
	io_connSS_18_ctrl_stealReq_valid,
	io_connSS_18_ctrl_stealReq_ready,
	io_connSS_18_data_availableTask_ready,
	io_connSS_18_data_availableTask_valid,
	io_connSS_18_data_availableTask_bits,
	io_connSS_18_data_qOutTask_ready,
	io_connSS_18_data_qOutTask_valid,
	io_connSS_18_data_qOutTask_bits,
	io_connSS_19_ctrl_serveStealReq_valid,
	io_connSS_19_ctrl_serveStealReq_ready,
	io_connSS_19_ctrl_stealReq_valid,
	io_connSS_19_ctrl_stealReq_ready,
	io_connSS_19_data_availableTask_ready,
	io_connSS_19_data_availableTask_valid,
	io_connSS_19_data_availableTask_bits,
	io_connSS_19_data_qOutTask_ready,
	io_connSS_19_data_qOutTask_valid,
	io_connSS_19_data_qOutTask_bits,
	io_connSS_20_ctrl_serveStealReq_valid,
	io_connSS_20_ctrl_serveStealReq_ready,
	io_connSS_20_ctrl_stealReq_valid,
	io_connSS_20_ctrl_stealReq_ready,
	io_connSS_20_data_availableTask_ready,
	io_connSS_20_data_availableTask_valid,
	io_connSS_20_data_availableTask_bits,
	io_connSS_20_data_qOutTask_ready,
	io_connSS_20_data_qOutTask_valid,
	io_connSS_20_data_qOutTask_bits,
	io_connSS_21_ctrl_serveStealReq_valid,
	io_connSS_21_ctrl_serveStealReq_ready,
	io_connSS_21_ctrl_stealReq_valid,
	io_connSS_21_ctrl_stealReq_ready,
	io_connSS_21_data_availableTask_ready,
	io_connSS_21_data_availableTask_valid,
	io_connSS_21_data_availableTask_bits,
	io_connSS_21_data_qOutTask_ready,
	io_connSS_21_data_qOutTask_valid,
	io_connSS_21_data_qOutTask_bits,
	io_connSS_22_ctrl_serveStealReq_valid,
	io_connSS_22_ctrl_serveStealReq_ready,
	io_connSS_22_ctrl_stealReq_valid,
	io_connSS_22_ctrl_stealReq_ready,
	io_connSS_22_data_availableTask_ready,
	io_connSS_22_data_availableTask_valid,
	io_connSS_22_data_availableTask_bits,
	io_connSS_22_data_qOutTask_ready,
	io_connSS_22_data_qOutTask_valid,
	io_connSS_22_data_qOutTask_bits,
	io_connSS_23_ctrl_serveStealReq_valid,
	io_connSS_23_ctrl_serveStealReq_ready,
	io_connSS_23_ctrl_stealReq_valid,
	io_connSS_23_ctrl_stealReq_ready,
	io_connSS_23_data_availableTask_ready,
	io_connSS_23_data_availableTask_valid,
	io_connSS_23_data_availableTask_bits,
	io_connSS_23_data_qOutTask_ready,
	io_connSS_23_data_qOutTask_valid,
	io_connSS_23_data_qOutTask_bits,
	io_connSS_24_ctrl_serveStealReq_valid,
	io_connSS_24_ctrl_serveStealReq_ready,
	io_connSS_24_ctrl_stealReq_valid,
	io_connSS_24_ctrl_stealReq_ready,
	io_connSS_24_data_availableTask_ready,
	io_connSS_24_data_availableTask_valid,
	io_connSS_24_data_availableTask_bits,
	io_connSS_24_data_qOutTask_ready,
	io_connSS_24_data_qOutTask_valid,
	io_connSS_24_data_qOutTask_bits,
	io_connSS_25_ctrl_serveStealReq_valid,
	io_connSS_25_ctrl_serveStealReq_ready,
	io_connSS_25_ctrl_stealReq_valid,
	io_connSS_25_ctrl_stealReq_ready,
	io_connSS_25_data_availableTask_ready,
	io_connSS_25_data_availableTask_valid,
	io_connSS_25_data_availableTask_bits,
	io_connSS_25_data_qOutTask_ready,
	io_connSS_25_data_qOutTask_valid,
	io_connSS_25_data_qOutTask_bits,
	io_connSS_26_ctrl_serveStealReq_valid,
	io_connSS_26_ctrl_serveStealReq_ready,
	io_connSS_26_ctrl_stealReq_valid,
	io_connSS_26_ctrl_stealReq_ready,
	io_connSS_26_data_availableTask_ready,
	io_connSS_26_data_availableTask_valid,
	io_connSS_26_data_availableTask_bits,
	io_connSS_26_data_qOutTask_ready,
	io_connSS_26_data_qOutTask_valid,
	io_connSS_26_data_qOutTask_bits,
	io_connSS_27_ctrl_serveStealReq_valid,
	io_connSS_27_ctrl_serveStealReq_ready,
	io_connSS_27_ctrl_stealReq_valid,
	io_connSS_27_ctrl_stealReq_ready,
	io_connSS_27_data_availableTask_ready,
	io_connSS_27_data_availableTask_valid,
	io_connSS_27_data_availableTask_bits,
	io_connSS_27_data_qOutTask_ready,
	io_connSS_27_data_qOutTask_valid,
	io_connSS_27_data_qOutTask_bits,
	io_connSS_28_ctrl_serveStealReq_valid,
	io_connSS_28_ctrl_serveStealReq_ready,
	io_connSS_28_ctrl_stealReq_valid,
	io_connSS_28_ctrl_stealReq_ready,
	io_connSS_28_data_availableTask_ready,
	io_connSS_28_data_availableTask_valid,
	io_connSS_28_data_availableTask_bits,
	io_connSS_28_data_qOutTask_ready,
	io_connSS_28_data_qOutTask_valid,
	io_connSS_28_data_qOutTask_bits,
	io_connSS_29_ctrl_serveStealReq_valid,
	io_connSS_29_ctrl_serveStealReq_ready,
	io_connSS_29_ctrl_stealReq_valid,
	io_connSS_29_ctrl_stealReq_ready,
	io_connSS_29_data_availableTask_ready,
	io_connSS_29_data_availableTask_valid,
	io_connSS_29_data_availableTask_bits,
	io_connSS_29_data_qOutTask_ready,
	io_connSS_29_data_qOutTask_valid,
	io_connSS_29_data_qOutTask_bits,
	io_connSS_30_ctrl_serveStealReq_valid,
	io_connSS_30_ctrl_serveStealReq_ready,
	io_connSS_30_ctrl_stealReq_valid,
	io_connSS_30_ctrl_stealReq_ready,
	io_connSS_30_data_availableTask_ready,
	io_connSS_30_data_availableTask_valid,
	io_connSS_30_data_availableTask_bits,
	io_connSS_30_data_qOutTask_ready,
	io_connSS_30_data_qOutTask_valid,
	io_connSS_30_data_qOutTask_bits,
	io_connSS_31_ctrl_serveStealReq_valid,
	io_connSS_31_ctrl_serveStealReq_ready,
	io_connSS_31_ctrl_stealReq_valid,
	io_connSS_31_ctrl_stealReq_ready,
	io_connSS_31_data_availableTask_ready,
	io_connSS_31_data_availableTask_valid,
	io_connSS_31_data_availableTask_bits,
	io_connSS_31_data_qOutTask_ready,
	io_connSS_31_data_qOutTask_valid,
	io_connSS_31_data_qOutTask_bits,
	io_connSS_32_ctrl_serveStealReq_valid,
	io_connSS_32_ctrl_serveStealReq_ready,
	io_connSS_32_ctrl_stealReq_valid,
	io_connSS_32_ctrl_stealReq_ready,
	io_connSS_32_data_availableTask_ready,
	io_connSS_32_data_availableTask_valid,
	io_connSS_32_data_availableTask_bits,
	io_connSS_32_data_qOutTask_ready,
	io_connSS_32_data_qOutTask_valid,
	io_connSS_32_data_qOutTask_bits,
	io_connSS_33_ctrl_serveStealReq_valid,
	io_connSS_33_ctrl_serveStealReq_ready,
	io_connSS_33_data_availableTask_ready,
	io_connSS_33_data_availableTask_valid,
	io_connSS_33_data_availableTask_bits,
	io_connSS_33_data_qOutTask_ready,
	io_connSS_33_data_qOutTask_valid,
	io_connSS_33_data_qOutTask_bits,
	io_connSS_34_ctrl_serveStealReq_valid,
	io_connSS_34_ctrl_serveStealReq_ready,
	io_connSS_34_ctrl_stealReq_valid,
	io_connSS_34_ctrl_stealReq_ready,
	io_connSS_34_data_availableTask_ready,
	io_connSS_34_data_availableTask_valid,
	io_connSS_34_data_availableTask_bits,
	io_connSS_34_data_qOutTask_ready,
	io_connSS_34_data_qOutTask_valid,
	io_connSS_34_data_qOutTask_bits,
	io_connSS_35_ctrl_serveStealReq_valid,
	io_connSS_35_ctrl_serveStealReq_ready,
	io_connSS_35_ctrl_stealReq_valid,
	io_connSS_35_ctrl_stealReq_ready,
	io_connSS_35_data_availableTask_ready,
	io_connSS_35_data_availableTask_valid,
	io_connSS_35_data_availableTask_bits,
	io_connSS_35_data_qOutTask_ready,
	io_connSS_35_data_qOutTask_valid,
	io_connSS_35_data_qOutTask_bits,
	io_connSS_36_ctrl_serveStealReq_valid,
	io_connSS_36_ctrl_serveStealReq_ready,
	io_connSS_36_ctrl_stealReq_valid,
	io_connSS_36_ctrl_stealReq_ready,
	io_connSS_36_data_availableTask_ready,
	io_connSS_36_data_availableTask_valid,
	io_connSS_36_data_availableTask_bits,
	io_connSS_36_data_qOutTask_ready,
	io_connSS_36_data_qOutTask_valid,
	io_connSS_36_data_qOutTask_bits,
	io_connSS_37_ctrl_serveStealReq_valid,
	io_connSS_37_ctrl_serveStealReq_ready,
	io_connSS_37_ctrl_stealReq_valid,
	io_connSS_37_ctrl_stealReq_ready,
	io_connSS_37_data_availableTask_ready,
	io_connSS_37_data_availableTask_valid,
	io_connSS_37_data_availableTask_bits,
	io_connSS_37_data_qOutTask_ready,
	io_connSS_37_data_qOutTask_valid,
	io_connSS_37_data_qOutTask_bits,
	io_connSS_38_ctrl_serveStealReq_valid,
	io_connSS_38_ctrl_serveStealReq_ready,
	io_connSS_38_ctrl_stealReq_valid,
	io_connSS_38_ctrl_stealReq_ready,
	io_connSS_38_data_availableTask_ready,
	io_connSS_38_data_availableTask_valid,
	io_connSS_38_data_availableTask_bits,
	io_connSS_38_data_qOutTask_ready,
	io_connSS_38_data_qOutTask_valid,
	io_connSS_38_data_qOutTask_bits,
	io_connSS_39_ctrl_serveStealReq_valid,
	io_connSS_39_ctrl_serveStealReq_ready,
	io_connSS_39_ctrl_stealReq_valid,
	io_connSS_39_ctrl_stealReq_ready,
	io_connSS_39_data_availableTask_ready,
	io_connSS_39_data_availableTask_valid,
	io_connSS_39_data_availableTask_bits,
	io_connSS_39_data_qOutTask_ready,
	io_connSS_39_data_qOutTask_valid,
	io_connSS_39_data_qOutTask_bits,
	io_connSS_40_ctrl_serveStealReq_valid,
	io_connSS_40_ctrl_serveStealReq_ready,
	io_connSS_40_ctrl_stealReq_valid,
	io_connSS_40_ctrl_stealReq_ready,
	io_connSS_40_data_availableTask_ready,
	io_connSS_40_data_availableTask_valid,
	io_connSS_40_data_availableTask_bits,
	io_connSS_40_data_qOutTask_ready,
	io_connSS_40_data_qOutTask_valid,
	io_connSS_40_data_qOutTask_bits,
	io_connSS_41_ctrl_serveStealReq_valid,
	io_connSS_41_ctrl_serveStealReq_ready,
	io_connSS_41_ctrl_stealReq_valid,
	io_connSS_41_ctrl_stealReq_ready,
	io_connSS_41_data_availableTask_ready,
	io_connSS_41_data_availableTask_valid,
	io_connSS_41_data_availableTask_bits,
	io_connSS_41_data_qOutTask_ready,
	io_connSS_41_data_qOutTask_valid,
	io_connSS_41_data_qOutTask_bits,
	io_connSS_42_ctrl_serveStealReq_valid,
	io_connSS_42_ctrl_serveStealReq_ready,
	io_connSS_42_ctrl_stealReq_valid,
	io_connSS_42_ctrl_stealReq_ready,
	io_connSS_42_data_availableTask_ready,
	io_connSS_42_data_availableTask_valid,
	io_connSS_42_data_availableTask_bits,
	io_connSS_42_data_qOutTask_ready,
	io_connSS_42_data_qOutTask_valid,
	io_connSS_42_data_qOutTask_bits,
	io_connSS_43_ctrl_serveStealReq_valid,
	io_connSS_43_ctrl_serveStealReq_ready,
	io_connSS_43_ctrl_stealReq_valid,
	io_connSS_43_ctrl_stealReq_ready,
	io_connSS_43_data_availableTask_ready,
	io_connSS_43_data_availableTask_valid,
	io_connSS_43_data_availableTask_bits,
	io_connSS_43_data_qOutTask_ready,
	io_connSS_43_data_qOutTask_valid,
	io_connSS_43_data_qOutTask_bits,
	io_connSS_44_ctrl_serveStealReq_valid,
	io_connSS_44_ctrl_serveStealReq_ready,
	io_connSS_44_ctrl_stealReq_valid,
	io_connSS_44_ctrl_stealReq_ready,
	io_connSS_44_data_availableTask_ready,
	io_connSS_44_data_availableTask_valid,
	io_connSS_44_data_availableTask_bits,
	io_connSS_44_data_qOutTask_ready,
	io_connSS_44_data_qOutTask_valid,
	io_connSS_44_data_qOutTask_bits,
	io_connSS_45_ctrl_serveStealReq_valid,
	io_connSS_45_ctrl_serveStealReq_ready,
	io_connSS_45_ctrl_stealReq_valid,
	io_connSS_45_ctrl_stealReq_ready,
	io_connSS_45_data_availableTask_ready,
	io_connSS_45_data_availableTask_valid,
	io_connSS_45_data_availableTask_bits,
	io_connSS_45_data_qOutTask_ready,
	io_connSS_45_data_qOutTask_valid,
	io_connSS_45_data_qOutTask_bits,
	io_connSS_46_ctrl_serveStealReq_valid,
	io_connSS_46_ctrl_serveStealReq_ready,
	io_connSS_46_ctrl_stealReq_valid,
	io_connSS_46_ctrl_stealReq_ready,
	io_connSS_46_data_availableTask_ready,
	io_connSS_46_data_availableTask_valid,
	io_connSS_46_data_availableTask_bits,
	io_connSS_46_data_qOutTask_ready,
	io_connSS_46_data_qOutTask_valid,
	io_connSS_46_data_qOutTask_bits,
	io_connSS_47_ctrl_serveStealReq_valid,
	io_connSS_47_ctrl_serveStealReq_ready,
	io_connSS_47_ctrl_stealReq_valid,
	io_connSS_47_ctrl_stealReq_ready,
	io_connSS_47_data_availableTask_ready,
	io_connSS_47_data_availableTask_valid,
	io_connSS_47_data_availableTask_bits,
	io_connSS_47_data_qOutTask_ready,
	io_connSS_47_data_qOutTask_valid,
	io_connSS_47_data_qOutTask_bits,
	io_connSS_48_ctrl_serveStealReq_valid,
	io_connSS_48_ctrl_serveStealReq_ready,
	io_connSS_48_ctrl_stealReq_valid,
	io_connSS_48_ctrl_stealReq_ready,
	io_connSS_48_data_availableTask_ready,
	io_connSS_48_data_availableTask_valid,
	io_connSS_48_data_availableTask_bits,
	io_connSS_48_data_qOutTask_ready,
	io_connSS_48_data_qOutTask_valid,
	io_connSS_48_data_qOutTask_bits,
	io_connSS_49_ctrl_serveStealReq_valid,
	io_connSS_49_ctrl_serveStealReq_ready,
	io_connSS_49_ctrl_stealReq_valid,
	io_connSS_49_ctrl_stealReq_ready,
	io_connSS_49_data_availableTask_ready,
	io_connSS_49_data_availableTask_valid,
	io_connSS_49_data_availableTask_bits,
	io_connSS_49_data_qOutTask_ready,
	io_connSS_49_data_qOutTask_valid,
	io_connSS_49_data_qOutTask_bits,
	io_connSS_50_ctrl_serveStealReq_valid,
	io_connSS_50_ctrl_serveStealReq_ready,
	io_connSS_50_ctrl_stealReq_valid,
	io_connSS_50_ctrl_stealReq_ready,
	io_connSS_50_data_availableTask_ready,
	io_connSS_50_data_availableTask_valid,
	io_connSS_50_data_availableTask_bits,
	io_connSS_50_data_qOutTask_ready,
	io_connSS_50_data_qOutTask_valid,
	io_connSS_50_data_qOutTask_bits,
	io_connSS_51_ctrl_serveStealReq_valid,
	io_connSS_51_ctrl_serveStealReq_ready,
	io_connSS_51_ctrl_stealReq_valid,
	io_connSS_51_ctrl_stealReq_ready,
	io_connSS_51_data_availableTask_ready,
	io_connSS_51_data_availableTask_valid,
	io_connSS_51_data_availableTask_bits,
	io_connSS_51_data_qOutTask_ready,
	io_connSS_51_data_qOutTask_valid,
	io_connSS_51_data_qOutTask_bits,
	io_connSS_52_ctrl_serveStealReq_valid,
	io_connSS_52_ctrl_serveStealReq_ready,
	io_connSS_52_ctrl_stealReq_valid,
	io_connSS_52_ctrl_stealReq_ready,
	io_connSS_52_data_availableTask_ready,
	io_connSS_52_data_availableTask_valid,
	io_connSS_52_data_availableTask_bits,
	io_connSS_52_data_qOutTask_ready,
	io_connSS_52_data_qOutTask_valid,
	io_connSS_52_data_qOutTask_bits,
	io_connSS_53_ctrl_serveStealReq_valid,
	io_connSS_53_ctrl_serveStealReq_ready,
	io_connSS_53_ctrl_stealReq_valid,
	io_connSS_53_ctrl_stealReq_ready,
	io_connSS_53_data_availableTask_ready,
	io_connSS_53_data_availableTask_valid,
	io_connSS_53_data_availableTask_bits,
	io_connSS_53_data_qOutTask_ready,
	io_connSS_53_data_qOutTask_valid,
	io_connSS_53_data_qOutTask_bits,
	io_connSS_54_ctrl_serveStealReq_valid,
	io_connSS_54_ctrl_serveStealReq_ready,
	io_connSS_54_ctrl_stealReq_valid,
	io_connSS_54_ctrl_stealReq_ready,
	io_connSS_54_data_availableTask_ready,
	io_connSS_54_data_availableTask_valid,
	io_connSS_54_data_availableTask_bits,
	io_connSS_54_data_qOutTask_ready,
	io_connSS_54_data_qOutTask_valid,
	io_connSS_54_data_qOutTask_bits,
	io_connSS_55_ctrl_serveStealReq_valid,
	io_connSS_55_ctrl_serveStealReq_ready,
	io_connSS_55_ctrl_stealReq_valid,
	io_connSS_55_ctrl_stealReq_ready,
	io_connSS_55_data_availableTask_ready,
	io_connSS_55_data_availableTask_valid,
	io_connSS_55_data_availableTask_bits,
	io_connSS_55_data_qOutTask_ready,
	io_connSS_55_data_qOutTask_valid,
	io_connSS_55_data_qOutTask_bits,
	io_connSS_56_ctrl_serveStealReq_valid,
	io_connSS_56_ctrl_serveStealReq_ready,
	io_connSS_56_ctrl_stealReq_valid,
	io_connSS_56_ctrl_stealReq_ready,
	io_connSS_56_data_availableTask_ready,
	io_connSS_56_data_availableTask_valid,
	io_connSS_56_data_availableTask_bits,
	io_connSS_56_data_qOutTask_ready,
	io_connSS_56_data_qOutTask_valid,
	io_connSS_56_data_qOutTask_bits,
	io_connSS_57_ctrl_serveStealReq_valid,
	io_connSS_57_ctrl_serveStealReq_ready,
	io_connSS_57_ctrl_stealReq_valid,
	io_connSS_57_ctrl_stealReq_ready,
	io_connSS_57_data_availableTask_ready,
	io_connSS_57_data_availableTask_valid,
	io_connSS_57_data_availableTask_bits,
	io_connSS_57_data_qOutTask_ready,
	io_connSS_57_data_qOutTask_valid,
	io_connSS_57_data_qOutTask_bits,
	io_connSS_58_ctrl_serveStealReq_valid,
	io_connSS_58_ctrl_serveStealReq_ready,
	io_connSS_58_ctrl_stealReq_valid,
	io_connSS_58_ctrl_stealReq_ready,
	io_connSS_58_data_availableTask_ready,
	io_connSS_58_data_availableTask_valid,
	io_connSS_58_data_availableTask_bits,
	io_connSS_58_data_qOutTask_ready,
	io_connSS_58_data_qOutTask_valid,
	io_connSS_58_data_qOutTask_bits,
	io_connSS_59_ctrl_serveStealReq_valid,
	io_connSS_59_ctrl_serveStealReq_ready,
	io_connSS_59_ctrl_stealReq_valid,
	io_connSS_59_ctrl_stealReq_ready,
	io_connSS_59_data_availableTask_ready,
	io_connSS_59_data_availableTask_valid,
	io_connSS_59_data_availableTask_bits,
	io_connSS_59_data_qOutTask_ready,
	io_connSS_59_data_qOutTask_valid,
	io_connSS_59_data_qOutTask_bits,
	io_connSS_60_ctrl_serveStealReq_valid,
	io_connSS_60_ctrl_serveStealReq_ready,
	io_connSS_60_ctrl_stealReq_valid,
	io_connSS_60_ctrl_stealReq_ready,
	io_connSS_60_data_availableTask_ready,
	io_connSS_60_data_availableTask_valid,
	io_connSS_60_data_availableTask_bits,
	io_connSS_60_data_qOutTask_ready,
	io_connSS_60_data_qOutTask_valid,
	io_connSS_60_data_qOutTask_bits,
	io_connSS_61_ctrl_serveStealReq_valid,
	io_connSS_61_ctrl_serveStealReq_ready,
	io_connSS_61_ctrl_stealReq_valid,
	io_connSS_61_ctrl_stealReq_ready,
	io_connSS_61_data_availableTask_ready,
	io_connSS_61_data_availableTask_valid,
	io_connSS_61_data_availableTask_bits,
	io_connSS_61_data_qOutTask_ready,
	io_connSS_61_data_qOutTask_valid,
	io_connSS_61_data_qOutTask_bits,
	io_connSS_62_ctrl_serveStealReq_valid,
	io_connSS_62_ctrl_serveStealReq_ready,
	io_connSS_62_ctrl_stealReq_valid,
	io_connSS_62_ctrl_stealReq_ready,
	io_connSS_62_data_availableTask_ready,
	io_connSS_62_data_availableTask_valid,
	io_connSS_62_data_availableTask_bits,
	io_connSS_62_data_qOutTask_ready,
	io_connSS_62_data_qOutTask_valid,
	io_connSS_62_data_qOutTask_bits,
	io_connSS_63_ctrl_serveStealReq_valid,
	io_connSS_63_ctrl_serveStealReq_ready,
	io_connSS_63_ctrl_stealReq_valid,
	io_connSS_63_ctrl_stealReq_ready,
	io_connSS_63_data_availableTask_ready,
	io_connSS_63_data_availableTask_valid,
	io_connSS_63_data_availableTask_bits,
	io_connSS_63_data_qOutTask_ready,
	io_connSS_63_data_qOutTask_valid,
	io_connSS_63_data_qOutTask_bits,
	io_connSS_64_ctrl_serveStealReq_valid,
	io_connSS_64_ctrl_serveStealReq_ready,
	io_connSS_64_ctrl_stealReq_valid,
	io_connSS_64_ctrl_stealReq_ready,
	io_connSS_64_data_availableTask_ready,
	io_connSS_64_data_availableTask_valid,
	io_connSS_64_data_availableTask_bits,
	io_connSS_64_data_qOutTask_ready,
	io_connSS_64_data_qOutTask_valid,
	io_connSS_64_data_qOutTask_bits,
	io_connSS_65_ctrl_serveStealReq_valid,
	io_connSS_65_ctrl_serveStealReq_ready,
	io_connSS_65_ctrl_stealReq_valid,
	io_connSS_65_ctrl_stealReq_ready,
	io_connSS_65_data_availableTask_ready,
	io_connSS_65_data_availableTask_valid,
	io_connSS_65_data_availableTask_bits,
	io_connSS_65_data_qOutTask_ready,
	io_connSS_65_data_qOutTask_valid,
	io_connSS_65_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0,
	io_ntwDataUnitOccupancyVSS_1
);
	input clock;
	input reset;
	input io_connSS_0_ctrl_serveStealReq_valid;
	output wire io_connSS_0_ctrl_serveStealReq_ready;
	input io_connSS_0_data_availableTask_ready;
	output wire io_connSS_0_data_availableTask_valid;
	output wire [127:0] io_connSS_0_data_availableTask_bits;
	output wire io_connSS_0_data_qOutTask_ready;
	input io_connSS_0_data_qOutTask_valid;
	input [127:0] io_connSS_0_data_qOutTask_bits;
	input io_connSS_1_ctrl_serveStealReq_valid;
	output wire io_connSS_1_ctrl_serveStealReq_ready;
	input io_connSS_1_ctrl_stealReq_valid;
	output wire io_connSS_1_ctrl_stealReq_ready;
	input io_connSS_1_data_availableTask_ready;
	output wire io_connSS_1_data_availableTask_valid;
	output wire [127:0] io_connSS_1_data_availableTask_bits;
	output wire io_connSS_1_data_qOutTask_ready;
	input io_connSS_1_data_qOutTask_valid;
	input [127:0] io_connSS_1_data_qOutTask_bits;
	input io_connSS_2_ctrl_serveStealReq_valid;
	output wire io_connSS_2_ctrl_serveStealReq_ready;
	input io_connSS_2_ctrl_stealReq_valid;
	output wire io_connSS_2_ctrl_stealReq_ready;
	input io_connSS_2_data_availableTask_ready;
	output wire io_connSS_2_data_availableTask_valid;
	output wire [127:0] io_connSS_2_data_availableTask_bits;
	output wire io_connSS_2_data_qOutTask_ready;
	input io_connSS_2_data_qOutTask_valid;
	input [127:0] io_connSS_2_data_qOutTask_bits;
	input io_connSS_3_ctrl_serveStealReq_valid;
	output wire io_connSS_3_ctrl_serveStealReq_ready;
	input io_connSS_3_ctrl_stealReq_valid;
	output wire io_connSS_3_ctrl_stealReq_ready;
	input io_connSS_3_data_availableTask_ready;
	output wire io_connSS_3_data_availableTask_valid;
	output wire [127:0] io_connSS_3_data_availableTask_bits;
	output wire io_connSS_3_data_qOutTask_ready;
	input io_connSS_3_data_qOutTask_valid;
	input [127:0] io_connSS_3_data_qOutTask_bits;
	input io_connSS_4_ctrl_serveStealReq_valid;
	output wire io_connSS_4_ctrl_serveStealReq_ready;
	input io_connSS_4_ctrl_stealReq_valid;
	output wire io_connSS_4_ctrl_stealReq_ready;
	input io_connSS_4_data_availableTask_ready;
	output wire io_connSS_4_data_availableTask_valid;
	output wire [127:0] io_connSS_4_data_availableTask_bits;
	output wire io_connSS_4_data_qOutTask_ready;
	input io_connSS_4_data_qOutTask_valid;
	input [127:0] io_connSS_4_data_qOutTask_bits;
	input io_connSS_5_ctrl_serveStealReq_valid;
	output wire io_connSS_5_ctrl_serveStealReq_ready;
	input io_connSS_5_ctrl_stealReq_valid;
	output wire io_connSS_5_ctrl_stealReq_ready;
	input io_connSS_5_data_availableTask_ready;
	output wire io_connSS_5_data_availableTask_valid;
	output wire [127:0] io_connSS_5_data_availableTask_bits;
	output wire io_connSS_5_data_qOutTask_ready;
	input io_connSS_5_data_qOutTask_valid;
	input [127:0] io_connSS_5_data_qOutTask_bits;
	input io_connSS_6_ctrl_serveStealReq_valid;
	output wire io_connSS_6_ctrl_serveStealReq_ready;
	input io_connSS_6_ctrl_stealReq_valid;
	output wire io_connSS_6_ctrl_stealReq_ready;
	input io_connSS_6_data_availableTask_ready;
	output wire io_connSS_6_data_availableTask_valid;
	output wire [127:0] io_connSS_6_data_availableTask_bits;
	output wire io_connSS_6_data_qOutTask_ready;
	input io_connSS_6_data_qOutTask_valid;
	input [127:0] io_connSS_6_data_qOutTask_bits;
	input io_connSS_7_ctrl_serveStealReq_valid;
	output wire io_connSS_7_ctrl_serveStealReq_ready;
	input io_connSS_7_ctrl_stealReq_valid;
	output wire io_connSS_7_ctrl_stealReq_ready;
	input io_connSS_7_data_availableTask_ready;
	output wire io_connSS_7_data_availableTask_valid;
	output wire [127:0] io_connSS_7_data_availableTask_bits;
	output wire io_connSS_7_data_qOutTask_ready;
	input io_connSS_7_data_qOutTask_valid;
	input [127:0] io_connSS_7_data_qOutTask_bits;
	input io_connSS_8_ctrl_serveStealReq_valid;
	output wire io_connSS_8_ctrl_serveStealReq_ready;
	input io_connSS_8_ctrl_stealReq_valid;
	output wire io_connSS_8_ctrl_stealReq_ready;
	input io_connSS_8_data_availableTask_ready;
	output wire io_connSS_8_data_availableTask_valid;
	output wire [127:0] io_connSS_8_data_availableTask_bits;
	output wire io_connSS_8_data_qOutTask_ready;
	input io_connSS_8_data_qOutTask_valid;
	input [127:0] io_connSS_8_data_qOutTask_bits;
	input io_connSS_9_ctrl_serveStealReq_valid;
	output wire io_connSS_9_ctrl_serveStealReq_ready;
	input io_connSS_9_ctrl_stealReq_valid;
	output wire io_connSS_9_ctrl_stealReq_ready;
	input io_connSS_9_data_availableTask_ready;
	output wire io_connSS_9_data_availableTask_valid;
	output wire [127:0] io_connSS_9_data_availableTask_bits;
	output wire io_connSS_9_data_qOutTask_ready;
	input io_connSS_9_data_qOutTask_valid;
	input [127:0] io_connSS_9_data_qOutTask_bits;
	input io_connSS_10_ctrl_serveStealReq_valid;
	output wire io_connSS_10_ctrl_serveStealReq_ready;
	input io_connSS_10_ctrl_stealReq_valid;
	output wire io_connSS_10_ctrl_stealReq_ready;
	input io_connSS_10_data_availableTask_ready;
	output wire io_connSS_10_data_availableTask_valid;
	output wire [127:0] io_connSS_10_data_availableTask_bits;
	output wire io_connSS_10_data_qOutTask_ready;
	input io_connSS_10_data_qOutTask_valid;
	input [127:0] io_connSS_10_data_qOutTask_bits;
	input io_connSS_11_ctrl_serveStealReq_valid;
	output wire io_connSS_11_ctrl_serveStealReq_ready;
	input io_connSS_11_ctrl_stealReq_valid;
	output wire io_connSS_11_ctrl_stealReq_ready;
	input io_connSS_11_data_availableTask_ready;
	output wire io_connSS_11_data_availableTask_valid;
	output wire [127:0] io_connSS_11_data_availableTask_bits;
	output wire io_connSS_11_data_qOutTask_ready;
	input io_connSS_11_data_qOutTask_valid;
	input [127:0] io_connSS_11_data_qOutTask_bits;
	input io_connSS_12_ctrl_serveStealReq_valid;
	output wire io_connSS_12_ctrl_serveStealReq_ready;
	input io_connSS_12_ctrl_stealReq_valid;
	output wire io_connSS_12_ctrl_stealReq_ready;
	input io_connSS_12_data_availableTask_ready;
	output wire io_connSS_12_data_availableTask_valid;
	output wire [127:0] io_connSS_12_data_availableTask_bits;
	output wire io_connSS_12_data_qOutTask_ready;
	input io_connSS_12_data_qOutTask_valid;
	input [127:0] io_connSS_12_data_qOutTask_bits;
	input io_connSS_13_ctrl_serveStealReq_valid;
	output wire io_connSS_13_ctrl_serveStealReq_ready;
	input io_connSS_13_ctrl_stealReq_valid;
	output wire io_connSS_13_ctrl_stealReq_ready;
	input io_connSS_13_data_availableTask_ready;
	output wire io_connSS_13_data_availableTask_valid;
	output wire [127:0] io_connSS_13_data_availableTask_bits;
	output wire io_connSS_13_data_qOutTask_ready;
	input io_connSS_13_data_qOutTask_valid;
	input [127:0] io_connSS_13_data_qOutTask_bits;
	input io_connSS_14_ctrl_serveStealReq_valid;
	output wire io_connSS_14_ctrl_serveStealReq_ready;
	input io_connSS_14_ctrl_stealReq_valid;
	output wire io_connSS_14_ctrl_stealReq_ready;
	input io_connSS_14_data_availableTask_ready;
	output wire io_connSS_14_data_availableTask_valid;
	output wire [127:0] io_connSS_14_data_availableTask_bits;
	output wire io_connSS_14_data_qOutTask_ready;
	input io_connSS_14_data_qOutTask_valid;
	input [127:0] io_connSS_14_data_qOutTask_bits;
	input io_connSS_15_ctrl_serveStealReq_valid;
	output wire io_connSS_15_ctrl_serveStealReq_ready;
	input io_connSS_15_ctrl_stealReq_valid;
	output wire io_connSS_15_ctrl_stealReq_ready;
	input io_connSS_15_data_availableTask_ready;
	output wire io_connSS_15_data_availableTask_valid;
	output wire [127:0] io_connSS_15_data_availableTask_bits;
	output wire io_connSS_15_data_qOutTask_ready;
	input io_connSS_15_data_qOutTask_valid;
	input [127:0] io_connSS_15_data_qOutTask_bits;
	input io_connSS_16_ctrl_serveStealReq_valid;
	output wire io_connSS_16_ctrl_serveStealReq_ready;
	input io_connSS_16_ctrl_stealReq_valid;
	output wire io_connSS_16_ctrl_stealReq_ready;
	input io_connSS_16_data_availableTask_ready;
	output wire io_connSS_16_data_availableTask_valid;
	output wire [127:0] io_connSS_16_data_availableTask_bits;
	output wire io_connSS_16_data_qOutTask_ready;
	input io_connSS_16_data_qOutTask_valid;
	input [127:0] io_connSS_16_data_qOutTask_bits;
	input io_connSS_17_ctrl_serveStealReq_valid;
	output wire io_connSS_17_ctrl_serveStealReq_ready;
	input io_connSS_17_ctrl_stealReq_valid;
	output wire io_connSS_17_ctrl_stealReq_ready;
	input io_connSS_17_data_availableTask_ready;
	output wire io_connSS_17_data_availableTask_valid;
	output wire [127:0] io_connSS_17_data_availableTask_bits;
	output wire io_connSS_17_data_qOutTask_ready;
	input io_connSS_17_data_qOutTask_valid;
	input [127:0] io_connSS_17_data_qOutTask_bits;
	input io_connSS_18_ctrl_serveStealReq_valid;
	output wire io_connSS_18_ctrl_serveStealReq_ready;
	input io_connSS_18_ctrl_stealReq_valid;
	output wire io_connSS_18_ctrl_stealReq_ready;
	input io_connSS_18_data_availableTask_ready;
	output wire io_connSS_18_data_availableTask_valid;
	output wire [127:0] io_connSS_18_data_availableTask_bits;
	output wire io_connSS_18_data_qOutTask_ready;
	input io_connSS_18_data_qOutTask_valid;
	input [127:0] io_connSS_18_data_qOutTask_bits;
	input io_connSS_19_ctrl_serveStealReq_valid;
	output wire io_connSS_19_ctrl_serveStealReq_ready;
	input io_connSS_19_ctrl_stealReq_valid;
	output wire io_connSS_19_ctrl_stealReq_ready;
	input io_connSS_19_data_availableTask_ready;
	output wire io_connSS_19_data_availableTask_valid;
	output wire [127:0] io_connSS_19_data_availableTask_bits;
	output wire io_connSS_19_data_qOutTask_ready;
	input io_connSS_19_data_qOutTask_valid;
	input [127:0] io_connSS_19_data_qOutTask_bits;
	input io_connSS_20_ctrl_serveStealReq_valid;
	output wire io_connSS_20_ctrl_serveStealReq_ready;
	input io_connSS_20_ctrl_stealReq_valid;
	output wire io_connSS_20_ctrl_stealReq_ready;
	input io_connSS_20_data_availableTask_ready;
	output wire io_connSS_20_data_availableTask_valid;
	output wire [127:0] io_connSS_20_data_availableTask_bits;
	output wire io_connSS_20_data_qOutTask_ready;
	input io_connSS_20_data_qOutTask_valid;
	input [127:0] io_connSS_20_data_qOutTask_bits;
	input io_connSS_21_ctrl_serveStealReq_valid;
	output wire io_connSS_21_ctrl_serveStealReq_ready;
	input io_connSS_21_ctrl_stealReq_valid;
	output wire io_connSS_21_ctrl_stealReq_ready;
	input io_connSS_21_data_availableTask_ready;
	output wire io_connSS_21_data_availableTask_valid;
	output wire [127:0] io_connSS_21_data_availableTask_bits;
	output wire io_connSS_21_data_qOutTask_ready;
	input io_connSS_21_data_qOutTask_valid;
	input [127:0] io_connSS_21_data_qOutTask_bits;
	input io_connSS_22_ctrl_serveStealReq_valid;
	output wire io_connSS_22_ctrl_serveStealReq_ready;
	input io_connSS_22_ctrl_stealReq_valid;
	output wire io_connSS_22_ctrl_stealReq_ready;
	input io_connSS_22_data_availableTask_ready;
	output wire io_connSS_22_data_availableTask_valid;
	output wire [127:0] io_connSS_22_data_availableTask_bits;
	output wire io_connSS_22_data_qOutTask_ready;
	input io_connSS_22_data_qOutTask_valid;
	input [127:0] io_connSS_22_data_qOutTask_bits;
	input io_connSS_23_ctrl_serveStealReq_valid;
	output wire io_connSS_23_ctrl_serveStealReq_ready;
	input io_connSS_23_ctrl_stealReq_valid;
	output wire io_connSS_23_ctrl_stealReq_ready;
	input io_connSS_23_data_availableTask_ready;
	output wire io_connSS_23_data_availableTask_valid;
	output wire [127:0] io_connSS_23_data_availableTask_bits;
	output wire io_connSS_23_data_qOutTask_ready;
	input io_connSS_23_data_qOutTask_valid;
	input [127:0] io_connSS_23_data_qOutTask_bits;
	input io_connSS_24_ctrl_serveStealReq_valid;
	output wire io_connSS_24_ctrl_serveStealReq_ready;
	input io_connSS_24_ctrl_stealReq_valid;
	output wire io_connSS_24_ctrl_stealReq_ready;
	input io_connSS_24_data_availableTask_ready;
	output wire io_connSS_24_data_availableTask_valid;
	output wire [127:0] io_connSS_24_data_availableTask_bits;
	output wire io_connSS_24_data_qOutTask_ready;
	input io_connSS_24_data_qOutTask_valid;
	input [127:0] io_connSS_24_data_qOutTask_bits;
	input io_connSS_25_ctrl_serveStealReq_valid;
	output wire io_connSS_25_ctrl_serveStealReq_ready;
	input io_connSS_25_ctrl_stealReq_valid;
	output wire io_connSS_25_ctrl_stealReq_ready;
	input io_connSS_25_data_availableTask_ready;
	output wire io_connSS_25_data_availableTask_valid;
	output wire [127:0] io_connSS_25_data_availableTask_bits;
	output wire io_connSS_25_data_qOutTask_ready;
	input io_connSS_25_data_qOutTask_valid;
	input [127:0] io_connSS_25_data_qOutTask_bits;
	input io_connSS_26_ctrl_serveStealReq_valid;
	output wire io_connSS_26_ctrl_serveStealReq_ready;
	input io_connSS_26_ctrl_stealReq_valid;
	output wire io_connSS_26_ctrl_stealReq_ready;
	input io_connSS_26_data_availableTask_ready;
	output wire io_connSS_26_data_availableTask_valid;
	output wire [127:0] io_connSS_26_data_availableTask_bits;
	output wire io_connSS_26_data_qOutTask_ready;
	input io_connSS_26_data_qOutTask_valid;
	input [127:0] io_connSS_26_data_qOutTask_bits;
	input io_connSS_27_ctrl_serveStealReq_valid;
	output wire io_connSS_27_ctrl_serveStealReq_ready;
	input io_connSS_27_ctrl_stealReq_valid;
	output wire io_connSS_27_ctrl_stealReq_ready;
	input io_connSS_27_data_availableTask_ready;
	output wire io_connSS_27_data_availableTask_valid;
	output wire [127:0] io_connSS_27_data_availableTask_bits;
	output wire io_connSS_27_data_qOutTask_ready;
	input io_connSS_27_data_qOutTask_valid;
	input [127:0] io_connSS_27_data_qOutTask_bits;
	input io_connSS_28_ctrl_serveStealReq_valid;
	output wire io_connSS_28_ctrl_serveStealReq_ready;
	input io_connSS_28_ctrl_stealReq_valid;
	output wire io_connSS_28_ctrl_stealReq_ready;
	input io_connSS_28_data_availableTask_ready;
	output wire io_connSS_28_data_availableTask_valid;
	output wire [127:0] io_connSS_28_data_availableTask_bits;
	output wire io_connSS_28_data_qOutTask_ready;
	input io_connSS_28_data_qOutTask_valid;
	input [127:0] io_connSS_28_data_qOutTask_bits;
	input io_connSS_29_ctrl_serveStealReq_valid;
	output wire io_connSS_29_ctrl_serveStealReq_ready;
	input io_connSS_29_ctrl_stealReq_valid;
	output wire io_connSS_29_ctrl_stealReq_ready;
	input io_connSS_29_data_availableTask_ready;
	output wire io_connSS_29_data_availableTask_valid;
	output wire [127:0] io_connSS_29_data_availableTask_bits;
	output wire io_connSS_29_data_qOutTask_ready;
	input io_connSS_29_data_qOutTask_valid;
	input [127:0] io_connSS_29_data_qOutTask_bits;
	input io_connSS_30_ctrl_serveStealReq_valid;
	output wire io_connSS_30_ctrl_serveStealReq_ready;
	input io_connSS_30_ctrl_stealReq_valid;
	output wire io_connSS_30_ctrl_stealReq_ready;
	input io_connSS_30_data_availableTask_ready;
	output wire io_connSS_30_data_availableTask_valid;
	output wire [127:0] io_connSS_30_data_availableTask_bits;
	output wire io_connSS_30_data_qOutTask_ready;
	input io_connSS_30_data_qOutTask_valid;
	input [127:0] io_connSS_30_data_qOutTask_bits;
	input io_connSS_31_ctrl_serveStealReq_valid;
	output wire io_connSS_31_ctrl_serveStealReq_ready;
	input io_connSS_31_ctrl_stealReq_valid;
	output wire io_connSS_31_ctrl_stealReq_ready;
	input io_connSS_31_data_availableTask_ready;
	output wire io_connSS_31_data_availableTask_valid;
	output wire [127:0] io_connSS_31_data_availableTask_bits;
	output wire io_connSS_31_data_qOutTask_ready;
	input io_connSS_31_data_qOutTask_valid;
	input [127:0] io_connSS_31_data_qOutTask_bits;
	input io_connSS_32_ctrl_serveStealReq_valid;
	output wire io_connSS_32_ctrl_serveStealReq_ready;
	input io_connSS_32_ctrl_stealReq_valid;
	output wire io_connSS_32_ctrl_stealReq_ready;
	input io_connSS_32_data_availableTask_ready;
	output wire io_connSS_32_data_availableTask_valid;
	output wire [127:0] io_connSS_32_data_availableTask_bits;
	output wire io_connSS_32_data_qOutTask_ready;
	input io_connSS_32_data_qOutTask_valid;
	input [127:0] io_connSS_32_data_qOutTask_bits;
	input io_connSS_33_ctrl_serveStealReq_valid;
	output wire io_connSS_33_ctrl_serveStealReq_ready;
	input io_connSS_33_data_availableTask_ready;
	output wire io_connSS_33_data_availableTask_valid;
	output wire [127:0] io_connSS_33_data_availableTask_bits;
	output wire io_connSS_33_data_qOutTask_ready;
	input io_connSS_33_data_qOutTask_valid;
	input [127:0] io_connSS_33_data_qOutTask_bits;
	input io_connSS_34_ctrl_serveStealReq_valid;
	output wire io_connSS_34_ctrl_serveStealReq_ready;
	input io_connSS_34_ctrl_stealReq_valid;
	output wire io_connSS_34_ctrl_stealReq_ready;
	input io_connSS_34_data_availableTask_ready;
	output wire io_connSS_34_data_availableTask_valid;
	output wire [127:0] io_connSS_34_data_availableTask_bits;
	output wire io_connSS_34_data_qOutTask_ready;
	input io_connSS_34_data_qOutTask_valid;
	input [127:0] io_connSS_34_data_qOutTask_bits;
	input io_connSS_35_ctrl_serveStealReq_valid;
	output wire io_connSS_35_ctrl_serveStealReq_ready;
	input io_connSS_35_ctrl_stealReq_valid;
	output wire io_connSS_35_ctrl_stealReq_ready;
	input io_connSS_35_data_availableTask_ready;
	output wire io_connSS_35_data_availableTask_valid;
	output wire [127:0] io_connSS_35_data_availableTask_bits;
	output wire io_connSS_35_data_qOutTask_ready;
	input io_connSS_35_data_qOutTask_valid;
	input [127:0] io_connSS_35_data_qOutTask_bits;
	input io_connSS_36_ctrl_serveStealReq_valid;
	output wire io_connSS_36_ctrl_serveStealReq_ready;
	input io_connSS_36_ctrl_stealReq_valid;
	output wire io_connSS_36_ctrl_stealReq_ready;
	input io_connSS_36_data_availableTask_ready;
	output wire io_connSS_36_data_availableTask_valid;
	output wire [127:0] io_connSS_36_data_availableTask_bits;
	output wire io_connSS_36_data_qOutTask_ready;
	input io_connSS_36_data_qOutTask_valid;
	input [127:0] io_connSS_36_data_qOutTask_bits;
	input io_connSS_37_ctrl_serveStealReq_valid;
	output wire io_connSS_37_ctrl_serveStealReq_ready;
	input io_connSS_37_ctrl_stealReq_valid;
	output wire io_connSS_37_ctrl_stealReq_ready;
	input io_connSS_37_data_availableTask_ready;
	output wire io_connSS_37_data_availableTask_valid;
	output wire [127:0] io_connSS_37_data_availableTask_bits;
	output wire io_connSS_37_data_qOutTask_ready;
	input io_connSS_37_data_qOutTask_valid;
	input [127:0] io_connSS_37_data_qOutTask_bits;
	input io_connSS_38_ctrl_serveStealReq_valid;
	output wire io_connSS_38_ctrl_serveStealReq_ready;
	input io_connSS_38_ctrl_stealReq_valid;
	output wire io_connSS_38_ctrl_stealReq_ready;
	input io_connSS_38_data_availableTask_ready;
	output wire io_connSS_38_data_availableTask_valid;
	output wire [127:0] io_connSS_38_data_availableTask_bits;
	output wire io_connSS_38_data_qOutTask_ready;
	input io_connSS_38_data_qOutTask_valid;
	input [127:0] io_connSS_38_data_qOutTask_bits;
	input io_connSS_39_ctrl_serveStealReq_valid;
	output wire io_connSS_39_ctrl_serveStealReq_ready;
	input io_connSS_39_ctrl_stealReq_valid;
	output wire io_connSS_39_ctrl_stealReq_ready;
	input io_connSS_39_data_availableTask_ready;
	output wire io_connSS_39_data_availableTask_valid;
	output wire [127:0] io_connSS_39_data_availableTask_bits;
	output wire io_connSS_39_data_qOutTask_ready;
	input io_connSS_39_data_qOutTask_valid;
	input [127:0] io_connSS_39_data_qOutTask_bits;
	input io_connSS_40_ctrl_serveStealReq_valid;
	output wire io_connSS_40_ctrl_serveStealReq_ready;
	input io_connSS_40_ctrl_stealReq_valid;
	output wire io_connSS_40_ctrl_stealReq_ready;
	input io_connSS_40_data_availableTask_ready;
	output wire io_connSS_40_data_availableTask_valid;
	output wire [127:0] io_connSS_40_data_availableTask_bits;
	output wire io_connSS_40_data_qOutTask_ready;
	input io_connSS_40_data_qOutTask_valid;
	input [127:0] io_connSS_40_data_qOutTask_bits;
	input io_connSS_41_ctrl_serveStealReq_valid;
	output wire io_connSS_41_ctrl_serveStealReq_ready;
	input io_connSS_41_ctrl_stealReq_valid;
	output wire io_connSS_41_ctrl_stealReq_ready;
	input io_connSS_41_data_availableTask_ready;
	output wire io_connSS_41_data_availableTask_valid;
	output wire [127:0] io_connSS_41_data_availableTask_bits;
	output wire io_connSS_41_data_qOutTask_ready;
	input io_connSS_41_data_qOutTask_valid;
	input [127:0] io_connSS_41_data_qOutTask_bits;
	input io_connSS_42_ctrl_serveStealReq_valid;
	output wire io_connSS_42_ctrl_serveStealReq_ready;
	input io_connSS_42_ctrl_stealReq_valid;
	output wire io_connSS_42_ctrl_stealReq_ready;
	input io_connSS_42_data_availableTask_ready;
	output wire io_connSS_42_data_availableTask_valid;
	output wire [127:0] io_connSS_42_data_availableTask_bits;
	output wire io_connSS_42_data_qOutTask_ready;
	input io_connSS_42_data_qOutTask_valid;
	input [127:0] io_connSS_42_data_qOutTask_bits;
	input io_connSS_43_ctrl_serveStealReq_valid;
	output wire io_connSS_43_ctrl_serveStealReq_ready;
	input io_connSS_43_ctrl_stealReq_valid;
	output wire io_connSS_43_ctrl_stealReq_ready;
	input io_connSS_43_data_availableTask_ready;
	output wire io_connSS_43_data_availableTask_valid;
	output wire [127:0] io_connSS_43_data_availableTask_bits;
	output wire io_connSS_43_data_qOutTask_ready;
	input io_connSS_43_data_qOutTask_valid;
	input [127:0] io_connSS_43_data_qOutTask_bits;
	input io_connSS_44_ctrl_serveStealReq_valid;
	output wire io_connSS_44_ctrl_serveStealReq_ready;
	input io_connSS_44_ctrl_stealReq_valid;
	output wire io_connSS_44_ctrl_stealReq_ready;
	input io_connSS_44_data_availableTask_ready;
	output wire io_connSS_44_data_availableTask_valid;
	output wire [127:0] io_connSS_44_data_availableTask_bits;
	output wire io_connSS_44_data_qOutTask_ready;
	input io_connSS_44_data_qOutTask_valid;
	input [127:0] io_connSS_44_data_qOutTask_bits;
	input io_connSS_45_ctrl_serveStealReq_valid;
	output wire io_connSS_45_ctrl_serveStealReq_ready;
	input io_connSS_45_ctrl_stealReq_valid;
	output wire io_connSS_45_ctrl_stealReq_ready;
	input io_connSS_45_data_availableTask_ready;
	output wire io_connSS_45_data_availableTask_valid;
	output wire [127:0] io_connSS_45_data_availableTask_bits;
	output wire io_connSS_45_data_qOutTask_ready;
	input io_connSS_45_data_qOutTask_valid;
	input [127:0] io_connSS_45_data_qOutTask_bits;
	input io_connSS_46_ctrl_serveStealReq_valid;
	output wire io_connSS_46_ctrl_serveStealReq_ready;
	input io_connSS_46_ctrl_stealReq_valid;
	output wire io_connSS_46_ctrl_stealReq_ready;
	input io_connSS_46_data_availableTask_ready;
	output wire io_connSS_46_data_availableTask_valid;
	output wire [127:0] io_connSS_46_data_availableTask_bits;
	output wire io_connSS_46_data_qOutTask_ready;
	input io_connSS_46_data_qOutTask_valid;
	input [127:0] io_connSS_46_data_qOutTask_bits;
	input io_connSS_47_ctrl_serveStealReq_valid;
	output wire io_connSS_47_ctrl_serveStealReq_ready;
	input io_connSS_47_ctrl_stealReq_valid;
	output wire io_connSS_47_ctrl_stealReq_ready;
	input io_connSS_47_data_availableTask_ready;
	output wire io_connSS_47_data_availableTask_valid;
	output wire [127:0] io_connSS_47_data_availableTask_bits;
	output wire io_connSS_47_data_qOutTask_ready;
	input io_connSS_47_data_qOutTask_valid;
	input [127:0] io_connSS_47_data_qOutTask_bits;
	input io_connSS_48_ctrl_serveStealReq_valid;
	output wire io_connSS_48_ctrl_serveStealReq_ready;
	input io_connSS_48_ctrl_stealReq_valid;
	output wire io_connSS_48_ctrl_stealReq_ready;
	input io_connSS_48_data_availableTask_ready;
	output wire io_connSS_48_data_availableTask_valid;
	output wire [127:0] io_connSS_48_data_availableTask_bits;
	output wire io_connSS_48_data_qOutTask_ready;
	input io_connSS_48_data_qOutTask_valid;
	input [127:0] io_connSS_48_data_qOutTask_bits;
	input io_connSS_49_ctrl_serveStealReq_valid;
	output wire io_connSS_49_ctrl_serveStealReq_ready;
	input io_connSS_49_ctrl_stealReq_valid;
	output wire io_connSS_49_ctrl_stealReq_ready;
	input io_connSS_49_data_availableTask_ready;
	output wire io_connSS_49_data_availableTask_valid;
	output wire [127:0] io_connSS_49_data_availableTask_bits;
	output wire io_connSS_49_data_qOutTask_ready;
	input io_connSS_49_data_qOutTask_valid;
	input [127:0] io_connSS_49_data_qOutTask_bits;
	input io_connSS_50_ctrl_serveStealReq_valid;
	output wire io_connSS_50_ctrl_serveStealReq_ready;
	input io_connSS_50_ctrl_stealReq_valid;
	output wire io_connSS_50_ctrl_stealReq_ready;
	input io_connSS_50_data_availableTask_ready;
	output wire io_connSS_50_data_availableTask_valid;
	output wire [127:0] io_connSS_50_data_availableTask_bits;
	output wire io_connSS_50_data_qOutTask_ready;
	input io_connSS_50_data_qOutTask_valid;
	input [127:0] io_connSS_50_data_qOutTask_bits;
	input io_connSS_51_ctrl_serveStealReq_valid;
	output wire io_connSS_51_ctrl_serveStealReq_ready;
	input io_connSS_51_ctrl_stealReq_valid;
	output wire io_connSS_51_ctrl_stealReq_ready;
	input io_connSS_51_data_availableTask_ready;
	output wire io_connSS_51_data_availableTask_valid;
	output wire [127:0] io_connSS_51_data_availableTask_bits;
	output wire io_connSS_51_data_qOutTask_ready;
	input io_connSS_51_data_qOutTask_valid;
	input [127:0] io_connSS_51_data_qOutTask_bits;
	input io_connSS_52_ctrl_serveStealReq_valid;
	output wire io_connSS_52_ctrl_serveStealReq_ready;
	input io_connSS_52_ctrl_stealReq_valid;
	output wire io_connSS_52_ctrl_stealReq_ready;
	input io_connSS_52_data_availableTask_ready;
	output wire io_connSS_52_data_availableTask_valid;
	output wire [127:0] io_connSS_52_data_availableTask_bits;
	output wire io_connSS_52_data_qOutTask_ready;
	input io_connSS_52_data_qOutTask_valid;
	input [127:0] io_connSS_52_data_qOutTask_bits;
	input io_connSS_53_ctrl_serveStealReq_valid;
	output wire io_connSS_53_ctrl_serveStealReq_ready;
	input io_connSS_53_ctrl_stealReq_valid;
	output wire io_connSS_53_ctrl_stealReq_ready;
	input io_connSS_53_data_availableTask_ready;
	output wire io_connSS_53_data_availableTask_valid;
	output wire [127:0] io_connSS_53_data_availableTask_bits;
	output wire io_connSS_53_data_qOutTask_ready;
	input io_connSS_53_data_qOutTask_valid;
	input [127:0] io_connSS_53_data_qOutTask_bits;
	input io_connSS_54_ctrl_serveStealReq_valid;
	output wire io_connSS_54_ctrl_serveStealReq_ready;
	input io_connSS_54_ctrl_stealReq_valid;
	output wire io_connSS_54_ctrl_stealReq_ready;
	input io_connSS_54_data_availableTask_ready;
	output wire io_connSS_54_data_availableTask_valid;
	output wire [127:0] io_connSS_54_data_availableTask_bits;
	output wire io_connSS_54_data_qOutTask_ready;
	input io_connSS_54_data_qOutTask_valid;
	input [127:0] io_connSS_54_data_qOutTask_bits;
	input io_connSS_55_ctrl_serveStealReq_valid;
	output wire io_connSS_55_ctrl_serveStealReq_ready;
	input io_connSS_55_ctrl_stealReq_valid;
	output wire io_connSS_55_ctrl_stealReq_ready;
	input io_connSS_55_data_availableTask_ready;
	output wire io_connSS_55_data_availableTask_valid;
	output wire [127:0] io_connSS_55_data_availableTask_bits;
	output wire io_connSS_55_data_qOutTask_ready;
	input io_connSS_55_data_qOutTask_valid;
	input [127:0] io_connSS_55_data_qOutTask_bits;
	input io_connSS_56_ctrl_serveStealReq_valid;
	output wire io_connSS_56_ctrl_serveStealReq_ready;
	input io_connSS_56_ctrl_stealReq_valid;
	output wire io_connSS_56_ctrl_stealReq_ready;
	input io_connSS_56_data_availableTask_ready;
	output wire io_connSS_56_data_availableTask_valid;
	output wire [127:0] io_connSS_56_data_availableTask_bits;
	output wire io_connSS_56_data_qOutTask_ready;
	input io_connSS_56_data_qOutTask_valid;
	input [127:0] io_connSS_56_data_qOutTask_bits;
	input io_connSS_57_ctrl_serveStealReq_valid;
	output wire io_connSS_57_ctrl_serveStealReq_ready;
	input io_connSS_57_ctrl_stealReq_valid;
	output wire io_connSS_57_ctrl_stealReq_ready;
	input io_connSS_57_data_availableTask_ready;
	output wire io_connSS_57_data_availableTask_valid;
	output wire [127:0] io_connSS_57_data_availableTask_bits;
	output wire io_connSS_57_data_qOutTask_ready;
	input io_connSS_57_data_qOutTask_valid;
	input [127:0] io_connSS_57_data_qOutTask_bits;
	input io_connSS_58_ctrl_serveStealReq_valid;
	output wire io_connSS_58_ctrl_serveStealReq_ready;
	input io_connSS_58_ctrl_stealReq_valid;
	output wire io_connSS_58_ctrl_stealReq_ready;
	input io_connSS_58_data_availableTask_ready;
	output wire io_connSS_58_data_availableTask_valid;
	output wire [127:0] io_connSS_58_data_availableTask_bits;
	output wire io_connSS_58_data_qOutTask_ready;
	input io_connSS_58_data_qOutTask_valid;
	input [127:0] io_connSS_58_data_qOutTask_bits;
	input io_connSS_59_ctrl_serveStealReq_valid;
	output wire io_connSS_59_ctrl_serveStealReq_ready;
	input io_connSS_59_ctrl_stealReq_valid;
	output wire io_connSS_59_ctrl_stealReq_ready;
	input io_connSS_59_data_availableTask_ready;
	output wire io_connSS_59_data_availableTask_valid;
	output wire [127:0] io_connSS_59_data_availableTask_bits;
	output wire io_connSS_59_data_qOutTask_ready;
	input io_connSS_59_data_qOutTask_valid;
	input [127:0] io_connSS_59_data_qOutTask_bits;
	input io_connSS_60_ctrl_serveStealReq_valid;
	output wire io_connSS_60_ctrl_serveStealReq_ready;
	input io_connSS_60_ctrl_stealReq_valid;
	output wire io_connSS_60_ctrl_stealReq_ready;
	input io_connSS_60_data_availableTask_ready;
	output wire io_connSS_60_data_availableTask_valid;
	output wire [127:0] io_connSS_60_data_availableTask_bits;
	output wire io_connSS_60_data_qOutTask_ready;
	input io_connSS_60_data_qOutTask_valid;
	input [127:0] io_connSS_60_data_qOutTask_bits;
	input io_connSS_61_ctrl_serveStealReq_valid;
	output wire io_connSS_61_ctrl_serveStealReq_ready;
	input io_connSS_61_ctrl_stealReq_valid;
	output wire io_connSS_61_ctrl_stealReq_ready;
	input io_connSS_61_data_availableTask_ready;
	output wire io_connSS_61_data_availableTask_valid;
	output wire [127:0] io_connSS_61_data_availableTask_bits;
	output wire io_connSS_61_data_qOutTask_ready;
	input io_connSS_61_data_qOutTask_valid;
	input [127:0] io_connSS_61_data_qOutTask_bits;
	input io_connSS_62_ctrl_serveStealReq_valid;
	output wire io_connSS_62_ctrl_serveStealReq_ready;
	input io_connSS_62_ctrl_stealReq_valid;
	output wire io_connSS_62_ctrl_stealReq_ready;
	input io_connSS_62_data_availableTask_ready;
	output wire io_connSS_62_data_availableTask_valid;
	output wire [127:0] io_connSS_62_data_availableTask_bits;
	output wire io_connSS_62_data_qOutTask_ready;
	input io_connSS_62_data_qOutTask_valid;
	input [127:0] io_connSS_62_data_qOutTask_bits;
	input io_connSS_63_ctrl_serveStealReq_valid;
	output wire io_connSS_63_ctrl_serveStealReq_ready;
	input io_connSS_63_ctrl_stealReq_valid;
	output wire io_connSS_63_ctrl_stealReq_ready;
	input io_connSS_63_data_availableTask_ready;
	output wire io_connSS_63_data_availableTask_valid;
	output wire [127:0] io_connSS_63_data_availableTask_bits;
	output wire io_connSS_63_data_qOutTask_ready;
	input io_connSS_63_data_qOutTask_valid;
	input [127:0] io_connSS_63_data_qOutTask_bits;
	input io_connSS_64_ctrl_serveStealReq_valid;
	output wire io_connSS_64_ctrl_serveStealReq_ready;
	input io_connSS_64_ctrl_stealReq_valid;
	output wire io_connSS_64_ctrl_stealReq_ready;
	input io_connSS_64_data_availableTask_ready;
	output wire io_connSS_64_data_availableTask_valid;
	output wire [127:0] io_connSS_64_data_availableTask_bits;
	output wire io_connSS_64_data_qOutTask_ready;
	input io_connSS_64_data_qOutTask_valid;
	input [127:0] io_connSS_64_data_qOutTask_bits;
	input io_connSS_65_ctrl_serveStealReq_valid;
	output wire io_connSS_65_ctrl_serveStealReq_ready;
	input io_connSS_65_ctrl_stealReq_valid;
	output wire io_connSS_65_ctrl_stealReq_ready;
	input io_connSS_65_data_availableTask_ready;
	output wire io_connSS_65_data_availableTask_valid;
	output wire [127:0] io_connSS_65_data_availableTask_bits;
	output wire io_connSS_65_data_qOutTask_ready;
	input io_connSS_65_data_qOutTask_valid;
	input [127:0] io_connSS_65_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	output wire io_ntwDataUnitOccupancyVSS_1;
	wire _ctrlunits_65_io_reqTaskOut;
	wire _ctrlunits_64_io_reqTaskOut;
	wire _ctrlunits_63_io_reqTaskOut;
	wire _ctrlunits_62_io_reqTaskOut;
	wire _ctrlunits_61_io_reqTaskOut;
	wire _ctrlunits_60_io_reqTaskOut;
	wire _ctrlunits_59_io_reqTaskOut;
	wire _ctrlunits_58_io_reqTaskOut;
	wire _ctrlunits_57_io_reqTaskOut;
	wire _ctrlunits_56_io_reqTaskOut;
	wire _ctrlunits_55_io_reqTaskOut;
	wire _ctrlunits_54_io_reqTaskOut;
	wire _ctrlunits_53_io_reqTaskOut;
	wire _ctrlunits_52_io_reqTaskOut;
	wire _ctrlunits_51_io_reqTaskOut;
	wire _ctrlunits_50_io_reqTaskOut;
	wire _ctrlunits_49_io_reqTaskOut;
	wire _ctrlunits_48_io_reqTaskOut;
	wire _ctrlunits_47_io_reqTaskOut;
	wire _ctrlunits_46_io_reqTaskOut;
	wire _ctrlunits_45_io_reqTaskOut;
	wire _ctrlunits_44_io_reqTaskOut;
	wire _ctrlunits_43_io_reqTaskOut;
	wire _ctrlunits_42_io_reqTaskOut;
	wire _ctrlunits_41_io_reqTaskOut;
	wire _ctrlunits_40_io_reqTaskOut;
	wire _ctrlunits_39_io_reqTaskOut;
	wire _ctrlunits_38_io_reqTaskOut;
	wire _ctrlunits_37_io_reqTaskOut;
	wire _ctrlunits_36_io_reqTaskOut;
	wire _ctrlunits_35_io_reqTaskOut;
	wire _ctrlunits_34_io_reqTaskOut;
	wire _ctrlunits_33_io_reqTaskOut;
	wire _ctrlunits_32_io_reqTaskOut;
	wire _ctrlunits_31_io_reqTaskOut;
	wire _ctrlunits_30_io_reqTaskOut;
	wire _ctrlunits_29_io_reqTaskOut;
	wire _ctrlunits_28_io_reqTaskOut;
	wire _ctrlunits_27_io_reqTaskOut;
	wire _ctrlunits_26_io_reqTaskOut;
	wire _ctrlunits_25_io_reqTaskOut;
	wire _ctrlunits_24_io_reqTaskOut;
	wire _ctrlunits_23_io_reqTaskOut;
	wire _ctrlunits_22_io_reqTaskOut;
	wire _ctrlunits_21_io_reqTaskOut;
	wire _ctrlunits_20_io_reqTaskOut;
	wire _ctrlunits_19_io_reqTaskOut;
	wire _ctrlunits_18_io_reqTaskOut;
	wire _ctrlunits_17_io_reqTaskOut;
	wire _ctrlunits_16_io_reqTaskOut;
	wire _ctrlunits_15_io_reqTaskOut;
	wire _ctrlunits_14_io_reqTaskOut;
	wire _ctrlunits_13_io_reqTaskOut;
	wire _ctrlunits_12_io_reqTaskOut;
	wire _ctrlunits_11_io_reqTaskOut;
	wire _ctrlunits_10_io_reqTaskOut;
	wire _ctrlunits_9_io_reqTaskOut;
	wire _ctrlunits_8_io_reqTaskOut;
	wire _ctrlunits_7_io_reqTaskOut;
	wire _ctrlunits_6_io_reqTaskOut;
	wire _ctrlunits_5_io_reqTaskOut;
	wire _ctrlunits_4_io_reqTaskOut;
	wire _ctrlunits_3_io_reqTaskOut;
	wire _ctrlunits_2_io_reqTaskOut;
	wire _ctrlunits_1_io_reqTaskOut;
	wire _ctrlunits_0_io_reqTaskOut;
	wire [127:0] _dataUnits_65_io_taskOut;
	wire _dataUnits_65_io_validOut;
	wire [127:0] _dataUnits_64_io_taskOut;
	wire _dataUnits_64_io_validOut;
	wire [127:0] _dataUnits_63_io_taskOut;
	wire _dataUnits_63_io_validOut;
	wire [127:0] _dataUnits_62_io_taskOut;
	wire _dataUnits_62_io_validOut;
	wire [127:0] _dataUnits_61_io_taskOut;
	wire _dataUnits_61_io_validOut;
	wire [127:0] _dataUnits_60_io_taskOut;
	wire _dataUnits_60_io_validOut;
	wire [127:0] _dataUnits_59_io_taskOut;
	wire _dataUnits_59_io_validOut;
	wire [127:0] _dataUnits_58_io_taskOut;
	wire _dataUnits_58_io_validOut;
	wire [127:0] _dataUnits_57_io_taskOut;
	wire _dataUnits_57_io_validOut;
	wire [127:0] _dataUnits_56_io_taskOut;
	wire _dataUnits_56_io_validOut;
	wire [127:0] _dataUnits_55_io_taskOut;
	wire _dataUnits_55_io_validOut;
	wire [127:0] _dataUnits_54_io_taskOut;
	wire _dataUnits_54_io_validOut;
	wire [127:0] _dataUnits_53_io_taskOut;
	wire _dataUnits_53_io_validOut;
	wire [127:0] _dataUnits_52_io_taskOut;
	wire _dataUnits_52_io_validOut;
	wire [127:0] _dataUnits_51_io_taskOut;
	wire _dataUnits_51_io_validOut;
	wire [127:0] _dataUnits_50_io_taskOut;
	wire _dataUnits_50_io_validOut;
	wire [127:0] _dataUnits_49_io_taskOut;
	wire _dataUnits_49_io_validOut;
	wire [127:0] _dataUnits_48_io_taskOut;
	wire _dataUnits_48_io_validOut;
	wire [127:0] _dataUnits_47_io_taskOut;
	wire _dataUnits_47_io_validOut;
	wire [127:0] _dataUnits_46_io_taskOut;
	wire _dataUnits_46_io_validOut;
	wire [127:0] _dataUnits_45_io_taskOut;
	wire _dataUnits_45_io_validOut;
	wire [127:0] _dataUnits_44_io_taskOut;
	wire _dataUnits_44_io_validOut;
	wire [127:0] _dataUnits_43_io_taskOut;
	wire _dataUnits_43_io_validOut;
	wire [127:0] _dataUnits_42_io_taskOut;
	wire _dataUnits_42_io_validOut;
	wire [127:0] _dataUnits_41_io_taskOut;
	wire _dataUnits_41_io_validOut;
	wire [127:0] _dataUnits_40_io_taskOut;
	wire _dataUnits_40_io_validOut;
	wire [127:0] _dataUnits_39_io_taskOut;
	wire _dataUnits_39_io_validOut;
	wire [127:0] _dataUnits_38_io_taskOut;
	wire _dataUnits_38_io_validOut;
	wire [127:0] _dataUnits_37_io_taskOut;
	wire _dataUnits_37_io_validOut;
	wire [127:0] _dataUnits_36_io_taskOut;
	wire _dataUnits_36_io_validOut;
	wire [127:0] _dataUnits_35_io_taskOut;
	wire _dataUnits_35_io_validOut;
	wire [127:0] _dataUnits_34_io_taskOut;
	wire _dataUnits_34_io_validOut;
	wire [127:0] _dataUnits_33_io_taskOut;
	wire _dataUnits_33_io_validOut;
	wire [127:0] _dataUnits_32_io_taskOut;
	wire _dataUnits_32_io_validOut;
	wire [127:0] _dataUnits_31_io_taskOut;
	wire _dataUnits_31_io_validOut;
	wire [127:0] _dataUnits_30_io_taskOut;
	wire _dataUnits_30_io_validOut;
	wire [127:0] _dataUnits_29_io_taskOut;
	wire _dataUnits_29_io_validOut;
	wire [127:0] _dataUnits_28_io_taskOut;
	wire _dataUnits_28_io_validOut;
	wire [127:0] _dataUnits_27_io_taskOut;
	wire _dataUnits_27_io_validOut;
	wire [127:0] _dataUnits_26_io_taskOut;
	wire _dataUnits_26_io_validOut;
	wire [127:0] _dataUnits_25_io_taskOut;
	wire _dataUnits_25_io_validOut;
	wire [127:0] _dataUnits_24_io_taskOut;
	wire _dataUnits_24_io_validOut;
	wire [127:0] _dataUnits_23_io_taskOut;
	wire _dataUnits_23_io_validOut;
	wire [127:0] _dataUnits_22_io_taskOut;
	wire _dataUnits_22_io_validOut;
	wire [127:0] _dataUnits_21_io_taskOut;
	wire _dataUnits_21_io_validOut;
	wire [127:0] _dataUnits_20_io_taskOut;
	wire _dataUnits_20_io_validOut;
	wire [127:0] _dataUnits_19_io_taskOut;
	wire _dataUnits_19_io_validOut;
	wire [127:0] _dataUnits_18_io_taskOut;
	wire _dataUnits_18_io_validOut;
	wire [127:0] _dataUnits_17_io_taskOut;
	wire _dataUnits_17_io_validOut;
	wire [127:0] _dataUnits_16_io_taskOut;
	wire _dataUnits_16_io_validOut;
	wire [127:0] _dataUnits_15_io_taskOut;
	wire _dataUnits_15_io_validOut;
	wire [127:0] _dataUnits_14_io_taskOut;
	wire _dataUnits_14_io_validOut;
	wire [127:0] _dataUnits_13_io_taskOut;
	wire _dataUnits_13_io_validOut;
	wire [127:0] _dataUnits_12_io_taskOut;
	wire _dataUnits_12_io_validOut;
	wire [127:0] _dataUnits_11_io_taskOut;
	wire _dataUnits_11_io_validOut;
	wire [127:0] _dataUnits_10_io_taskOut;
	wire _dataUnits_10_io_validOut;
	wire [127:0] _dataUnits_9_io_taskOut;
	wire _dataUnits_9_io_validOut;
	wire [127:0] _dataUnits_8_io_taskOut;
	wire _dataUnits_8_io_validOut;
	wire [127:0] _dataUnits_7_io_taskOut;
	wire _dataUnits_7_io_validOut;
	wire [127:0] _dataUnits_6_io_taskOut;
	wire _dataUnits_6_io_validOut;
	wire [127:0] _dataUnits_5_io_taskOut;
	wire _dataUnits_5_io_validOut;
	wire [127:0] _dataUnits_4_io_taskOut;
	wire _dataUnits_4_io_validOut;
	wire [127:0] _dataUnits_3_io_taskOut;
	wire _dataUnits_3_io_validOut;
	wire [127:0] _dataUnits_2_io_taskOut;
	wire _dataUnits_2_io_validOut;
	wire [127:0] _dataUnits_1_io_taskOut;
	wire _dataUnits_1_io_validOut;
	wire [127:0] _dataUnits_0_io_taskOut;
	wire _dataUnits_0_io_validOut;
	SchedulerNetworkDataUnit dataUnits_0(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_65_io_taskOut),
		.io_taskOut(_dataUnits_0_io_taskOut),
		.io_validIn(_dataUnits_65_io_validOut),
		.io_validOut(_dataUnits_0_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_0_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_0_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_0_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_0_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_0_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_0_data_qOutTask_bits),
		.io_occupied(io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerNetworkDataUnit dataUnits_1(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_0_io_taskOut),
		.io_taskOut(_dataUnits_1_io_taskOut),
		.io_validIn(_dataUnits_0_io_validOut),
		.io_validOut(_dataUnits_1_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_1_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_1_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_1_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_1_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_1_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_1_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_2(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_1_io_taskOut),
		.io_taskOut(_dataUnits_2_io_taskOut),
		.io_validIn(_dataUnits_1_io_validOut),
		.io_validOut(_dataUnits_2_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_2_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_2_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_2_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_2_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_2_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_2_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_3(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_2_io_taskOut),
		.io_taskOut(_dataUnits_3_io_taskOut),
		.io_validIn(_dataUnits_2_io_validOut),
		.io_validOut(_dataUnits_3_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_3_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_3_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_3_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_3_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_3_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_3_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_4(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_3_io_taskOut),
		.io_taskOut(_dataUnits_4_io_taskOut),
		.io_validIn(_dataUnits_3_io_validOut),
		.io_validOut(_dataUnits_4_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_4_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_4_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_4_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_4_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_4_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_4_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_5(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_4_io_taskOut),
		.io_taskOut(_dataUnits_5_io_taskOut),
		.io_validIn(_dataUnits_4_io_validOut),
		.io_validOut(_dataUnits_5_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_5_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_5_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_5_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_5_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_5_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_5_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_6(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_5_io_taskOut),
		.io_taskOut(_dataUnits_6_io_taskOut),
		.io_validIn(_dataUnits_5_io_validOut),
		.io_validOut(_dataUnits_6_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_6_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_6_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_6_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_6_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_6_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_6_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_7(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_6_io_taskOut),
		.io_taskOut(_dataUnits_7_io_taskOut),
		.io_validIn(_dataUnits_6_io_validOut),
		.io_validOut(_dataUnits_7_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_7_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_7_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_7_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_7_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_7_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_7_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_8(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_7_io_taskOut),
		.io_taskOut(_dataUnits_8_io_taskOut),
		.io_validIn(_dataUnits_7_io_validOut),
		.io_validOut(_dataUnits_8_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_8_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_8_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_8_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_8_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_8_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_8_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_9(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_8_io_taskOut),
		.io_taskOut(_dataUnits_9_io_taskOut),
		.io_validIn(_dataUnits_8_io_validOut),
		.io_validOut(_dataUnits_9_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_9_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_9_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_9_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_9_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_9_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_9_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_10(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_9_io_taskOut),
		.io_taskOut(_dataUnits_10_io_taskOut),
		.io_validIn(_dataUnits_9_io_validOut),
		.io_validOut(_dataUnits_10_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_10_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_10_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_10_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_10_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_10_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_10_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_11(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_10_io_taskOut),
		.io_taskOut(_dataUnits_11_io_taskOut),
		.io_validIn(_dataUnits_10_io_validOut),
		.io_validOut(_dataUnits_11_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_11_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_11_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_11_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_11_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_11_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_11_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_12(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_11_io_taskOut),
		.io_taskOut(_dataUnits_12_io_taskOut),
		.io_validIn(_dataUnits_11_io_validOut),
		.io_validOut(_dataUnits_12_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_12_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_12_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_12_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_12_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_12_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_12_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_13(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_12_io_taskOut),
		.io_taskOut(_dataUnits_13_io_taskOut),
		.io_validIn(_dataUnits_12_io_validOut),
		.io_validOut(_dataUnits_13_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_13_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_13_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_13_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_13_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_13_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_13_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_14(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_13_io_taskOut),
		.io_taskOut(_dataUnits_14_io_taskOut),
		.io_validIn(_dataUnits_13_io_validOut),
		.io_validOut(_dataUnits_14_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_14_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_14_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_14_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_14_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_14_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_14_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_15(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_14_io_taskOut),
		.io_taskOut(_dataUnits_15_io_taskOut),
		.io_validIn(_dataUnits_14_io_validOut),
		.io_validOut(_dataUnits_15_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_15_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_15_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_15_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_15_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_15_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_15_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_16(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_15_io_taskOut),
		.io_taskOut(_dataUnits_16_io_taskOut),
		.io_validIn(_dataUnits_15_io_validOut),
		.io_validOut(_dataUnits_16_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_16_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_16_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_16_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_16_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_16_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_16_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_17(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_16_io_taskOut),
		.io_taskOut(_dataUnits_17_io_taskOut),
		.io_validIn(_dataUnits_16_io_validOut),
		.io_validOut(_dataUnits_17_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_17_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_17_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_17_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_17_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_17_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_17_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_18(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_17_io_taskOut),
		.io_taskOut(_dataUnits_18_io_taskOut),
		.io_validIn(_dataUnits_17_io_validOut),
		.io_validOut(_dataUnits_18_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_18_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_18_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_18_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_18_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_18_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_18_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_19(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_18_io_taskOut),
		.io_taskOut(_dataUnits_19_io_taskOut),
		.io_validIn(_dataUnits_18_io_validOut),
		.io_validOut(_dataUnits_19_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_19_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_19_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_19_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_19_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_19_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_19_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_20(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_19_io_taskOut),
		.io_taskOut(_dataUnits_20_io_taskOut),
		.io_validIn(_dataUnits_19_io_validOut),
		.io_validOut(_dataUnits_20_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_20_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_20_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_20_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_20_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_20_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_20_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_21(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_20_io_taskOut),
		.io_taskOut(_dataUnits_21_io_taskOut),
		.io_validIn(_dataUnits_20_io_validOut),
		.io_validOut(_dataUnits_21_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_21_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_21_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_21_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_21_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_21_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_21_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_22(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_21_io_taskOut),
		.io_taskOut(_dataUnits_22_io_taskOut),
		.io_validIn(_dataUnits_21_io_validOut),
		.io_validOut(_dataUnits_22_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_22_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_22_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_22_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_22_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_22_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_22_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_23(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_22_io_taskOut),
		.io_taskOut(_dataUnits_23_io_taskOut),
		.io_validIn(_dataUnits_22_io_validOut),
		.io_validOut(_dataUnits_23_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_23_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_23_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_23_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_23_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_23_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_23_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_24(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_23_io_taskOut),
		.io_taskOut(_dataUnits_24_io_taskOut),
		.io_validIn(_dataUnits_23_io_validOut),
		.io_validOut(_dataUnits_24_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_24_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_24_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_24_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_24_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_24_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_24_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_25(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_24_io_taskOut),
		.io_taskOut(_dataUnits_25_io_taskOut),
		.io_validIn(_dataUnits_24_io_validOut),
		.io_validOut(_dataUnits_25_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_25_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_25_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_25_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_25_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_25_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_25_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_26(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_25_io_taskOut),
		.io_taskOut(_dataUnits_26_io_taskOut),
		.io_validIn(_dataUnits_25_io_validOut),
		.io_validOut(_dataUnits_26_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_26_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_26_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_26_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_26_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_26_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_26_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_27(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_26_io_taskOut),
		.io_taskOut(_dataUnits_27_io_taskOut),
		.io_validIn(_dataUnits_26_io_validOut),
		.io_validOut(_dataUnits_27_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_27_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_27_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_27_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_27_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_27_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_27_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_28(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_27_io_taskOut),
		.io_taskOut(_dataUnits_28_io_taskOut),
		.io_validIn(_dataUnits_27_io_validOut),
		.io_validOut(_dataUnits_28_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_28_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_28_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_28_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_28_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_28_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_28_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_29(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_28_io_taskOut),
		.io_taskOut(_dataUnits_29_io_taskOut),
		.io_validIn(_dataUnits_28_io_validOut),
		.io_validOut(_dataUnits_29_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_29_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_29_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_29_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_29_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_29_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_29_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_30(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_29_io_taskOut),
		.io_taskOut(_dataUnits_30_io_taskOut),
		.io_validIn(_dataUnits_29_io_validOut),
		.io_validOut(_dataUnits_30_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_30_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_30_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_30_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_30_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_30_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_30_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_31(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_30_io_taskOut),
		.io_taskOut(_dataUnits_31_io_taskOut),
		.io_validIn(_dataUnits_30_io_validOut),
		.io_validOut(_dataUnits_31_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_31_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_31_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_31_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_31_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_31_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_31_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_32(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_31_io_taskOut),
		.io_taskOut(_dataUnits_32_io_taskOut),
		.io_validIn(_dataUnits_31_io_validOut),
		.io_validOut(_dataUnits_32_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_32_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_32_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_32_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_32_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_32_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_32_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_33(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_32_io_taskOut),
		.io_taskOut(_dataUnits_33_io_taskOut),
		.io_validIn(_dataUnits_32_io_validOut),
		.io_validOut(_dataUnits_33_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_33_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_33_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_33_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_33_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_33_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_33_data_qOutTask_bits),
		.io_occupied(io_ntwDataUnitOccupancyVSS_1)
	);
	SchedulerNetworkDataUnit dataUnits_34(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_33_io_taskOut),
		.io_taskOut(_dataUnits_34_io_taskOut),
		.io_validIn(_dataUnits_33_io_validOut),
		.io_validOut(_dataUnits_34_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_34_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_34_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_34_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_34_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_34_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_34_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_35(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_34_io_taskOut),
		.io_taskOut(_dataUnits_35_io_taskOut),
		.io_validIn(_dataUnits_34_io_validOut),
		.io_validOut(_dataUnits_35_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_35_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_35_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_35_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_35_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_35_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_35_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_36(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_35_io_taskOut),
		.io_taskOut(_dataUnits_36_io_taskOut),
		.io_validIn(_dataUnits_35_io_validOut),
		.io_validOut(_dataUnits_36_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_36_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_36_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_36_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_36_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_36_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_36_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_37(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_36_io_taskOut),
		.io_taskOut(_dataUnits_37_io_taskOut),
		.io_validIn(_dataUnits_36_io_validOut),
		.io_validOut(_dataUnits_37_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_37_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_37_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_37_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_37_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_37_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_37_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_38(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_37_io_taskOut),
		.io_taskOut(_dataUnits_38_io_taskOut),
		.io_validIn(_dataUnits_37_io_validOut),
		.io_validOut(_dataUnits_38_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_38_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_38_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_38_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_38_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_38_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_38_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_39(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_38_io_taskOut),
		.io_taskOut(_dataUnits_39_io_taskOut),
		.io_validIn(_dataUnits_38_io_validOut),
		.io_validOut(_dataUnits_39_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_39_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_39_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_39_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_39_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_39_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_39_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_40(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_39_io_taskOut),
		.io_taskOut(_dataUnits_40_io_taskOut),
		.io_validIn(_dataUnits_39_io_validOut),
		.io_validOut(_dataUnits_40_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_40_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_40_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_40_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_40_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_40_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_40_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_41(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_40_io_taskOut),
		.io_taskOut(_dataUnits_41_io_taskOut),
		.io_validIn(_dataUnits_40_io_validOut),
		.io_validOut(_dataUnits_41_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_41_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_41_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_41_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_41_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_41_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_41_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_42(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_41_io_taskOut),
		.io_taskOut(_dataUnits_42_io_taskOut),
		.io_validIn(_dataUnits_41_io_validOut),
		.io_validOut(_dataUnits_42_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_42_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_42_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_42_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_42_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_42_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_42_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_43(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_42_io_taskOut),
		.io_taskOut(_dataUnits_43_io_taskOut),
		.io_validIn(_dataUnits_42_io_validOut),
		.io_validOut(_dataUnits_43_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_43_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_43_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_43_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_43_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_43_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_43_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_44(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_43_io_taskOut),
		.io_taskOut(_dataUnits_44_io_taskOut),
		.io_validIn(_dataUnits_43_io_validOut),
		.io_validOut(_dataUnits_44_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_44_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_44_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_44_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_44_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_44_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_44_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_45(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_44_io_taskOut),
		.io_taskOut(_dataUnits_45_io_taskOut),
		.io_validIn(_dataUnits_44_io_validOut),
		.io_validOut(_dataUnits_45_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_45_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_45_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_45_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_45_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_45_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_45_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_46(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_45_io_taskOut),
		.io_taskOut(_dataUnits_46_io_taskOut),
		.io_validIn(_dataUnits_45_io_validOut),
		.io_validOut(_dataUnits_46_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_46_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_46_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_46_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_46_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_46_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_46_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_47(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_46_io_taskOut),
		.io_taskOut(_dataUnits_47_io_taskOut),
		.io_validIn(_dataUnits_46_io_validOut),
		.io_validOut(_dataUnits_47_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_47_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_47_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_47_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_47_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_47_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_47_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_48(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_47_io_taskOut),
		.io_taskOut(_dataUnits_48_io_taskOut),
		.io_validIn(_dataUnits_47_io_validOut),
		.io_validOut(_dataUnits_48_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_48_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_48_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_48_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_48_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_48_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_48_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_49(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_48_io_taskOut),
		.io_taskOut(_dataUnits_49_io_taskOut),
		.io_validIn(_dataUnits_48_io_validOut),
		.io_validOut(_dataUnits_49_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_49_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_49_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_49_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_49_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_49_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_49_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_50(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_49_io_taskOut),
		.io_taskOut(_dataUnits_50_io_taskOut),
		.io_validIn(_dataUnits_49_io_validOut),
		.io_validOut(_dataUnits_50_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_50_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_50_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_50_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_50_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_50_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_50_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_51(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_50_io_taskOut),
		.io_taskOut(_dataUnits_51_io_taskOut),
		.io_validIn(_dataUnits_50_io_validOut),
		.io_validOut(_dataUnits_51_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_51_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_51_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_51_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_51_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_51_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_51_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_52(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_51_io_taskOut),
		.io_taskOut(_dataUnits_52_io_taskOut),
		.io_validIn(_dataUnits_51_io_validOut),
		.io_validOut(_dataUnits_52_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_52_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_52_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_52_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_52_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_52_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_52_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_53(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_52_io_taskOut),
		.io_taskOut(_dataUnits_53_io_taskOut),
		.io_validIn(_dataUnits_52_io_validOut),
		.io_validOut(_dataUnits_53_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_53_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_53_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_53_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_53_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_53_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_53_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_54(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_53_io_taskOut),
		.io_taskOut(_dataUnits_54_io_taskOut),
		.io_validIn(_dataUnits_53_io_validOut),
		.io_validOut(_dataUnits_54_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_54_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_54_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_54_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_54_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_54_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_54_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_55(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_54_io_taskOut),
		.io_taskOut(_dataUnits_55_io_taskOut),
		.io_validIn(_dataUnits_54_io_validOut),
		.io_validOut(_dataUnits_55_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_55_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_55_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_55_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_55_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_55_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_55_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_56(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_55_io_taskOut),
		.io_taskOut(_dataUnits_56_io_taskOut),
		.io_validIn(_dataUnits_55_io_validOut),
		.io_validOut(_dataUnits_56_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_56_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_56_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_56_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_56_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_56_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_56_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_57(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_56_io_taskOut),
		.io_taskOut(_dataUnits_57_io_taskOut),
		.io_validIn(_dataUnits_56_io_validOut),
		.io_validOut(_dataUnits_57_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_57_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_57_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_57_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_57_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_57_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_57_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_58(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_57_io_taskOut),
		.io_taskOut(_dataUnits_58_io_taskOut),
		.io_validIn(_dataUnits_57_io_validOut),
		.io_validOut(_dataUnits_58_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_58_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_58_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_58_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_58_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_58_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_58_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_59(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_58_io_taskOut),
		.io_taskOut(_dataUnits_59_io_taskOut),
		.io_validIn(_dataUnits_58_io_validOut),
		.io_validOut(_dataUnits_59_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_59_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_59_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_59_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_59_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_59_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_59_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_60(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_59_io_taskOut),
		.io_taskOut(_dataUnits_60_io_taskOut),
		.io_validIn(_dataUnits_59_io_validOut),
		.io_validOut(_dataUnits_60_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_60_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_60_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_60_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_60_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_60_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_60_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_61(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_60_io_taskOut),
		.io_taskOut(_dataUnits_61_io_taskOut),
		.io_validIn(_dataUnits_60_io_validOut),
		.io_validOut(_dataUnits_61_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_61_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_61_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_61_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_61_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_61_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_61_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_62(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_61_io_taskOut),
		.io_taskOut(_dataUnits_62_io_taskOut),
		.io_validIn(_dataUnits_61_io_validOut),
		.io_validOut(_dataUnits_62_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_62_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_62_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_62_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_62_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_62_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_62_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_63(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_62_io_taskOut),
		.io_taskOut(_dataUnits_63_io_taskOut),
		.io_validIn(_dataUnits_62_io_validOut),
		.io_validOut(_dataUnits_63_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_63_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_63_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_63_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_63_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_63_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_63_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_64(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_63_io_taskOut),
		.io_taskOut(_dataUnits_64_io_taskOut),
		.io_validIn(_dataUnits_63_io_validOut),
		.io_validOut(_dataUnits_64_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_64_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_64_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_64_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_64_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_64_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_64_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_65(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_64_io_taskOut),
		.io_taskOut(_dataUnits_65_io_taskOut),
		.io_validIn(_dataUnits_64_io_validOut),
		.io_validOut(_dataUnits_65_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_65_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_65_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_65_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_65_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_65_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_65_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkControlUnit ctrlunits_0(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_1_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_0_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_0_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_0_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_1(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_2_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_1_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_1_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_1_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_1_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_1_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_2(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_3_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_2_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_2_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_2_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_2_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_2_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_3(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_4_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_3_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_3_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_3_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_3_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_3_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_4(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_5_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_4_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_4_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_4_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_4_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_4_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_5(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_6_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_5_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_5_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_5_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_5_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_5_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_6(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_7_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_6_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_6_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_6_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_6_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_6_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_7(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_8_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_7_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_7_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_7_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_7_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_7_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_8(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_9_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_8_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_8_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_8_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_8_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_8_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_9(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_10_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_9_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_9_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_9_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_9_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_9_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_10(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_11_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_10_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_10_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_10_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_10_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_10_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_11(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_12_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_11_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_11_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_11_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_11_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_11_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_12(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_13_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_12_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_12_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_12_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_12_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_12_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_13(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_14_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_13_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_13_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_13_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_13_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_13_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_14(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_15_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_14_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_14_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_14_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_14_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_14_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_15(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_16_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_15_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_15_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_15_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_15_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_15_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_16(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_17_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_16_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_16_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_16_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_16_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_16_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_17(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_18_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_17_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_17_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_17_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_17_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_18(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_19_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_18_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_18_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_18_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_18_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_19(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_20_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_19_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_19_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_19_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_19_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_20(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_21_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_20_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_20_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_20_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_20_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_21(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_22_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_21_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_21_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_21_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_21_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_22(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_23_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_22_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_22_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_22_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_22_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_23(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_24_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_23_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_23_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_23_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_23_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_24(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_25_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_24_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_24_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_24_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_24_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_25(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_26_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_25_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_25_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_25_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_25_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_26(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_27_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_26_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_26_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_26_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_26_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_27(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_28_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_27_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_27_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_27_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_27_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_28(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_29_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_28_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_28_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_28_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_28_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_29(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_30_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_29_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_29_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_29_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_29_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_30(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_31_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_30_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_30_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_30_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_30_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_31(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_32_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_31_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_31_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_31_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_31_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_32(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_33_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_32_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_32_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_32_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_32_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_33(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_34_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_33_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_33_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_33_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_34(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_35_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_34_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_34_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_34_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_34_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_34_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_35(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_36_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_35_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_35_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_35_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_35_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_35_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_36(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_37_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_36_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_36_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_36_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_36_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_36_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_37(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_38_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_37_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_37_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_37_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_37_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_37_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_38(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_39_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_38_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_38_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_38_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_38_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_38_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_39(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_40_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_39_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_39_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_39_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_39_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_39_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_40(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_41_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_40_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_40_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_40_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_40_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_40_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_41(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_42_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_41_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_41_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_41_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_41_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_41_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_42(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_43_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_42_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_42_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_42_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_42_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_42_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_43(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_44_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_43_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_43_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_43_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_43_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_43_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_44(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_45_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_44_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_44_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_44_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_44_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_44_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_45(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_46_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_45_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_45_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_45_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_45_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_45_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_46(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_47_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_46_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_46_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_46_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_46_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_46_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_47(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_48_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_47_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_47_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_47_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_47_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_47_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_48(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_49_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_48_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_48_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_48_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_48_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_48_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_49(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_50_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_49_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_49_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_49_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_49_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_49_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_50(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_51_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_50_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_50_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_50_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_50_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_50_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_51(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_52_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_51_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_51_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_51_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_51_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_51_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_52(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_53_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_52_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_52_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_52_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_52_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_52_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_53(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_54_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_53_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_53_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_53_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_53_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_53_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_54(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_55_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_54_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_54_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_54_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_54_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_54_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_55(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_56_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_55_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_55_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_55_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_55_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_55_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_56(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_57_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_56_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_56_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_56_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_56_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_56_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_57(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_58_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_57_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_57_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_57_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_57_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_57_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_58(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_59_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_58_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_58_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_58_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_58_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_58_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_59(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_60_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_59_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_59_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_59_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_59_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_59_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_60(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_61_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_60_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_60_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_60_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_60_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_60_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_61(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_62_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_61_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_61_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_61_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_61_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_61_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_62(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_63_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_62_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_62_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_62_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_62_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_62_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_63(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_64_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_63_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_63_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_63_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_63_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_63_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_64(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_65_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_64_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_64_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_64_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_64_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_64_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_65(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_0_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_65_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_65_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_65_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_65_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_65_ctrl_stealReq_ready)
	);
endmodule
module SchedulerClient (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_ctrl_stealReq_valid,
	io_connNetwork_ctrl_stealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_connQ_currLength,
	io_connQ_push_ready,
	io_connQ_push_valid,
	io_connQ_push_bits,
	io_connQ_pop_ready,
	io_connQ_pop_valid,
	io_connQ_pop_bits
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_ctrl_stealReq_valid;
	input io_connNetwork_ctrl_stealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [127:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [127:0] io_connNetwork_data_qOutTask_bits;
	input [3:0] io_connQ_currLength;
	input io_connQ_push_ready;
	output wire io_connQ_push_valid;
	output wire [127:0] io_connQ_push_bits;
	output wire io_connQ_pop_ready;
	input io_connQ_pop_valid;
	input [127:0] io_connQ_pop_bits;
	reg [2:0] stateReg;
	reg [127:0] stolenTaskReg;
	reg [127:0] giveTaskReg;
	reg [1:0] taskRequestCount;
	reg [31:0] tasksGivenAwayCount;
	reg [31:0] requestKilledCount;
	reg [31:0] requestFullCount;
	wire _GEN = stateReg == 3'h0;
	wire _GEN_0 = stateReg == 3'h1;
	wire _GEN_1 = io_connNetwork_ctrl_stealReq_ready & (taskRequestCount == 2'h1);
	wire _GEN_2 = io_connNetwork_ctrl_stealReq_ready & (taskRequestCount == 2'h2);
	wire _GEN_3 = _GEN_2 | (|io_connQ_currLength);
	wire _GEN_4 = _GEN_1 | _GEN_3;
	wire _GEN_5 = stateReg == 3'h2;
	wire _GEN_6 = _GEN | _GEN_0;
	wire _GEN_7 = stateReg == 3'h3;
	wire _GEN_8 = (_GEN | _GEN_0) | _GEN_5;
	wire _GEN_9 = stateReg == 3'h4;
	wire _GEN_10 = stateReg == 3'h5;
	wire _GEN_11 = (_GEN_5 | _GEN_7) | _GEN_9;
	wire _GEN_12 = (_GEN | _GEN_0) | _GEN_11;
	wire _GEN_13 = stateReg == 3'h6;
	wire _GEN_14 = ((_GEN_5 | _GEN_7) | _GEN_9) | _GEN_10;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 3'h0;
			stolenTaskReg <= 128'h00000000000000000000000000000000;
			giveTaskReg <= 128'h00000000000000000000000000000000;
			taskRequestCount <= 2'h1;
			tasksGivenAwayCount <= 32'h00000000;
			requestKilledCount <= 32'h00000042;
			requestFullCount <= 32'h00000042;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_15;
			reg _GEN_16;
			reg _GEN_17;
			reg _GEN_18;
			reg [31:0] _GEN_19;
			reg _GEN_20;
			reg _GEN_21;
			reg _GEN_22;
			reg [1:0] _GEN_23;
			reg [23:0] _GEN_24;
			reg [15:0] _GEN_25;
			reg [255:0] _GEN_26;
			_GEN_16 = io_connQ_currLength > 4'h5;
			_GEN_19 = (_GEN_11 | ~(_GEN_10 & io_connNetwork_data_qOutTask_ready) ? tasksGivenAwayCount : tasksGivenAwayCount + 32'h00000001);
			_GEN_26 = {_GEN_19, _GEN_19, _GEN_19, tasksGivenAwayCount, tasksGivenAwayCount, tasksGivenAwayCount, (_GEN_4 | ~(|tasksGivenAwayCount) ? tasksGivenAwayCount : tasksGivenAwayCount - 32'h00000001), tasksGivenAwayCount};
			_GEN_15 = io_connQ_currLength == 4'h0;
			_GEN_17 = requestKilledCount == 32'h00000000;
			_GEN_18 = io_connQ_currLength > 4'h4;
			_GEN_20 = _GEN_16 | (io_connNetwork_ctrl_serveStealReq_ready & |io_connQ_currLength);
			_GEN_21 = _GEN_15 & io_connNetwork_ctrl_serveStealReq_ready;
			_GEN_22 = _GEN_21 | _GEN_15;
			_GEN_23 = ((_GEN_14 | ~_GEN_13) | _GEN_20 ? taskRequestCount : (_GEN_21 ? 2'h2 : (_GEN_15 ? 2'h1 : taskRequestCount)));
			_GEN_24 = {stateReg, (_GEN_20 ? 3'h4 : (_GEN_22 ? 3'h1 : 3'h6)), (io_connNetwork_data_qOutTask_ready ? 3'h0 : 3'h5), (io_connQ_pop_valid ? 3'h5 : (_GEN_15 ? 3'h1 : 3'h4)), (io_connQ_push_ready ? 3'h0 : (_GEN_18 ? 3'h5 : 3'h3)), (io_connNetwork_data_availableTask_valid ? 3'h3 : (|io_connQ_currLength ? 3'h0 : (_GEN_17 ? 3'h1 : 3'h2))), (_GEN_1 ? 3'h2 : (_GEN_2 ? 3'h1 : (|io_connQ_currLength ? 3'h6 : (|tasksGivenAwayCount | (requestFullCount == 32'h00000000) ? 3'h2 : 3'h1)))), (_GEN_15 ? 3'h1 : (_GEN_16 ? 3'h4 : (|io_connQ_currLength[3:1] ? 3'h6 : 3'h0)))};
			stateReg <= _GEN_24[stateReg * 3+:3];
			if (_GEN_6 | ~(_GEN_5 & io_connNetwork_data_availableTask_valid))
				;
			else
				stolenTaskReg <= io_connNetwork_data_availableTask_bits;
			if (~_GEN_8) begin
				if (_GEN_7) begin
					if (io_connQ_push_ready | ~_GEN_18)
						;
					else
						giveTaskReg <= stolenTaskReg;
				end
				else if (_GEN_9 & io_connQ_pop_valid)
					giveTaskReg <= io_connQ_pop_bits;
			end
			_GEN_25 = {_GEN_23, _GEN_23, taskRequestCount, taskRequestCount, taskRequestCount, taskRequestCount, (_GEN_1 | ~_GEN_2 ? taskRequestCount : 2'h1), taskRequestCount};
			taskRequestCount <= _GEN_25[stateReg * 2+:2];
			tasksGivenAwayCount <= _GEN_26[stateReg * 32+:32];
			if (_GEN) begin
				if (_GEN_15)
					requestFullCount <= 32'h00000042;
			end
			else if (_GEN_0) begin
				if (_GEN_1 | ~(_GEN_3 | ~(|tasksGivenAwayCount)))
					requestKilledCount <= 32'h00000042;
				if (io_connNetwork_ctrl_serveStealReq_ready)
					requestFullCount <= requestFullCount - 32'h00000001;
				else
					requestFullCount <= 32'h00000042;
			end
			else begin
				if (_GEN_5) begin
					if (io_connNetwork_ctrl_serveStealReq_ready)
						requestKilledCount <= 32'h00000042;
					else
						requestKilledCount <= requestKilledCount - 32'h00000001;
				end
				if ((_GEN_5 ? (io_connNetwork_data_availableTask_valid | (|io_connQ_currLength)) | ~_GEN_17 : _GEN_7 | (_GEN_9 ? io_connQ_pop_valid | ~_GEN_15 : ((_GEN_10 | ~_GEN_13) | _GEN_20) | ~_GEN_22)))
					;
				else
					requestFullCount <= 32'h00000042;
			end
		end
	assign io_connNetwork_ctrl_serveStealReq_valid = ~_GEN & (_GEN_0 ? ~_GEN_4 & |tasksGivenAwayCount : ~_GEN_14 & _GEN_13);
	assign io_connNetwork_ctrl_stealReq_valid = ~_GEN & _GEN_0;
	assign io_connNetwork_data_availableTask_ready = ~_GEN_6 & _GEN_5;
	assign io_connNetwork_data_qOutTask_valid = ~_GEN_12 & _GEN_10;
	assign io_connNetwork_data_qOutTask_bits = (_GEN_12 | ~_GEN_10 ? 128'h00000000000000000000000000000000 : giveTaskReg);
	assign io_connQ_push_valid = ~_GEN_8 & _GEN_7;
	assign io_connQ_push_bits = (_GEN_8 | ~_GEN_7 ? 128'h00000000000000000000000000000000 : stolenTaskReg);
	assign io_connQ_pop_ready = ~(((_GEN | _GEN_0) | _GEN_5) | _GEN_7) & _GEN_9;
endmodule
module hw_deque (
	clock,
	reset,
	io_connVec_0_push_ready,
	io_connVec_0_push_valid,
	io_connVec_0_push_bits,
	io_connVec_0_pop_ready,
	io_connVec_0_pop_valid,
	io_connVec_0_pop_bits,
	io_connVec_1_currLength,
	io_connVec_1_push_ready,
	io_connVec_1_push_valid,
	io_connVec_1_push_bits,
	io_connVec_1_pop_ready,
	io_connVec_1_pop_valid,
	io_connVec_1_pop_bits
);
	input clock;
	input reset;
	output wire io_connVec_0_push_ready;
	input io_connVec_0_push_valid;
	input [127:0] io_connVec_0_push_bits;
	input io_connVec_0_pop_ready;
	output wire io_connVec_0_pop_valid;
	output wire [127:0] io_connVec_0_pop_bits;
	output wire [4:0] io_connVec_1_currLength;
	output wire io_connVec_1_push_ready;
	input io_connVec_1_push_valid;
	input [127:0] io_connVec_1_push_bits;
	input io_connVec_1_pop_ready;
	output wire io_connVec_1_pop_valid;
	output wire [127:0] io_connVec_1_pop_bits;
	wire [127:0] _bramMem_a_dout;
	wire [127:0] _bramMem_b_dout;
	reg [4:0] sideReg_0;
	reg [4:0] sideReg_1;
	reg readLatency_0;
	reg readLatency_1;
	reg writeLatency_0;
	reg writeLatency_1;
	reg [2:0] stateRegs_0;
	reg [2:0] stateRegs_1;
	wire _GEN = stateRegs_0 == 3'h0;
	wire _GEN_0 = stateRegs_1 == 3'h0;
	wire _GEN_1 = stateRegs_0 == 3'h1;
	wire _GEN_2 = stateRegs_0 == 3'h2;
	wire _GEN_3 = sideReg_0 == 5'h09;
	wire _GEN_4 = stateRegs_0 == 3'h4;
	wire [4:0] _bramMem_io_a_addr_T_2 = sideReg_0 + 5'h01;
	wire _GEN_5 = (_GEN | _GEN_1) | _GEN_2;
	wire _GEN_6 = stateRegs_0 == 3'h3;
	wire _GEN_7 = stateRegs_1 == 3'h1;
	wire _GEN_8 = stateRegs_1 == 3'h2;
	wire _GEN_9 = sideReg_1 == 5'h00;
	wire _GEN_10 = stateRegs_1 == 3'h4;
	wire [4:0] _bramMem_io_b_addr_T_6 = sideReg_1 - 5'h01;
	wire _GEN_11 = (_GEN_0 | _GEN_7) | _GEN_8;
	wire _GEN_12 = stateRegs_1 == 3'h3;
	wire [4:0] currLen = (sideReg_0 > sideReg_1 ? ((sideReg_1 + 5'h0a) - sideReg_0) - 5'h01 : (sideReg_1 - sideReg_0) - 5'h01);
	always @(posedge clock)
		if (reset) begin
			sideReg_0 <= 5'h00;
			sideReg_1 <= 5'h01;
			readLatency_0 <= 1'h0;
			readLatency_1 <= 1'h0;
			writeLatency_0 <= 1'h0;
			writeLatency_1 <= 1'h0;
			stateRegs_0 <= 3'h0;
			stateRegs_1 <= 3'h0;
		end
		else begin : sv2v_autoblock_1
			reg [23:0] _GEN_13;
			reg [23:0] _GEN_14;
			_GEN_13 = {stateRegs_0, stateRegs_0, stateRegs_0, 6'h00, (readLatency_0 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_0, 1'h1, ((io_connVec_0_pop_ready & |currLen[4:1]) | ((io_connVec_0_pop_ready & _GEN_0) & |currLen) ? 3'h2 : {2'h0, io_connVec_0_push_valid & (currLen < 5'h0a)})};
			_GEN_14 = {stateRegs_1, stateRegs_1, stateRegs_1, 6'h00, (readLatency_1 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_1, 1'h1, (io_connVec_1_push_valid & (currLen < 5'h09) ? 3'h1 : {1'h0, (io_connVec_1_pop_ready & |currLen[4:1]) | (((io_connVec_1_pop_ready & ~io_connVec_0_pop_ready) & |currLen) & (stateRegs_0 != 3'h4)), 1'h0})};
			if (~_GEN_5) begin
				if (_GEN_4) begin
					if (_GEN_3)
						sideReg_0 <= 5'h00;
					else
						sideReg_0 <= _bramMem_io_a_addr_T_2;
				end
				else if (_GEN_6) begin
					if (sideReg_0 == 5'h00)
						sideReg_0 <= 5'h09;
					else
						sideReg_0 <= sideReg_0 - 5'h01;
				end
			end
			if (~_GEN_11) begin
				if (_GEN_10) begin
					if (_GEN_9)
						sideReg_1 <= 5'h09;
					else
						sideReg_1 <= _bramMem_io_b_addr_T_6;
				end
				else if (_GEN_12) begin
					if (sideReg_1 == 5'h09)
						sideReg_1 <= 5'h00;
					else
						sideReg_1 <= sideReg_1 + 5'h01;
				end
			end
			readLatency_0 <= (((_GEN | _GEN_1) | ~_GEN_2) | (readLatency_0 - 1'h1)) & readLatency_0;
			readLatency_1 <= (((_GEN_0 | _GEN_7) | ~_GEN_8) | (readLatency_1 - 1'h1)) & readLatency_1;
			writeLatency_0 <= ((_GEN | ~_GEN_1) | (writeLatency_0 - 1'h1)) & writeLatency_0;
			writeLatency_1 <= ((_GEN_0 | ~_GEN_7) | (writeLatency_1 - 1'h1)) & writeLatency_1;
			stateRegs_0 <= _GEN_13[stateRegs_0 * 3+:3];
			stateRegs_1 <= _GEN_14[stateRegs_1 * 3+:3];
		end
	DualPortBRAM #(
		.ADDR(6),
		.DATA(128)
	) bramMem(
		.clk(clock),
		.rst(reset),
		.a_addr((_GEN ? 6'h3f : (_GEN_1 ? {1'h0, sideReg_0} : (_GEN_2 ? (_GEN_3 ? 6'h00 : {1'h0, sideReg_0 + 5'h01}) : (_GEN_4 ? (_GEN_3 ? 6'h00 : {1'h0, _bramMem_io_a_addr_T_2}) : 6'h3f))))),
		.a_din(io_connVec_0_push_bits),
		.a_wr(~_GEN & _GEN_1),
		.a_dout(_bramMem_a_dout),
		.b_addr((_GEN_0 ? 6'h3f : (_GEN_7 ? {1'h0, sideReg_1} : (_GEN_8 ? (_GEN_9 ? 6'h09 : {1'h0, sideReg_1 - 5'h01}) : (_GEN_10 ? (_GEN_9 ? 6'h09 : {1'h0, _bramMem_io_b_addr_T_6}) : 6'h3f))))),
		.b_din(io_connVec_1_push_bits),
		.b_wr(~_GEN_0 & _GEN_7),
		.b_dout(_bramMem_b_dout)
	);
	assign io_connVec_0_push_ready = ~(((_GEN | _GEN_1) | _GEN_2) | _GEN_4) & _GEN_6;
	assign io_connVec_0_pop_valid = ~_GEN_5 & _GEN_4;
	assign io_connVec_0_pop_bits = (_GEN_5 | ~_GEN_4 ? 128'h00000000000000000000000000000000 : _bramMem_a_dout);
	assign io_connVec_1_currLength = currLen;
	assign io_connVec_1_push_ready = ~(((_GEN_0 | _GEN_7) | _GEN_8) | _GEN_10) & _GEN_12;
	assign io_connVec_1_pop_valid = ~_GEN_11 & _GEN_10;
	assign io_connVec_1_pop_bits = (_GEN_11 | ~_GEN_10 ? 128'h00000000000000000000000000000000 : _bramMem_b_dout);
endmodule
module SchedulerLocalNetwork (
	clock,
	reset,
	io_connPE_0_push_ready,
	io_connPE_0_push_valid,
	io_connPE_0_push_bits,
	io_connPE_0_pop_ready,
	io_connPE_0_pop_valid,
	io_connPE_0_pop_bits,
	io_connPE_1_push_ready,
	io_connPE_1_push_valid,
	io_connPE_1_push_bits,
	io_connPE_1_pop_ready,
	io_connPE_1_pop_valid,
	io_connPE_1_pop_bits,
	io_connPE_2_push_ready,
	io_connPE_2_push_valid,
	io_connPE_2_push_bits,
	io_connPE_2_pop_ready,
	io_connPE_2_pop_valid,
	io_connPE_2_pop_bits,
	io_connPE_3_push_ready,
	io_connPE_3_push_valid,
	io_connPE_3_push_bits,
	io_connPE_3_pop_ready,
	io_connPE_3_pop_valid,
	io_connPE_3_pop_bits,
	io_connPE_4_push_ready,
	io_connPE_4_push_valid,
	io_connPE_4_push_bits,
	io_connPE_4_pop_ready,
	io_connPE_4_pop_valid,
	io_connPE_4_pop_bits,
	io_connPE_5_push_ready,
	io_connPE_5_push_valid,
	io_connPE_5_push_bits,
	io_connPE_5_pop_ready,
	io_connPE_5_pop_valid,
	io_connPE_5_pop_bits,
	io_connPE_6_push_ready,
	io_connPE_6_push_valid,
	io_connPE_6_push_bits,
	io_connPE_6_pop_ready,
	io_connPE_6_pop_valid,
	io_connPE_6_pop_bits,
	io_connPE_7_push_ready,
	io_connPE_7_push_valid,
	io_connPE_7_push_bits,
	io_connPE_7_pop_ready,
	io_connPE_7_pop_valid,
	io_connPE_7_pop_bits,
	io_connPE_8_push_ready,
	io_connPE_8_push_valid,
	io_connPE_8_push_bits,
	io_connPE_8_pop_ready,
	io_connPE_8_pop_valid,
	io_connPE_8_pop_bits,
	io_connPE_9_push_ready,
	io_connPE_9_push_valid,
	io_connPE_9_push_bits,
	io_connPE_9_pop_ready,
	io_connPE_9_pop_valid,
	io_connPE_9_pop_bits,
	io_connPE_10_push_ready,
	io_connPE_10_push_valid,
	io_connPE_10_push_bits,
	io_connPE_10_pop_ready,
	io_connPE_10_pop_valid,
	io_connPE_10_pop_bits,
	io_connPE_11_push_ready,
	io_connPE_11_push_valid,
	io_connPE_11_push_bits,
	io_connPE_11_pop_ready,
	io_connPE_11_pop_valid,
	io_connPE_11_pop_bits,
	io_connPE_12_push_ready,
	io_connPE_12_push_valid,
	io_connPE_12_push_bits,
	io_connPE_12_pop_ready,
	io_connPE_12_pop_valid,
	io_connPE_12_pop_bits,
	io_connPE_13_push_ready,
	io_connPE_13_push_valid,
	io_connPE_13_push_bits,
	io_connPE_13_pop_ready,
	io_connPE_13_pop_valid,
	io_connPE_13_pop_bits,
	io_connPE_14_push_ready,
	io_connPE_14_push_valid,
	io_connPE_14_push_bits,
	io_connPE_14_pop_ready,
	io_connPE_14_pop_valid,
	io_connPE_14_pop_bits,
	io_connPE_15_push_ready,
	io_connPE_15_push_valid,
	io_connPE_15_push_bits,
	io_connPE_15_pop_ready,
	io_connPE_15_pop_valid,
	io_connPE_15_pop_bits,
	io_connPE_16_push_ready,
	io_connPE_16_push_valid,
	io_connPE_16_push_bits,
	io_connPE_16_pop_ready,
	io_connPE_16_pop_valid,
	io_connPE_16_pop_bits,
	io_connPE_17_push_ready,
	io_connPE_17_push_valid,
	io_connPE_17_push_bits,
	io_connPE_17_pop_ready,
	io_connPE_17_pop_valid,
	io_connPE_17_pop_bits,
	io_connPE_18_push_ready,
	io_connPE_18_push_valid,
	io_connPE_18_push_bits,
	io_connPE_18_pop_ready,
	io_connPE_18_pop_valid,
	io_connPE_18_pop_bits,
	io_connPE_19_push_ready,
	io_connPE_19_push_valid,
	io_connPE_19_push_bits,
	io_connPE_19_pop_ready,
	io_connPE_19_pop_valid,
	io_connPE_19_pop_bits,
	io_connPE_20_push_ready,
	io_connPE_20_push_valid,
	io_connPE_20_push_bits,
	io_connPE_20_pop_ready,
	io_connPE_20_pop_valid,
	io_connPE_20_pop_bits,
	io_connPE_21_push_ready,
	io_connPE_21_push_valid,
	io_connPE_21_push_bits,
	io_connPE_21_pop_ready,
	io_connPE_21_pop_valid,
	io_connPE_21_pop_bits,
	io_connPE_22_push_ready,
	io_connPE_22_push_valid,
	io_connPE_22_push_bits,
	io_connPE_22_pop_ready,
	io_connPE_22_pop_valid,
	io_connPE_22_pop_bits,
	io_connPE_23_push_ready,
	io_connPE_23_push_valid,
	io_connPE_23_push_bits,
	io_connPE_23_pop_ready,
	io_connPE_23_pop_valid,
	io_connPE_23_pop_bits,
	io_connPE_24_push_ready,
	io_connPE_24_push_valid,
	io_connPE_24_push_bits,
	io_connPE_24_pop_ready,
	io_connPE_24_pop_valid,
	io_connPE_24_pop_bits,
	io_connPE_25_push_ready,
	io_connPE_25_push_valid,
	io_connPE_25_push_bits,
	io_connPE_25_pop_ready,
	io_connPE_25_pop_valid,
	io_connPE_25_pop_bits,
	io_connPE_26_push_ready,
	io_connPE_26_push_valid,
	io_connPE_26_push_bits,
	io_connPE_26_pop_ready,
	io_connPE_26_pop_valid,
	io_connPE_26_pop_bits,
	io_connPE_27_push_ready,
	io_connPE_27_push_valid,
	io_connPE_27_push_bits,
	io_connPE_27_pop_ready,
	io_connPE_27_pop_valid,
	io_connPE_27_pop_bits,
	io_connPE_28_push_ready,
	io_connPE_28_push_valid,
	io_connPE_28_push_bits,
	io_connPE_28_pop_ready,
	io_connPE_28_pop_valid,
	io_connPE_28_pop_bits,
	io_connPE_29_push_ready,
	io_connPE_29_push_valid,
	io_connPE_29_push_bits,
	io_connPE_29_pop_ready,
	io_connPE_29_pop_valid,
	io_connPE_29_pop_bits,
	io_connPE_30_push_ready,
	io_connPE_30_push_valid,
	io_connPE_30_push_bits,
	io_connPE_30_pop_ready,
	io_connPE_30_pop_valid,
	io_connPE_30_pop_bits,
	io_connPE_31_push_ready,
	io_connPE_31_push_valid,
	io_connPE_31_push_bits,
	io_connPE_31_pop_ready,
	io_connPE_31_pop_valid,
	io_connPE_31_pop_bits,
	io_connPE_32_push_ready,
	io_connPE_32_push_valid,
	io_connPE_32_push_bits,
	io_connPE_32_pop_ready,
	io_connPE_32_pop_valid,
	io_connPE_32_pop_bits,
	io_connPE_33_push_ready,
	io_connPE_33_push_valid,
	io_connPE_33_push_bits,
	io_connPE_33_pop_ready,
	io_connPE_33_pop_valid,
	io_connPE_33_pop_bits,
	io_connPE_34_push_ready,
	io_connPE_34_push_valid,
	io_connPE_34_push_bits,
	io_connPE_34_pop_ready,
	io_connPE_34_pop_valid,
	io_connPE_34_pop_bits,
	io_connPE_35_push_ready,
	io_connPE_35_push_valid,
	io_connPE_35_push_bits,
	io_connPE_35_pop_ready,
	io_connPE_35_pop_valid,
	io_connPE_35_pop_bits,
	io_connPE_36_push_ready,
	io_connPE_36_push_valid,
	io_connPE_36_push_bits,
	io_connPE_36_pop_ready,
	io_connPE_36_pop_valid,
	io_connPE_36_pop_bits,
	io_connPE_37_push_ready,
	io_connPE_37_push_valid,
	io_connPE_37_push_bits,
	io_connPE_37_pop_ready,
	io_connPE_37_pop_valid,
	io_connPE_37_pop_bits,
	io_connPE_38_push_ready,
	io_connPE_38_push_valid,
	io_connPE_38_push_bits,
	io_connPE_38_pop_ready,
	io_connPE_38_pop_valid,
	io_connPE_38_pop_bits,
	io_connPE_39_push_ready,
	io_connPE_39_push_valid,
	io_connPE_39_push_bits,
	io_connPE_39_pop_ready,
	io_connPE_39_pop_valid,
	io_connPE_39_pop_bits,
	io_connPE_40_push_ready,
	io_connPE_40_push_valid,
	io_connPE_40_push_bits,
	io_connPE_40_pop_ready,
	io_connPE_40_pop_valid,
	io_connPE_40_pop_bits,
	io_connPE_41_push_ready,
	io_connPE_41_push_valid,
	io_connPE_41_push_bits,
	io_connPE_41_pop_ready,
	io_connPE_41_pop_valid,
	io_connPE_41_pop_bits,
	io_connPE_42_push_ready,
	io_connPE_42_push_valid,
	io_connPE_42_push_bits,
	io_connPE_42_pop_ready,
	io_connPE_42_pop_valid,
	io_connPE_42_pop_bits,
	io_connPE_43_push_ready,
	io_connPE_43_push_valid,
	io_connPE_43_push_bits,
	io_connPE_43_pop_ready,
	io_connPE_43_pop_valid,
	io_connPE_43_pop_bits,
	io_connPE_44_push_ready,
	io_connPE_44_push_valid,
	io_connPE_44_push_bits,
	io_connPE_44_pop_ready,
	io_connPE_44_pop_valid,
	io_connPE_44_pop_bits,
	io_connPE_45_push_ready,
	io_connPE_45_push_valid,
	io_connPE_45_push_bits,
	io_connPE_45_pop_ready,
	io_connPE_45_pop_valid,
	io_connPE_45_pop_bits,
	io_connPE_46_push_ready,
	io_connPE_46_push_valid,
	io_connPE_46_push_bits,
	io_connPE_46_pop_ready,
	io_connPE_46_pop_valid,
	io_connPE_46_pop_bits,
	io_connPE_47_push_ready,
	io_connPE_47_push_valid,
	io_connPE_47_push_bits,
	io_connPE_47_pop_ready,
	io_connPE_47_pop_valid,
	io_connPE_47_pop_bits,
	io_connPE_48_push_ready,
	io_connPE_48_push_valid,
	io_connPE_48_push_bits,
	io_connPE_48_pop_ready,
	io_connPE_48_pop_valid,
	io_connPE_48_pop_bits,
	io_connPE_49_push_ready,
	io_connPE_49_push_valid,
	io_connPE_49_push_bits,
	io_connPE_49_pop_ready,
	io_connPE_49_pop_valid,
	io_connPE_49_pop_bits,
	io_connPE_50_push_ready,
	io_connPE_50_push_valid,
	io_connPE_50_push_bits,
	io_connPE_50_pop_ready,
	io_connPE_50_pop_valid,
	io_connPE_50_pop_bits,
	io_connPE_51_push_ready,
	io_connPE_51_push_valid,
	io_connPE_51_push_bits,
	io_connPE_51_pop_ready,
	io_connPE_51_pop_valid,
	io_connPE_51_pop_bits,
	io_connPE_52_push_ready,
	io_connPE_52_push_valid,
	io_connPE_52_push_bits,
	io_connPE_52_pop_ready,
	io_connPE_52_pop_valid,
	io_connPE_52_pop_bits,
	io_connPE_53_push_ready,
	io_connPE_53_push_valid,
	io_connPE_53_push_bits,
	io_connPE_53_pop_ready,
	io_connPE_53_pop_valid,
	io_connPE_53_pop_bits,
	io_connPE_54_push_ready,
	io_connPE_54_push_valid,
	io_connPE_54_push_bits,
	io_connPE_54_pop_ready,
	io_connPE_54_pop_valid,
	io_connPE_54_pop_bits,
	io_connPE_55_push_ready,
	io_connPE_55_push_valid,
	io_connPE_55_push_bits,
	io_connPE_55_pop_ready,
	io_connPE_55_pop_valid,
	io_connPE_55_pop_bits,
	io_connPE_56_push_ready,
	io_connPE_56_push_valid,
	io_connPE_56_push_bits,
	io_connPE_56_pop_ready,
	io_connPE_56_pop_valid,
	io_connPE_56_pop_bits,
	io_connPE_57_push_ready,
	io_connPE_57_push_valid,
	io_connPE_57_push_bits,
	io_connPE_57_pop_ready,
	io_connPE_57_pop_valid,
	io_connPE_57_pop_bits,
	io_connPE_58_push_ready,
	io_connPE_58_push_valid,
	io_connPE_58_push_bits,
	io_connPE_58_pop_ready,
	io_connPE_58_pop_valid,
	io_connPE_58_pop_bits,
	io_connPE_59_push_ready,
	io_connPE_59_push_valid,
	io_connPE_59_push_bits,
	io_connPE_59_pop_ready,
	io_connPE_59_pop_valid,
	io_connPE_59_pop_bits,
	io_connPE_60_push_ready,
	io_connPE_60_push_valid,
	io_connPE_60_push_bits,
	io_connPE_60_pop_ready,
	io_connPE_60_pop_valid,
	io_connPE_60_pop_bits,
	io_connPE_61_push_ready,
	io_connPE_61_push_valid,
	io_connPE_61_push_bits,
	io_connPE_61_pop_ready,
	io_connPE_61_pop_valid,
	io_connPE_61_pop_bits,
	io_connPE_62_push_ready,
	io_connPE_62_push_valid,
	io_connPE_62_push_bits,
	io_connPE_62_pop_ready,
	io_connPE_62_pop_valid,
	io_connPE_62_pop_bits,
	io_connPE_63_push_ready,
	io_connPE_63_push_valid,
	io_connPE_63_push_bits,
	io_connPE_63_pop_ready,
	io_connPE_63_pop_valid,
	io_connPE_63_pop_bits,
	io_connVSS_0_ctrl_serveStealReq_valid,
	io_connVSS_0_ctrl_serveStealReq_ready,
	io_connVSS_0_data_availableTask_ready,
	io_connVSS_0_data_availableTask_valid,
	io_connVSS_0_data_availableTask_bits,
	io_connVSS_0_data_qOutTask_ready,
	io_connVSS_0_data_qOutTask_valid,
	io_connVSS_0_data_qOutTask_bits,
	io_connVSS_1_ctrl_serveStealReq_valid,
	io_connVSS_1_ctrl_serveStealReq_ready,
	io_connVSS_1_data_availableTask_ready,
	io_connVSS_1_data_availableTask_valid,
	io_connVSS_1_data_availableTask_bits,
	io_connVSS_1_data_qOutTask_ready,
	io_connVSS_1_data_qOutTask_valid,
	io_connVSS_1_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0,
	io_ntwDataUnitOccupancyVSS_1
);
	input clock;
	input reset;
	output wire io_connPE_0_push_ready;
	input io_connPE_0_push_valid;
	input [127:0] io_connPE_0_push_bits;
	input io_connPE_0_pop_ready;
	output wire io_connPE_0_pop_valid;
	output wire [127:0] io_connPE_0_pop_bits;
	output wire io_connPE_1_push_ready;
	input io_connPE_1_push_valid;
	input [127:0] io_connPE_1_push_bits;
	input io_connPE_1_pop_ready;
	output wire io_connPE_1_pop_valid;
	output wire [127:0] io_connPE_1_pop_bits;
	output wire io_connPE_2_push_ready;
	input io_connPE_2_push_valid;
	input [127:0] io_connPE_2_push_bits;
	input io_connPE_2_pop_ready;
	output wire io_connPE_2_pop_valid;
	output wire [127:0] io_connPE_2_pop_bits;
	output wire io_connPE_3_push_ready;
	input io_connPE_3_push_valid;
	input [127:0] io_connPE_3_push_bits;
	input io_connPE_3_pop_ready;
	output wire io_connPE_3_pop_valid;
	output wire [127:0] io_connPE_3_pop_bits;
	output wire io_connPE_4_push_ready;
	input io_connPE_4_push_valid;
	input [127:0] io_connPE_4_push_bits;
	input io_connPE_4_pop_ready;
	output wire io_connPE_4_pop_valid;
	output wire [127:0] io_connPE_4_pop_bits;
	output wire io_connPE_5_push_ready;
	input io_connPE_5_push_valid;
	input [127:0] io_connPE_5_push_bits;
	input io_connPE_5_pop_ready;
	output wire io_connPE_5_pop_valid;
	output wire [127:0] io_connPE_5_pop_bits;
	output wire io_connPE_6_push_ready;
	input io_connPE_6_push_valid;
	input [127:0] io_connPE_6_push_bits;
	input io_connPE_6_pop_ready;
	output wire io_connPE_6_pop_valid;
	output wire [127:0] io_connPE_6_pop_bits;
	output wire io_connPE_7_push_ready;
	input io_connPE_7_push_valid;
	input [127:0] io_connPE_7_push_bits;
	input io_connPE_7_pop_ready;
	output wire io_connPE_7_pop_valid;
	output wire [127:0] io_connPE_7_pop_bits;
	output wire io_connPE_8_push_ready;
	input io_connPE_8_push_valid;
	input [127:0] io_connPE_8_push_bits;
	input io_connPE_8_pop_ready;
	output wire io_connPE_8_pop_valid;
	output wire [127:0] io_connPE_8_pop_bits;
	output wire io_connPE_9_push_ready;
	input io_connPE_9_push_valid;
	input [127:0] io_connPE_9_push_bits;
	input io_connPE_9_pop_ready;
	output wire io_connPE_9_pop_valid;
	output wire [127:0] io_connPE_9_pop_bits;
	output wire io_connPE_10_push_ready;
	input io_connPE_10_push_valid;
	input [127:0] io_connPE_10_push_bits;
	input io_connPE_10_pop_ready;
	output wire io_connPE_10_pop_valid;
	output wire [127:0] io_connPE_10_pop_bits;
	output wire io_connPE_11_push_ready;
	input io_connPE_11_push_valid;
	input [127:0] io_connPE_11_push_bits;
	input io_connPE_11_pop_ready;
	output wire io_connPE_11_pop_valid;
	output wire [127:0] io_connPE_11_pop_bits;
	output wire io_connPE_12_push_ready;
	input io_connPE_12_push_valid;
	input [127:0] io_connPE_12_push_bits;
	input io_connPE_12_pop_ready;
	output wire io_connPE_12_pop_valid;
	output wire [127:0] io_connPE_12_pop_bits;
	output wire io_connPE_13_push_ready;
	input io_connPE_13_push_valid;
	input [127:0] io_connPE_13_push_bits;
	input io_connPE_13_pop_ready;
	output wire io_connPE_13_pop_valid;
	output wire [127:0] io_connPE_13_pop_bits;
	output wire io_connPE_14_push_ready;
	input io_connPE_14_push_valid;
	input [127:0] io_connPE_14_push_bits;
	input io_connPE_14_pop_ready;
	output wire io_connPE_14_pop_valid;
	output wire [127:0] io_connPE_14_pop_bits;
	output wire io_connPE_15_push_ready;
	input io_connPE_15_push_valid;
	input [127:0] io_connPE_15_push_bits;
	input io_connPE_15_pop_ready;
	output wire io_connPE_15_pop_valid;
	output wire [127:0] io_connPE_15_pop_bits;
	output wire io_connPE_16_push_ready;
	input io_connPE_16_push_valid;
	input [127:0] io_connPE_16_push_bits;
	input io_connPE_16_pop_ready;
	output wire io_connPE_16_pop_valid;
	output wire [127:0] io_connPE_16_pop_bits;
	output wire io_connPE_17_push_ready;
	input io_connPE_17_push_valid;
	input [127:0] io_connPE_17_push_bits;
	input io_connPE_17_pop_ready;
	output wire io_connPE_17_pop_valid;
	output wire [127:0] io_connPE_17_pop_bits;
	output wire io_connPE_18_push_ready;
	input io_connPE_18_push_valid;
	input [127:0] io_connPE_18_push_bits;
	input io_connPE_18_pop_ready;
	output wire io_connPE_18_pop_valid;
	output wire [127:0] io_connPE_18_pop_bits;
	output wire io_connPE_19_push_ready;
	input io_connPE_19_push_valid;
	input [127:0] io_connPE_19_push_bits;
	input io_connPE_19_pop_ready;
	output wire io_connPE_19_pop_valid;
	output wire [127:0] io_connPE_19_pop_bits;
	output wire io_connPE_20_push_ready;
	input io_connPE_20_push_valid;
	input [127:0] io_connPE_20_push_bits;
	input io_connPE_20_pop_ready;
	output wire io_connPE_20_pop_valid;
	output wire [127:0] io_connPE_20_pop_bits;
	output wire io_connPE_21_push_ready;
	input io_connPE_21_push_valid;
	input [127:0] io_connPE_21_push_bits;
	input io_connPE_21_pop_ready;
	output wire io_connPE_21_pop_valid;
	output wire [127:0] io_connPE_21_pop_bits;
	output wire io_connPE_22_push_ready;
	input io_connPE_22_push_valid;
	input [127:0] io_connPE_22_push_bits;
	input io_connPE_22_pop_ready;
	output wire io_connPE_22_pop_valid;
	output wire [127:0] io_connPE_22_pop_bits;
	output wire io_connPE_23_push_ready;
	input io_connPE_23_push_valid;
	input [127:0] io_connPE_23_push_bits;
	input io_connPE_23_pop_ready;
	output wire io_connPE_23_pop_valid;
	output wire [127:0] io_connPE_23_pop_bits;
	output wire io_connPE_24_push_ready;
	input io_connPE_24_push_valid;
	input [127:0] io_connPE_24_push_bits;
	input io_connPE_24_pop_ready;
	output wire io_connPE_24_pop_valid;
	output wire [127:0] io_connPE_24_pop_bits;
	output wire io_connPE_25_push_ready;
	input io_connPE_25_push_valid;
	input [127:0] io_connPE_25_push_bits;
	input io_connPE_25_pop_ready;
	output wire io_connPE_25_pop_valid;
	output wire [127:0] io_connPE_25_pop_bits;
	output wire io_connPE_26_push_ready;
	input io_connPE_26_push_valid;
	input [127:0] io_connPE_26_push_bits;
	input io_connPE_26_pop_ready;
	output wire io_connPE_26_pop_valid;
	output wire [127:0] io_connPE_26_pop_bits;
	output wire io_connPE_27_push_ready;
	input io_connPE_27_push_valid;
	input [127:0] io_connPE_27_push_bits;
	input io_connPE_27_pop_ready;
	output wire io_connPE_27_pop_valid;
	output wire [127:0] io_connPE_27_pop_bits;
	output wire io_connPE_28_push_ready;
	input io_connPE_28_push_valid;
	input [127:0] io_connPE_28_push_bits;
	input io_connPE_28_pop_ready;
	output wire io_connPE_28_pop_valid;
	output wire [127:0] io_connPE_28_pop_bits;
	output wire io_connPE_29_push_ready;
	input io_connPE_29_push_valid;
	input [127:0] io_connPE_29_push_bits;
	input io_connPE_29_pop_ready;
	output wire io_connPE_29_pop_valid;
	output wire [127:0] io_connPE_29_pop_bits;
	output wire io_connPE_30_push_ready;
	input io_connPE_30_push_valid;
	input [127:0] io_connPE_30_push_bits;
	input io_connPE_30_pop_ready;
	output wire io_connPE_30_pop_valid;
	output wire [127:0] io_connPE_30_pop_bits;
	output wire io_connPE_31_push_ready;
	input io_connPE_31_push_valid;
	input [127:0] io_connPE_31_push_bits;
	input io_connPE_31_pop_ready;
	output wire io_connPE_31_pop_valid;
	output wire [127:0] io_connPE_31_pop_bits;
	output wire io_connPE_32_push_ready;
	input io_connPE_32_push_valid;
	input [127:0] io_connPE_32_push_bits;
	input io_connPE_32_pop_ready;
	output wire io_connPE_32_pop_valid;
	output wire [127:0] io_connPE_32_pop_bits;
	output wire io_connPE_33_push_ready;
	input io_connPE_33_push_valid;
	input [127:0] io_connPE_33_push_bits;
	input io_connPE_33_pop_ready;
	output wire io_connPE_33_pop_valid;
	output wire [127:0] io_connPE_33_pop_bits;
	output wire io_connPE_34_push_ready;
	input io_connPE_34_push_valid;
	input [127:0] io_connPE_34_push_bits;
	input io_connPE_34_pop_ready;
	output wire io_connPE_34_pop_valid;
	output wire [127:0] io_connPE_34_pop_bits;
	output wire io_connPE_35_push_ready;
	input io_connPE_35_push_valid;
	input [127:0] io_connPE_35_push_bits;
	input io_connPE_35_pop_ready;
	output wire io_connPE_35_pop_valid;
	output wire [127:0] io_connPE_35_pop_bits;
	output wire io_connPE_36_push_ready;
	input io_connPE_36_push_valid;
	input [127:0] io_connPE_36_push_bits;
	input io_connPE_36_pop_ready;
	output wire io_connPE_36_pop_valid;
	output wire [127:0] io_connPE_36_pop_bits;
	output wire io_connPE_37_push_ready;
	input io_connPE_37_push_valid;
	input [127:0] io_connPE_37_push_bits;
	input io_connPE_37_pop_ready;
	output wire io_connPE_37_pop_valid;
	output wire [127:0] io_connPE_37_pop_bits;
	output wire io_connPE_38_push_ready;
	input io_connPE_38_push_valid;
	input [127:0] io_connPE_38_push_bits;
	input io_connPE_38_pop_ready;
	output wire io_connPE_38_pop_valid;
	output wire [127:0] io_connPE_38_pop_bits;
	output wire io_connPE_39_push_ready;
	input io_connPE_39_push_valid;
	input [127:0] io_connPE_39_push_bits;
	input io_connPE_39_pop_ready;
	output wire io_connPE_39_pop_valid;
	output wire [127:0] io_connPE_39_pop_bits;
	output wire io_connPE_40_push_ready;
	input io_connPE_40_push_valid;
	input [127:0] io_connPE_40_push_bits;
	input io_connPE_40_pop_ready;
	output wire io_connPE_40_pop_valid;
	output wire [127:0] io_connPE_40_pop_bits;
	output wire io_connPE_41_push_ready;
	input io_connPE_41_push_valid;
	input [127:0] io_connPE_41_push_bits;
	input io_connPE_41_pop_ready;
	output wire io_connPE_41_pop_valid;
	output wire [127:0] io_connPE_41_pop_bits;
	output wire io_connPE_42_push_ready;
	input io_connPE_42_push_valid;
	input [127:0] io_connPE_42_push_bits;
	input io_connPE_42_pop_ready;
	output wire io_connPE_42_pop_valid;
	output wire [127:0] io_connPE_42_pop_bits;
	output wire io_connPE_43_push_ready;
	input io_connPE_43_push_valid;
	input [127:0] io_connPE_43_push_bits;
	input io_connPE_43_pop_ready;
	output wire io_connPE_43_pop_valid;
	output wire [127:0] io_connPE_43_pop_bits;
	output wire io_connPE_44_push_ready;
	input io_connPE_44_push_valid;
	input [127:0] io_connPE_44_push_bits;
	input io_connPE_44_pop_ready;
	output wire io_connPE_44_pop_valid;
	output wire [127:0] io_connPE_44_pop_bits;
	output wire io_connPE_45_push_ready;
	input io_connPE_45_push_valid;
	input [127:0] io_connPE_45_push_bits;
	input io_connPE_45_pop_ready;
	output wire io_connPE_45_pop_valid;
	output wire [127:0] io_connPE_45_pop_bits;
	output wire io_connPE_46_push_ready;
	input io_connPE_46_push_valid;
	input [127:0] io_connPE_46_push_bits;
	input io_connPE_46_pop_ready;
	output wire io_connPE_46_pop_valid;
	output wire [127:0] io_connPE_46_pop_bits;
	output wire io_connPE_47_push_ready;
	input io_connPE_47_push_valid;
	input [127:0] io_connPE_47_push_bits;
	input io_connPE_47_pop_ready;
	output wire io_connPE_47_pop_valid;
	output wire [127:0] io_connPE_47_pop_bits;
	output wire io_connPE_48_push_ready;
	input io_connPE_48_push_valid;
	input [127:0] io_connPE_48_push_bits;
	input io_connPE_48_pop_ready;
	output wire io_connPE_48_pop_valid;
	output wire [127:0] io_connPE_48_pop_bits;
	output wire io_connPE_49_push_ready;
	input io_connPE_49_push_valid;
	input [127:0] io_connPE_49_push_bits;
	input io_connPE_49_pop_ready;
	output wire io_connPE_49_pop_valid;
	output wire [127:0] io_connPE_49_pop_bits;
	output wire io_connPE_50_push_ready;
	input io_connPE_50_push_valid;
	input [127:0] io_connPE_50_push_bits;
	input io_connPE_50_pop_ready;
	output wire io_connPE_50_pop_valid;
	output wire [127:0] io_connPE_50_pop_bits;
	output wire io_connPE_51_push_ready;
	input io_connPE_51_push_valid;
	input [127:0] io_connPE_51_push_bits;
	input io_connPE_51_pop_ready;
	output wire io_connPE_51_pop_valid;
	output wire [127:0] io_connPE_51_pop_bits;
	output wire io_connPE_52_push_ready;
	input io_connPE_52_push_valid;
	input [127:0] io_connPE_52_push_bits;
	input io_connPE_52_pop_ready;
	output wire io_connPE_52_pop_valid;
	output wire [127:0] io_connPE_52_pop_bits;
	output wire io_connPE_53_push_ready;
	input io_connPE_53_push_valid;
	input [127:0] io_connPE_53_push_bits;
	input io_connPE_53_pop_ready;
	output wire io_connPE_53_pop_valid;
	output wire [127:0] io_connPE_53_pop_bits;
	output wire io_connPE_54_push_ready;
	input io_connPE_54_push_valid;
	input [127:0] io_connPE_54_push_bits;
	input io_connPE_54_pop_ready;
	output wire io_connPE_54_pop_valid;
	output wire [127:0] io_connPE_54_pop_bits;
	output wire io_connPE_55_push_ready;
	input io_connPE_55_push_valid;
	input [127:0] io_connPE_55_push_bits;
	input io_connPE_55_pop_ready;
	output wire io_connPE_55_pop_valid;
	output wire [127:0] io_connPE_55_pop_bits;
	output wire io_connPE_56_push_ready;
	input io_connPE_56_push_valid;
	input [127:0] io_connPE_56_push_bits;
	input io_connPE_56_pop_ready;
	output wire io_connPE_56_pop_valid;
	output wire [127:0] io_connPE_56_pop_bits;
	output wire io_connPE_57_push_ready;
	input io_connPE_57_push_valid;
	input [127:0] io_connPE_57_push_bits;
	input io_connPE_57_pop_ready;
	output wire io_connPE_57_pop_valid;
	output wire [127:0] io_connPE_57_pop_bits;
	output wire io_connPE_58_push_ready;
	input io_connPE_58_push_valid;
	input [127:0] io_connPE_58_push_bits;
	input io_connPE_58_pop_ready;
	output wire io_connPE_58_pop_valid;
	output wire [127:0] io_connPE_58_pop_bits;
	output wire io_connPE_59_push_ready;
	input io_connPE_59_push_valid;
	input [127:0] io_connPE_59_push_bits;
	input io_connPE_59_pop_ready;
	output wire io_connPE_59_pop_valid;
	output wire [127:0] io_connPE_59_pop_bits;
	output wire io_connPE_60_push_ready;
	input io_connPE_60_push_valid;
	input [127:0] io_connPE_60_push_bits;
	input io_connPE_60_pop_ready;
	output wire io_connPE_60_pop_valid;
	output wire [127:0] io_connPE_60_pop_bits;
	output wire io_connPE_61_push_ready;
	input io_connPE_61_push_valid;
	input [127:0] io_connPE_61_push_bits;
	input io_connPE_61_pop_ready;
	output wire io_connPE_61_pop_valid;
	output wire [127:0] io_connPE_61_pop_bits;
	output wire io_connPE_62_push_ready;
	input io_connPE_62_push_valid;
	input [127:0] io_connPE_62_push_bits;
	input io_connPE_62_pop_ready;
	output wire io_connPE_62_pop_valid;
	output wire [127:0] io_connPE_62_pop_bits;
	output wire io_connPE_63_push_ready;
	input io_connPE_63_push_valid;
	input [127:0] io_connPE_63_push_bits;
	input io_connPE_63_pop_ready;
	output wire io_connPE_63_pop_valid;
	output wire [127:0] io_connPE_63_pop_bits;
	input io_connVSS_0_ctrl_serveStealReq_valid;
	output wire io_connVSS_0_ctrl_serveStealReq_ready;
	input io_connVSS_0_data_availableTask_ready;
	output wire io_connVSS_0_data_availableTask_valid;
	output wire [127:0] io_connVSS_0_data_availableTask_bits;
	output wire io_connVSS_0_data_qOutTask_ready;
	input io_connVSS_0_data_qOutTask_valid;
	input [127:0] io_connVSS_0_data_qOutTask_bits;
	input io_connVSS_1_ctrl_serveStealReq_valid;
	output wire io_connVSS_1_ctrl_serveStealReq_ready;
	input io_connVSS_1_data_availableTask_ready;
	output wire io_connVSS_1_data_availableTask_valid;
	output wire [127:0] io_connVSS_1_data_availableTask_bits;
	output wire io_connVSS_1_data_qOutTask_ready;
	input io_connVSS_1_data_qOutTask_valid;
	input [127:0] io_connVSS_1_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	output wire io_ntwDataUnitOccupancyVSS_1;
	wire [4:0] _taskQueues_63_io_connVec_1_currLength;
	wire _taskQueues_63_io_connVec_1_push_ready;
	wire _taskQueues_63_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_63_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_62_io_connVec_1_currLength;
	wire _taskQueues_62_io_connVec_1_push_ready;
	wire _taskQueues_62_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_62_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_61_io_connVec_1_currLength;
	wire _taskQueues_61_io_connVec_1_push_ready;
	wire _taskQueues_61_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_61_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_60_io_connVec_1_currLength;
	wire _taskQueues_60_io_connVec_1_push_ready;
	wire _taskQueues_60_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_60_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_59_io_connVec_1_currLength;
	wire _taskQueues_59_io_connVec_1_push_ready;
	wire _taskQueues_59_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_59_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_58_io_connVec_1_currLength;
	wire _taskQueues_58_io_connVec_1_push_ready;
	wire _taskQueues_58_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_58_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_57_io_connVec_1_currLength;
	wire _taskQueues_57_io_connVec_1_push_ready;
	wire _taskQueues_57_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_57_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_56_io_connVec_1_currLength;
	wire _taskQueues_56_io_connVec_1_push_ready;
	wire _taskQueues_56_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_56_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_55_io_connVec_1_currLength;
	wire _taskQueues_55_io_connVec_1_push_ready;
	wire _taskQueues_55_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_55_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_54_io_connVec_1_currLength;
	wire _taskQueues_54_io_connVec_1_push_ready;
	wire _taskQueues_54_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_54_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_53_io_connVec_1_currLength;
	wire _taskQueues_53_io_connVec_1_push_ready;
	wire _taskQueues_53_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_53_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_52_io_connVec_1_currLength;
	wire _taskQueues_52_io_connVec_1_push_ready;
	wire _taskQueues_52_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_52_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_51_io_connVec_1_currLength;
	wire _taskQueues_51_io_connVec_1_push_ready;
	wire _taskQueues_51_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_51_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_50_io_connVec_1_currLength;
	wire _taskQueues_50_io_connVec_1_push_ready;
	wire _taskQueues_50_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_50_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_49_io_connVec_1_currLength;
	wire _taskQueues_49_io_connVec_1_push_ready;
	wire _taskQueues_49_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_49_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_48_io_connVec_1_currLength;
	wire _taskQueues_48_io_connVec_1_push_ready;
	wire _taskQueues_48_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_48_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_47_io_connVec_1_currLength;
	wire _taskQueues_47_io_connVec_1_push_ready;
	wire _taskQueues_47_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_47_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_46_io_connVec_1_currLength;
	wire _taskQueues_46_io_connVec_1_push_ready;
	wire _taskQueues_46_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_46_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_45_io_connVec_1_currLength;
	wire _taskQueues_45_io_connVec_1_push_ready;
	wire _taskQueues_45_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_45_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_44_io_connVec_1_currLength;
	wire _taskQueues_44_io_connVec_1_push_ready;
	wire _taskQueues_44_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_44_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_43_io_connVec_1_currLength;
	wire _taskQueues_43_io_connVec_1_push_ready;
	wire _taskQueues_43_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_43_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_42_io_connVec_1_currLength;
	wire _taskQueues_42_io_connVec_1_push_ready;
	wire _taskQueues_42_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_42_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_41_io_connVec_1_currLength;
	wire _taskQueues_41_io_connVec_1_push_ready;
	wire _taskQueues_41_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_41_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_40_io_connVec_1_currLength;
	wire _taskQueues_40_io_connVec_1_push_ready;
	wire _taskQueues_40_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_40_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_39_io_connVec_1_currLength;
	wire _taskQueues_39_io_connVec_1_push_ready;
	wire _taskQueues_39_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_39_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_38_io_connVec_1_currLength;
	wire _taskQueues_38_io_connVec_1_push_ready;
	wire _taskQueues_38_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_38_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_37_io_connVec_1_currLength;
	wire _taskQueues_37_io_connVec_1_push_ready;
	wire _taskQueues_37_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_37_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_36_io_connVec_1_currLength;
	wire _taskQueues_36_io_connVec_1_push_ready;
	wire _taskQueues_36_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_36_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_35_io_connVec_1_currLength;
	wire _taskQueues_35_io_connVec_1_push_ready;
	wire _taskQueues_35_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_35_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_34_io_connVec_1_currLength;
	wire _taskQueues_34_io_connVec_1_push_ready;
	wire _taskQueues_34_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_34_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_33_io_connVec_1_currLength;
	wire _taskQueues_33_io_connVec_1_push_ready;
	wire _taskQueues_33_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_33_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_32_io_connVec_1_currLength;
	wire _taskQueues_32_io_connVec_1_push_ready;
	wire _taskQueues_32_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_32_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_31_io_connVec_1_currLength;
	wire _taskQueues_31_io_connVec_1_push_ready;
	wire _taskQueues_31_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_31_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_30_io_connVec_1_currLength;
	wire _taskQueues_30_io_connVec_1_push_ready;
	wire _taskQueues_30_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_30_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_29_io_connVec_1_currLength;
	wire _taskQueues_29_io_connVec_1_push_ready;
	wire _taskQueues_29_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_29_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_28_io_connVec_1_currLength;
	wire _taskQueues_28_io_connVec_1_push_ready;
	wire _taskQueues_28_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_28_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_27_io_connVec_1_currLength;
	wire _taskQueues_27_io_connVec_1_push_ready;
	wire _taskQueues_27_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_27_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_26_io_connVec_1_currLength;
	wire _taskQueues_26_io_connVec_1_push_ready;
	wire _taskQueues_26_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_26_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_25_io_connVec_1_currLength;
	wire _taskQueues_25_io_connVec_1_push_ready;
	wire _taskQueues_25_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_25_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_24_io_connVec_1_currLength;
	wire _taskQueues_24_io_connVec_1_push_ready;
	wire _taskQueues_24_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_24_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_23_io_connVec_1_currLength;
	wire _taskQueues_23_io_connVec_1_push_ready;
	wire _taskQueues_23_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_23_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_22_io_connVec_1_currLength;
	wire _taskQueues_22_io_connVec_1_push_ready;
	wire _taskQueues_22_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_22_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_21_io_connVec_1_currLength;
	wire _taskQueues_21_io_connVec_1_push_ready;
	wire _taskQueues_21_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_21_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_20_io_connVec_1_currLength;
	wire _taskQueues_20_io_connVec_1_push_ready;
	wire _taskQueues_20_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_20_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_19_io_connVec_1_currLength;
	wire _taskQueues_19_io_connVec_1_push_ready;
	wire _taskQueues_19_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_19_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_18_io_connVec_1_currLength;
	wire _taskQueues_18_io_connVec_1_push_ready;
	wire _taskQueues_18_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_18_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_17_io_connVec_1_currLength;
	wire _taskQueues_17_io_connVec_1_push_ready;
	wire _taskQueues_17_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_17_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_16_io_connVec_1_currLength;
	wire _taskQueues_16_io_connVec_1_push_ready;
	wire _taskQueues_16_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_16_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_15_io_connVec_1_currLength;
	wire _taskQueues_15_io_connVec_1_push_ready;
	wire _taskQueues_15_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_15_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_14_io_connVec_1_currLength;
	wire _taskQueues_14_io_connVec_1_push_ready;
	wire _taskQueues_14_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_14_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_13_io_connVec_1_currLength;
	wire _taskQueues_13_io_connVec_1_push_ready;
	wire _taskQueues_13_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_13_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_12_io_connVec_1_currLength;
	wire _taskQueues_12_io_connVec_1_push_ready;
	wire _taskQueues_12_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_12_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_11_io_connVec_1_currLength;
	wire _taskQueues_11_io_connVec_1_push_ready;
	wire _taskQueues_11_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_11_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_10_io_connVec_1_currLength;
	wire _taskQueues_10_io_connVec_1_push_ready;
	wire _taskQueues_10_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_10_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_9_io_connVec_1_currLength;
	wire _taskQueues_9_io_connVec_1_push_ready;
	wire _taskQueues_9_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_9_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_8_io_connVec_1_currLength;
	wire _taskQueues_8_io_connVec_1_push_ready;
	wire _taskQueues_8_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_8_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_7_io_connVec_1_currLength;
	wire _taskQueues_7_io_connVec_1_push_ready;
	wire _taskQueues_7_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_7_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_6_io_connVec_1_currLength;
	wire _taskQueues_6_io_connVec_1_push_ready;
	wire _taskQueues_6_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_6_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_5_io_connVec_1_currLength;
	wire _taskQueues_5_io_connVec_1_push_ready;
	wire _taskQueues_5_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_5_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_4_io_connVec_1_currLength;
	wire _taskQueues_4_io_connVec_1_push_ready;
	wire _taskQueues_4_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_4_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_3_io_connVec_1_currLength;
	wire _taskQueues_3_io_connVec_1_push_ready;
	wire _taskQueues_3_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_3_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_2_io_connVec_1_currLength;
	wire _taskQueues_2_io_connVec_1_push_ready;
	wire _taskQueues_2_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_2_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_1_io_connVec_1_currLength;
	wire _taskQueues_1_io_connVec_1_push_ready;
	wire _taskQueues_1_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_1_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_0_io_connVec_1_currLength;
	wire _taskQueues_0_io_connVec_1_push_ready;
	wire _taskQueues_0_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_0_io_connVec_1_pop_bits;
	wire _stealServers_63_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_63_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_63_io_connNetwork_data_availableTask_ready;
	wire _stealServers_63_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_63_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_63_io_connQ_push_valid;
	wire [127:0] _stealServers_63_io_connQ_push_bits;
	wire _stealServers_63_io_connQ_pop_ready;
	wire _stealServers_62_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_62_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_62_io_connNetwork_data_availableTask_ready;
	wire _stealServers_62_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_62_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_62_io_connQ_push_valid;
	wire [127:0] _stealServers_62_io_connQ_push_bits;
	wire _stealServers_62_io_connQ_pop_ready;
	wire _stealServers_61_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_61_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_61_io_connNetwork_data_availableTask_ready;
	wire _stealServers_61_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_61_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_61_io_connQ_push_valid;
	wire [127:0] _stealServers_61_io_connQ_push_bits;
	wire _stealServers_61_io_connQ_pop_ready;
	wire _stealServers_60_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_60_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_60_io_connNetwork_data_availableTask_ready;
	wire _stealServers_60_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_60_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_60_io_connQ_push_valid;
	wire [127:0] _stealServers_60_io_connQ_push_bits;
	wire _stealServers_60_io_connQ_pop_ready;
	wire _stealServers_59_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_59_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_59_io_connNetwork_data_availableTask_ready;
	wire _stealServers_59_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_59_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_59_io_connQ_push_valid;
	wire [127:0] _stealServers_59_io_connQ_push_bits;
	wire _stealServers_59_io_connQ_pop_ready;
	wire _stealServers_58_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_58_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_58_io_connNetwork_data_availableTask_ready;
	wire _stealServers_58_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_58_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_58_io_connQ_push_valid;
	wire [127:0] _stealServers_58_io_connQ_push_bits;
	wire _stealServers_58_io_connQ_pop_ready;
	wire _stealServers_57_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_57_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_57_io_connNetwork_data_availableTask_ready;
	wire _stealServers_57_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_57_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_57_io_connQ_push_valid;
	wire [127:0] _stealServers_57_io_connQ_push_bits;
	wire _stealServers_57_io_connQ_pop_ready;
	wire _stealServers_56_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_56_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_56_io_connNetwork_data_availableTask_ready;
	wire _stealServers_56_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_56_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_56_io_connQ_push_valid;
	wire [127:0] _stealServers_56_io_connQ_push_bits;
	wire _stealServers_56_io_connQ_pop_ready;
	wire _stealServers_55_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_55_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_55_io_connNetwork_data_availableTask_ready;
	wire _stealServers_55_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_55_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_55_io_connQ_push_valid;
	wire [127:0] _stealServers_55_io_connQ_push_bits;
	wire _stealServers_55_io_connQ_pop_ready;
	wire _stealServers_54_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_54_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_54_io_connNetwork_data_availableTask_ready;
	wire _stealServers_54_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_54_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_54_io_connQ_push_valid;
	wire [127:0] _stealServers_54_io_connQ_push_bits;
	wire _stealServers_54_io_connQ_pop_ready;
	wire _stealServers_53_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_53_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_53_io_connNetwork_data_availableTask_ready;
	wire _stealServers_53_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_53_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_53_io_connQ_push_valid;
	wire [127:0] _stealServers_53_io_connQ_push_bits;
	wire _stealServers_53_io_connQ_pop_ready;
	wire _stealServers_52_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_52_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_52_io_connNetwork_data_availableTask_ready;
	wire _stealServers_52_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_52_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_52_io_connQ_push_valid;
	wire [127:0] _stealServers_52_io_connQ_push_bits;
	wire _stealServers_52_io_connQ_pop_ready;
	wire _stealServers_51_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_51_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_51_io_connNetwork_data_availableTask_ready;
	wire _stealServers_51_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_51_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_51_io_connQ_push_valid;
	wire [127:0] _stealServers_51_io_connQ_push_bits;
	wire _stealServers_51_io_connQ_pop_ready;
	wire _stealServers_50_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_50_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_50_io_connNetwork_data_availableTask_ready;
	wire _stealServers_50_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_50_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_50_io_connQ_push_valid;
	wire [127:0] _stealServers_50_io_connQ_push_bits;
	wire _stealServers_50_io_connQ_pop_ready;
	wire _stealServers_49_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_49_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_49_io_connNetwork_data_availableTask_ready;
	wire _stealServers_49_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_49_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_49_io_connQ_push_valid;
	wire [127:0] _stealServers_49_io_connQ_push_bits;
	wire _stealServers_49_io_connQ_pop_ready;
	wire _stealServers_48_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_48_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_48_io_connNetwork_data_availableTask_ready;
	wire _stealServers_48_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_48_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_48_io_connQ_push_valid;
	wire [127:0] _stealServers_48_io_connQ_push_bits;
	wire _stealServers_48_io_connQ_pop_ready;
	wire _stealServers_47_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_47_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_47_io_connNetwork_data_availableTask_ready;
	wire _stealServers_47_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_47_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_47_io_connQ_push_valid;
	wire [127:0] _stealServers_47_io_connQ_push_bits;
	wire _stealServers_47_io_connQ_pop_ready;
	wire _stealServers_46_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_46_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_46_io_connNetwork_data_availableTask_ready;
	wire _stealServers_46_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_46_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_46_io_connQ_push_valid;
	wire [127:0] _stealServers_46_io_connQ_push_bits;
	wire _stealServers_46_io_connQ_pop_ready;
	wire _stealServers_45_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_45_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_45_io_connNetwork_data_availableTask_ready;
	wire _stealServers_45_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_45_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_45_io_connQ_push_valid;
	wire [127:0] _stealServers_45_io_connQ_push_bits;
	wire _stealServers_45_io_connQ_pop_ready;
	wire _stealServers_44_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_44_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_44_io_connNetwork_data_availableTask_ready;
	wire _stealServers_44_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_44_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_44_io_connQ_push_valid;
	wire [127:0] _stealServers_44_io_connQ_push_bits;
	wire _stealServers_44_io_connQ_pop_ready;
	wire _stealServers_43_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_43_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_43_io_connNetwork_data_availableTask_ready;
	wire _stealServers_43_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_43_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_43_io_connQ_push_valid;
	wire [127:0] _stealServers_43_io_connQ_push_bits;
	wire _stealServers_43_io_connQ_pop_ready;
	wire _stealServers_42_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_42_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_42_io_connNetwork_data_availableTask_ready;
	wire _stealServers_42_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_42_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_42_io_connQ_push_valid;
	wire [127:0] _stealServers_42_io_connQ_push_bits;
	wire _stealServers_42_io_connQ_pop_ready;
	wire _stealServers_41_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_41_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_41_io_connNetwork_data_availableTask_ready;
	wire _stealServers_41_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_41_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_41_io_connQ_push_valid;
	wire [127:0] _stealServers_41_io_connQ_push_bits;
	wire _stealServers_41_io_connQ_pop_ready;
	wire _stealServers_40_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_40_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_40_io_connNetwork_data_availableTask_ready;
	wire _stealServers_40_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_40_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_40_io_connQ_push_valid;
	wire [127:0] _stealServers_40_io_connQ_push_bits;
	wire _stealServers_40_io_connQ_pop_ready;
	wire _stealServers_39_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_39_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_39_io_connNetwork_data_availableTask_ready;
	wire _stealServers_39_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_39_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_39_io_connQ_push_valid;
	wire [127:0] _stealServers_39_io_connQ_push_bits;
	wire _stealServers_39_io_connQ_pop_ready;
	wire _stealServers_38_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_38_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_38_io_connNetwork_data_availableTask_ready;
	wire _stealServers_38_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_38_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_38_io_connQ_push_valid;
	wire [127:0] _stealServers_38_io_connQ_push_bits;
	wire _stealServers_38_io_connQ_pop_ready;
	wire _stealServers_37_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_37_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_37_io_connNetwork_data_availableTask_ready;
	wire _stealServers_37_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_37_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_37_io_connQ_push_valid;
	wire [127:0] _stealServers_37_io_connQ_push_bits;
	wire _stealServers_37_io_connQ_pop_ready;
	wire _stealServers_36_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_36_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_36_io_connNetwork_data_availableTask_ready;
	wire _stealServers_36_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_36_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_36_io_connQ_push_valid;
	wire [127:0] _stealServers_36_io_connQ_push_bits;
	wire _stealServers_36_io_connQ_pop_ready;
	wire _stealServers_35_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_35_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_35_io_connNetwork_data_availableTask_ready;
	wire _stealServers_35_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_35_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_35_io_connQ_push_valid;
	wire [127:0] _stealServers_35_io_connQ_push_bits;
	wire _stealServers_35_io_connQ_pop_ready;
	wire _stealServers_34_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_34_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_34_io_connNetwork_data_availableTask_ready;
	wire _stealServers_34_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_34_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_34_io_connQ_push_valid;
	wire [127:0] _stealServers_34_io_connQ_push_bits;
	wire _stealServers_34_io_connQ_pop_ready;
	wire _stealServers_33_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_33_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_33_io_connNetwork_data_availableTask_ready;
	wire _stealServers_33_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_33_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_33_io_connQ_push_valid;
	wire [127:0] _stealServers_33_io_connQ_push_bits;
	wire _stealServers_33_io_connQ_pop_ready;
	wire _stealServers_32_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_32_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_32_io_connNetwork_data_availableTask_ready;
	wire _stealServers_32_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_32_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_32_io_connQ_push_valid;
	wire [127:0] _stealServers_32_io_connQ_push_bits;
	wire _stealServers_32_io_connQ_pop_ready;
	wire _stealServers_31_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_31_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_31_io_connNetwork_data_availableTask_ready;
	wire _stealServers_31_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_31_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_31_io_connQ_push_valid;
	wire [127:0] _stealServers_31_io_connQ_push_bits;
	wire _stealServers_31_io_connQ_pop_ready;
	wire _stealServers_30_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_30_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_30_io_connNetwork_data_availableTask_ready;
	wire _stealServers_30_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_30_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_30_io_connQ_push_valid;
	wire [127:0] _stealServers_30_io_connQ_push_bits;
	wire _stealServers_30_io_connQ_pop_ready;
	wire _stealServers_29_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_29_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_29_io_connNetwork_data_availableTask_ready;
	wire _stealServers_29_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_29_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_29_io_connQ_push_valid;
	wire [127:0] _stealServers_29_io_connQ_push_bits;
	wire _stealServers_29_io_connQ_pop_ready;
	wire _stealServers_28_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_28_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_28_io_connNetwork_data_availableTask_ready;
	wire _stealServers_28_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_28_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_28_io_connQ_push_valid;
	wire [127:0] _stealServers_28_io_connQ_push_bits;
	wire _stealServers_28_io_connQ_pop_ready;
	wire _stealServers_27_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_27_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_27_io_connNetwork_data_availableTask_ready;
	wire _stealServers_27_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_27_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_27_io_connQ_push_valid;
	wire [127:0] _stealServers_27_io_connQ_push_bits;
	wire _stealServers_27_io_connQ_pop_ready;
	wire _stealServers_26_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_26_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_26_io_connNetwork_data_availableTask_ready;
	wire _stealServers_26_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_26_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_26_io_connQ_push_valid;
	wire [127:0] _stealServers_26_io_connQ_push_bits;
	wire _stealServers_26_io_connQ_pop_ready;
	wire _stealServers_25_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_25_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_25_io_connNetwork_data_availableTask_ready;
	wire _stealServers_25_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_25_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_25_io_connQ_push_valid;
	wire [127:0] _stealServers_25_io_connQ_push_bits;
	wire _stealServers_25_io_connQ_pop_ready;
	wire _stealServers_24_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_24_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_24_io_connNetwork_data_availableTask_ready;
	wire _stealServers_24_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_24_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_24_io_connQ_push_valid;
	wire [127:0] _stealServers_24_io_connQ_push_bits;
	wire _stealServers_24_io_connQ_pop_ready;
	wire _stealServers_23_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_23_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_23_io_connNetwork_data_availableTask_ready;
	wire _stealServers_23_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_23_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_23_io_connQ_push_valid;
	wire [127:0] _stealServers_23_io_connQ_push_bits;
	wire _stealServers_23_io_connQ_pop_ready;
	wire _stealServers_22_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_22_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_22_io_connNetwork_data_availableTask_ready;
	wire _stealServers_22_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_22_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_22_io_connQ_push_valid;
	wire [127:0] _stealServers_22_io_connQ_push_bits;
	wire _stealServers_22_io_connQ_pop_ready;
	wire _stealServers_21_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_21_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_21_io_connNetwork_data_availableTask_ready;
	wire _stealServers_21_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_21_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_21_io_connQ_push_valid;
	wire [127:0] _stealServers_21_io_connQ_push_bits;
	wire _stealServers_21_io_connQ_pop_ready;
	wire _stealServers_20_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_20_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_20_io_connNetwork_data_availableTask_ready;
	wire _stealServers_20_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_20_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_20_io_connQ_push_valid;
	wire [127:0] _stealServers_20_io_connQ_push_bits;
	wire _stealServers_20_io_connQ_pop_ready;
	wire _stealServers_19_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_19_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_19_io_connNetwork_data_availableTask_ready;
	wire _stealServers_19_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_19_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_19_io_connQ_push_valid;
	wire [127:0] _stealServers_19_io_connQ_push_bits;
	wire _stealServers_19_io_connQ_pop_ready;
	wire _stealServers_18_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_18_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_18_io_connNetwork_data_availableTask_ready;
	wire _stealServers_18_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_18_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_18_io_connQ_push_valid;
	wire [127:0] _stealServers_18_io_connQ_push_bits;
	wire _stealServers_18_io_connQ_pop_ready;
	wire _stealServers_17_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_17_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_17_io_connNetwork_data_availableTask_ready;
	wire _stealServers_17_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_17_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_17_io_connQ_push_valid;
	wire [127:0] _stealServers_17_io_connQ_push_bits;
	wire _stealServers_17_io_connQ_pop_ready;
	wire _stealServers_16_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_16_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_16_io_connNetwork_data_availableTask_ready;
	wire _stealServers_16_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_16_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_16_io_connQ_push_valid;
	wire [127:0] _stealServers_16_io_connQ_push_bits;
	wire _stealServers_16_io_connQ_pop_ready;
	wire _stealServers_15_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_15_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_15_io_connNetwork_data_availableTask_ready;
	wire _stealServers_15_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_15_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_15_io_connQ_push_valid;
	wire [127:0] _stealServers_15_io_connQ_push_bits;
	wire _stealServers_15_io_connQ_pop_ready;
	wire _stealServers_14_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_14_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_14_io_connNetwork_data_availableTask_ready;
	wire _stealServers_14_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_14_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_14_io_connQ_push_valid;
	wire [127:0] _stealServers_14_io_connQ_push_bits;
	wire _stealServers_14_io_connQ_pop_ready;
	wire _stealServers_13_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_13_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_13_io_connNetwork_data_availableTask_ready;
	wire _stealServers_13_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_13_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_13_io_connQ_push_valid;
	wire [127:0] _stealServers_13_io_connQ_push_bits;
	wire _stealServers_13_io_connQ_pop_ready;
	wire _stealServers_12_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_12_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_12_io_connNetwork_data_availableTask_ready;
	wire _stealServers_12_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_12_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_12_io_connQ_push_valid;
	wire [127:0] _stealServers_12_io_connQ_push_bits;
	wire _stealServers_12_io_connQ_pop_ready;
	wire _stealServers_11_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_11_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_11_io_connNetwork_data_availableTask_ready;
	wire _stealServers_11_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_11_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_11_io_connQ_push_valid;
	wire [127:0] _stealServers_11_io_connQ_push_bits;
	wire _stealServers_11_io_connQ_pop_ready;
	wire _stealServers_10_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_10_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_10_io_connNetwork_data_availableTask_ready;
	wire _stealServers_10_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_10_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_10_io_connQ_push_valid;
	wire [127:0] _stealServers_10_io_connQ_push_bits;
	wire _stealServers_10_io_connQ_pop_ready;
	wire _stealServers_9_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_9_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_9_io_connNetwork_data_availableTask_ready;
	wire _stealServers_9_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_9_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_9_io_connQ_push_valid;
	wire [127:0] _stealServers_9_io_connQ_push_bits;
	wire _stealServers_9_io_connQ_pop_ready;
	wire _stealServers_8_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_8_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_8_io_connNetwork_data_availableTask_ready;
	wire _stealServers_8_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_8_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_8_io_connQ_push_valid;
	wire [127:0] _stealServers_8_io_connQ_push_bits;
	wire _stealServers_8_io_connQ_pop_ready;
	wire _stealServers_7_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_7_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_7_io_connNetwork_data_availableTask_ready;
	wire _stealServers_7_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_7_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_7_io_connQ_push_valid;
	wire [127:0] _stealServers_7_io_connQ_push_bits;
	wire _stealServers_7_io_connQ_pop_ready;
	wire _stealServers_6_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_6_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_6_io_connNetwork_data_availableTask_ready;
	wire _stealServers_6_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_6_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_6_io_connQ_push_valid;
	wire [127:0] _stealServers_6_io_connQ_push_bits;
	wire _stealServers_6_io_connQ_pop_ready;
	wire _stealServers_5_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_5_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_5_io_connNetwork_data_availableTask_ready;
	wire _stealServers_5_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_5_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_5_io_connQ_push_valid;
	wire [127:0] _stealServers_5_io_connQ_push_bits;
	wire _stealServers_5_io_connQ_pop_ready;
	wire _stealServers_4_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_4_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_4_io_connNetwork_data_availableTask_ready;
	wire _stealServers_4_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_4_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_4_io_connQ_push_valid;
	wire [127:0] _stealServers_4_io_connQ_push_bits;
	wire _stealServers_4_io_connQ_pop_ready;
	wire _stealServers_3_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_3_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_3_io_connNetwork_data_availableTask_ready;
	wire _stealServers_3_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_3_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_3_io_connQ_push_valid;
	wire [127:0] _stealServers_3_io_connQ_push_bits;
	wire _stealServers_3_io_connQ_pop_ready;
	wire _stealServers_2_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_2_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_2_io_connNetwork_data_availableTask_ready;
	wire _stealServers_2_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_2_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_2_io_connQ_push_valid;
	wire [127:0] _stealServers_2_io_connQ_push_bits;
	wire _stealServers_2_io_connQ_pop_ready;
	wire _stealServers_1_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_1_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_1_io_connNetwork_data_availableTask_ready;
	wire _stealServers_1_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_1_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_1_io_connQ_push_valid;
	wire [127:0] _stealServers_1_io_connQ_push_bits;
	wire _stealServers_1_io_connQ_pop_ready;
	wire _stealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_0_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_0_io_connNetwork_data_availableTask_ready;
	wire _stealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_0_io_connQ_push_valid;
	wire [127:0] _stealServers_0_io_connQ_push_bits;
	wire _stealServers_0_io_connQ_pop_ready;
	wire _stealNet_io_connSS_1_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_1_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_1_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_1_data_availableTask_bits;
	wire _stealNet_io_connSS_1_data_qOutTask_ready;
	wire _stealNet_io_connSS_2_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_2_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_2_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_2_data_availableTask_bits;
	wire _stealNet_io_connSS_2_data_qOutTask_ready;
	wire _stealNet_io_connSS_3_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_3_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_3_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_3_data_availableTask_bits;
	wire _stealNet_io_connSS_3_data_qOutTask_ready;
	wire _stealNet_io_connSS_4_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_4_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_4_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_4_data_availableTask_bits;
	wire _stealNet_io_connSS_4_data_qOutTask_ready;
	wire _stealNet_io_connSS_5_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_5_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_5_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_5_data_availableTask_bits;
	wire _stealNet_io_connSS_5_data_qOutTask_ready;
	wire _stealNet_io_connSS_6_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_6_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_6_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_6_data_availableTask_bits;
	wire _stealNet_io_connSS_6_data_qOutTask_ready;
	wire _stealNet_io_connSS_7_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_7_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_7_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_7_data_availableTask_bits;
	wire _stealNet_io_connSS_7_data_qOutTask_ready;
	wire _stealNet_io_connSS_8_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_8_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_8_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_8_data_availableTask_bits;
	wire _stealNet_io_connSS_8_data_qOutTask_ready;
	wire _stealNet_io_connSS_9_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_9_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_9_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_9_data_availableTask_bits;
	wire _stealNet_io_connSS_9_data_qOutTask_ready;
	wire _stealNet_io_connSS_10_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_10_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_10_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_10_data_availableTask_bits;
	wire _stealNet_io_connSS_10_data_qOutTask_ready;
	wire _stealNet_io_connSS_11_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_11_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_11_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_11_data_availableTask_bits;
	wire _stealNet_io_connSS_11_data_qOutTask_ready;
	wire _stealNet_io_connSS_12_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_12_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_12_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_12_data_availableTask_bits;
	wire _stealNet_io_connSS_12_data_qOutTask_ready;
	wire _stealNet_io_connSS_13_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_13_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_13_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_13_data_availableTask_bits;
	wire _stealNet_io_connSS_13_data_qOutTask_ready;
	wire _stealNet_io_connSS_14_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_14_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_14_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_14_data_availableTask_bits;
	wire _stealNet_io_connSS_14_data_qOutTask_ready;
	wire _stealNet_io_connSS_15_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_15_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_15_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_15_data_availableTask_bits;
	wire _stealNet_io_connSS_15_data_qOutTask_ready;
	wire _stealNet_io_connSS_16_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_16_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_16_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_16_data_availableTask_bits;
	wire _stealNet_io_connSS_16_data_qOutTask_ready;
	wire _stealNet_io_connSS_17_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_17_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_17_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_17_data_availableTask_bits;
	wire _stealNet_io_connSS_17_data_qOutTask_ready;
	wire _stealNet_io_connSS_18_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_18_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_18_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_18_data_availableTask_bits;
	wire _stealNet_io_connSS_18_data_qOutTask_ready;
	wire _stealNet_io_connSS_19_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_19_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_19_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_19_data_availableTask_bits;
	wire _stealNet_io_connSS_19_data_qOutTask_ready;
	wire _stealNet_io_connSS_20_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_20_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_20_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_20_data_availableTask_bits;
	wire _stealNet_io_connSS_20_data_qOutTask_ready;
	wire _stealNet_io_connSS_21_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_21_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_21_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_21_data_availableTask_bits;
	wire _stealNet_io_connSS_21_data_qOutTask_ready;
	wire _stealNet_io_connSS_22_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_22_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_22_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_22_data_availableTask_bits;
	wire _stealNet_io_connSS_22_data_qOutTask_ready;
	wire _stealNet_io_connSS_23_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_23_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_23_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_23_data_availableTask_bits;
	wire _stealNet_io_connSS_23_data_qOutTask_ready;
	wire _stealNet_io_connSS_24_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_24_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_24_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_24_data_availableTask_bits;
	wire _stealNet_io_connSS_24_data_qOutTask_ready;
	wire _stealNet_io_connSS_25_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_25_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_25_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_25_data_availableTask_bits;
	wire _stealNet_io_connSS_25_data_qOutTask_ready;
	wire _stealNet_io_connSS_26_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_26_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_26_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_26_data_availableTask_bits;
	wire _stealNet_io_connSS_26_data_qOutTask_ready;
	wire _stealNet_io_connSS_27_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_27_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_27_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_27_data_availableTask_bits;
	wire _stealNet_io_connSS_27_data_qOutTask_ready;
	wire _stealNet_io_connSS_28_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_28_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_28_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_28_data_availableTask_bits;
	wire _stealNet_io_connSS_28_data_qOutTask_ready;
	wire _stealNet_io_connSS_29_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_29_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_29_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_29_data_availableTask_bits;
	wire _stealNet_io_connSS_29_data_qOutTask_ready;
	wire _stealNet_io_connSS_30_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_30_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_30_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_30_data_availableTask_bits;
	wire _stealNet_io_connSS_30_data_qOutTask_ready;
	wire _stealNet_io_connSS_31_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_31_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_31_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_31_data_availableTask_bits;
	wire _stealNet_io_connSS_31_data_qOutTask_ready;
	wire _stealNet_io_connSS_32_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_32_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_32_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_32_data_availableTask_bits;
	wire _stealNet_io_connSS_32_data_qOutTask_ready;
	wire _stealNet_io_connSS_34_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_34_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_34_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_34_data_availableTask_bits;
	wire _stealNet_io_connSS_34_data_qOutTask_ready;
	wire _stealNet_io_connSS_35_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_35_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_35_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_35_data_availableTask_bits;
	wire _stealNet_io_connSS_35_data_qOutTask_ready;
	wire _stealNet_io_connSS_36_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_36_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_36_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_36_data_availableTask_bits;
	wire _stealNet_io_connSS_36_data_qOutTask_ready;
	wire _stealNet_io_connSS_37_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_37_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_37_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_37_data_availableTask_bits;
	wire _stealNet_io_connSS_37_data_qOutTask_ready;
	wire _stealNet_io_connSS_38_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_38_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_38_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_38_data_availableTask_bits;
	wire _stealNet_io_connSS_38_data_qOutTask_ready;
	wire _stealNet_io_connSS_39_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_39_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_39_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_39_data_availableTask_bits;
	wire _stealNet_io_connSS_39_data_qOutTask_ready;
	wire _stealNet_io_connSS_40_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_40_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_40_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_40_data_availableTask_bits;
	wire _stealNet_io_connSS_40_data_qOutTask_ready;
	wire _stealNet_io_connSS_41_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_41_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_41_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_41_data_availableTask_bits;
	wire _stealNet_io_connSS_41_data_qOutTask_ready;
	wire _stealNet_io_connSS_42_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_42_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_42_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_42_data_availableTask_bits;
	wire _stealNet_io_connSS_42_data_qOutTask_ready;
	wire _stealNet_io_connSS_43_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_43_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_43_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_43_data_availableTask_bits;
	wire _stealNet_io_connSS_43_data_qOutTask_ready;
	wire _stealNet_io_connSS_44_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_44_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_44_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_44_data_availableTask_bits;
	wire _stealNet_io_connSS_44_data_qOutTask_ready;
	wire _stealNet_io_connSS_45_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_45_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_45_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_45_data_availableTask_bits;
	wire _stealNet_io_connSS_45_data_qOutTask_ready;
	wire _stealNet_io_connSS_46_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_46_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_46_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_46_data_availableTask_bits;
	wire _stealNet_io_connSS_46_data_qOutTask_ready;
	wire _stealNet_io_connSS_47_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_47_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_47_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_47_data_availableTask_bits;
	wire _stealNet_io_connSS_47_data_qOutTask_ready;
	wire _stealNet_io_connSS_48_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_48_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_48_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_48_data_availableTask_bits;
	wire _stealNet_io_connSS_48_data_qOutTask_ready;
	wire _stealNet_io_connSS_49_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_49_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_49_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_49_data_availableTask_bits;
	wire _stealNet_io_connSS_49_data_qOutTask_ready;
	wire _stealNet_io_connSS_50_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_50_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_50_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_50_data_availableTask_bits;
	wire _stealNet_io_connSS_50_data_qOutTask_ready;
	wire _stealNet_io_connSS_51_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_51_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_51_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_51_data_availableTask_bits;
	wire _stealNet_io_connSS_51_data_qOutTask_ready;
	wire _stealNet_io_connSS_52_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_52_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_52_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_52_data_availableTask_bits;
	wire _stealNet_io_connSS_52_data_qOutTask_ready;
	wire _stealNet_io_connSS_53_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_53_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_53_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_53_data_availableTask_bits;
	wire _stealNet_io_connSS_53_data_qOutTask_ready;
	wire _stealNet_io_connSS_54_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_54_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_54_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_54_data_availableTask_bits;
	wire _stealNet_io_connSS_54_data_qOutTask_ready;
	wire _stealNet_io_connSS_55_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_55_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_55_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_55_data_availableTask_bits;
	wire _stealNet_io_connSS_55_data_qOutTask_ready;
	wire _stealNet_io_connSS_56_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_56_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_56_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_56_data_availableTask_bits;
	wire _stealNet_io_connSS_56_data_qOutTask_ready;
	wire _stealNet_io_connSS_57_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_57_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_57_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_57_data_availableTask_bits;
	wire _stealNet_io_connSS_57_data_qOutTask_ready;
	wire _stealNet_io_connSS_58_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_58_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_58_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_58_data_availableTask_bits;
	wire _stealNet_io_connSS_58_data_qOutTask_ready;
	wire _stealNet_io_connSS_59_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_59_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_59_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_59_data_availableTask_bits;
	wire _stealNet_io_connSS_59_data_qOutTask_ready;
	wire _stealNet_io_connSS_60_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_60_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_60_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_60_data_availableTask_bits;
	wire _stealNet_io_connSS_60_data_qOutTask_ready;
	wire _stealNet_io_connSS_61_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_61_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_61_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_61_data_availableTask_bits;
	wire _stealNet_io_connSS_61_data_qOutTask_ready;
	wire _stealNet_io_connSS_62_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_62_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_62_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_62_data_availableTask_bits;
	wire _stealNet_io_connSS_62_data_qOutTask_ready;
	wire _stealNet_io_connSS_63_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_63_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_63_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_63_data_availableTask_bits;
	wire _stealNet_io_connSS_63_data_qOutTask_ready;
	wire _stealNet_io_connSS_64_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_64_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_64_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_64_data_availableTask_bits;
	wire _stealNet_io_connSS_64_data_qOutTask_ready;
	wire _stealNet_io_connSS_65_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_65_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_65_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_65_data_availableTask_bits;
	wire _stealNet_io_connSS_65_data_qOutTask_ready;
	SchedulerNetwork stealNet(
		.clock(clock),
		.reset(reset),
		.io_connSS_0_ctrl_serveStealReq_valid(io_connVSS_0_ctrl_serveStealReq_valid),
		.io_connSS_0_ctrl_serveStealReq_ready(io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connSS_0_data_availableTask_ready(io_connVSS_0_data_availableTask_ready),
		.io_connSS_0_data_availableTask_valid(io_connVSS_0_data_availableTask_valid),
		.io_connSS_0_data_availableTask_bits(io_connVSS_0_data_availableTask_bits),
		.io_connSS_0_data_qOutTask_ready(io_connVSS_0_data_qOutTask_ready),
		.io_connSS_0_data_qOutTask_valid(io_connVSS_0_data_qOutTask_valid),
		.io_connSS_0_data_qOutTask_bits(io_connVSS_0_data_qOutTask_bits),
		.io_connSS_1_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_1_ctrl_serveStealReq_ready(_stealNet_io_connSS_1_ctrl_serveStealReq_ready),
		.io_connSS_1_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_1_ctrl_stealReq_ready(_stealNet_io_connSS_1_ctrl_stealReq_ready),
		.io_connSS_1_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connSS_1_data_availableTask_valid(_stealNet_io_connSS_1_data_availableTask_valid),
		.io_connSS_1_data_availableTask_bits(_stealNet_io_connSS_1_data_availableTask_bits),
		.io_connSS_1_data_qOutTask_ready(_stealNet_io_connSS_1_data_qOutTask_ready),
		.io_connSS_1_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connSS_1_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connSS_2_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_2_ctrl_serveStealReq_ready(_stealNet_io_connSS_2_ctrl_serveStealReq_ready),
		.io_connSS_2_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_2_ctrl_stealReq_ready(_stealNet_io_connSS_2_ctrl_stealReq_ready),
		.io_connSS_2_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connSS_2_data_availableTask_valid(_stealNet_io_connSS_2_data_availableTask_valid),
		.io_connSS_2_data_availableTask_bits(_stealNet_io_connSS_2_data_availableTask_bits),
		.io_connSS_2_data_qOutTask_ready(_stealNet_io_connSS_2_data_qOutTask_ready),
		.io_connSS_2_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connSS_2_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connSS_3_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_3_ctrl_serveStealReq_ready(_stealNet_io_connSS_3_ctrl_serveStealReq_ready),
		.io_connSS_3_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_3_ctrl_stealReq_ready(_stealNet_io_connSS_3_ctrl_stealReq_ready),
		.io_connSS_3_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connSS_3_data_availableTask_valid(_stealNet_io_connSS_3_data_availableTask_valid),
		.io_connSS_3_data_availableTask_bits(_stealNet_io_connSS_3_data_availableTask_bits),
		.io_connSS_3_data_qOutTask_ready(_stealNet_io_connSS_3_data_qOutTask_ready),
		.io_connSS_3_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connSS_3_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connSS_4_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_4_ctrl_serveStealReq_ready(_stealNet_io_connSS_4_ctrl_serveStealReq_ready),
		.io_connSS_4_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_4_ctrl_stealReq_ready(_stealNet_io_connSS_4_ctrl_stealReq_ready),
		.io_connSS_4_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connSS_4_data_availableTask_valid(_stealNet_io_connSS_4_data_availableTask_valid),
		.io_connSS_4_data_availableTask_bits(_stealNet_io_connSS_4_data_availableTask_bits),
		.io_connSS_4_data_qOutTask_ready(_stealNet_io_connSS_4_data_qOutTask_ready),
		.io_connSS_4_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connSS_4_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connSS_5_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_5_ctrl_serveStealReq_ready(_stealNet_io_connSS_5_ctrl_serveStealReq_ready),
		.io_connSS_5_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_5_ctrl_stealReq_ready(_stealNet_io_connSS_5_ctrl_stealReq_ready),
		.io_connSS_5_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connSS_5_data_availableTask_valid(_stealNet_io_connSS_5_data_availableTask_valid),
		.io_connSS_5_data_availableTask_bits(_stealNet_io_connSS_5_data_availableTask_bits),
		.io_connSS_5_data_qOutTask_ready(_stealNet_io_connSS_5_data_qOutTask_ready),
		.io_connSS_5_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connSS_5_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connSS_6_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_6_ctrl_serveStealReq_ready(_stealNet_io_connSS_6_ctrl_serveStealReq_ready),
		.io_connSS_6_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_6_ctrl_stealReq_ready(_stealNet_io_connSS_6_ctrl_stealReq_ready),
		.io_connSS_6_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connSS_6_data_availableTask_valid(_stealNet_io_connSS_6_data_availableTask_valid),
		.io_connSS_6_data_availableTask_bits(_stealNet_io_connSS_6_data_availableTask_bits),
		.io_connSS_6_data_qOutTask_ready(_stealNet_io_connSS_6_data_qOutTask_ready),
		.io_connSS_6_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connSS_6_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connSS_7_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_7_ctrl_serveStealReq_ready(_stealNet_io_connSS_7_ctrl_serveStealReq_ready),
		.io_connSS_7_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_7_ctrl_stealReq_ready(_stealNet_io_connSS_7_ctrl_stealReq_ready),
		.io_connSS_7_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connSS_7_data_availableTask_valid(_stealNet_io_connSS_7_data_availableTask_valid),
		.io_connSS_7_data_availableTask_bits(_stealNet_io_connSS_7_data_availableTask_bits),
		.io_connSS_7_data_qOutTask_ready(_stealNet_io_connSS_7_data_qOutTask_ready),
		.io_connSS_7_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connSS_7_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connSS_8_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_8_ctrl_serveStealReq_ready(_stealNet_io_connSS_8_ctrl_serveStealReq_ready),
		.io_connSS_8_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_8_ctrl_stealReq_ready(_stealNet_io_connSS_8_ctrl_stealReq_ready),
		.io_connSS_8_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connSS_8_data_availableTask_valid(_stealNet_io_connSS_8_data_availableTask_valid),
		.io_connSS_8_data_availableTask_bits(_stealNet_io_connSS_8_data_availableTask_bits),
		.io_connSS_8_data_qOutTask_ready(_stealNet_io_connSS_8_data_qOutTask_ready),
		.io_connSS_8_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connSS_8_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connSS_9_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_9_ctrl_serveStealReq_ready(_stealNet_io_connSS_9_ctrl_serveStealReq_ready),
		.io_connSS_9_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_9_ctrl_stealReq_ready(_stealNet_io_connSS_9_ctrl_stealReq_ready),
		.io_connSS_9_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connSS_9_data_availableTask_valid(_stealNet_io_connSS_9_data_availableTask_valid),
		.io_connSS_9_data_availableTask_bits(_stealNet_io_connSS_9_data_availableTask_bits),
		.io_connSS_9_data_qOutTask_ready(_stealNet_io_connSS_9_data_qOutTask_ready),
		.io_connSS_9_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connSS_9_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connSS_10_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_10_ctrl_serveStealReq_ready(_stealNet_io_connSS_10_ctrl_serveStealReq_ready),
		.io_connSS_10_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_10_ctrl_stealReq_ready(_stealNet_io_connSS_10_ctrl_stealReq_ready),
		.io_connSS_10_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connSS_10_data_availableTask_valid(_stealNet_io_connSS_10_data_availableTask_valid),
		.io_connSS_10_data_availableTask_bits(_stealNet_io_connSS_10_data_availableTask_bits),
		.io_connSS_10_data_qOutTask_ready(_stealNet_io_connSS_10_data_qOutTask_ready),
		.io_connSS_10_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connSS_10_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connSS_11_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_11_ctrl_serveStealReq_ready(_stealNet_io_connSS_11_ctrl_serveStealReq_ready),
		.io_connSS_11_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_11_ctrl_stealReq_ready(_stealNet_io_connSS_11_ctrl_stealReq_ready),
		.io_connSS_11_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connSS_11_data_availableTask_valid(_stealNet_io_connSS_11_data_availableTask_valid),
		.io_connSS_11_data_availableTask_bits(_stealNet_io_connSS_11_data_availableTask_bits),
		.io_connSS_11_data_qOutTask_ready(_stealNet_io_connSS_11_data_qOutTask_ready),
		.io_connSS_11_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connSS_11_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connSS_12_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_12_ctrl_serveStealReq_ready(_stealNet_io_connSS_12_ctrl_serveStealReq_ready),
		.io_connSS_12_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_12_ctrl_stealReq_ready(_stealNet_io_connSS_12_ctrl_stealReq_ready),
		.io_connSS_12_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connSS_12_data_availableTask_valid(_stealNet_io_connSS_12_data_availableTask_valid),
		.io_connSS_12_data_availableTask_bits(_stealNet_io_connSS_12_data_availableTask_bits),
		.io_connSS_12_data_qOutTask_ready(_stealNet_io_connSS_12_data_qOutTask_ready),
		.io_connSS_12_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connSS_12_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connSS_13_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_13_ctrl_serveStealReq_ready(_stealNet_io_connSS_13_ctrl_serveStealReq_ready),
		.io_connSS_13_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_13_ctrl_stealReq_ready(_stealNet_io_connSS_13_ctrl_stealReq_ready),
		.io_connSS_13_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connSS_13_data_availableTask_valid(_stealNet_io_connSS_13_data_availableTask_valid),
		.io_connSS_13_data_availableTask_bits(_stealNet_io_connSS_13_data_availableTask_bits),
		.io_connSS_13_data_qOutTask_ready(_stealNet_io_connSS_13_data_qOutTask_ready),
		.io_connSS_13_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connSS_13_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connSS_14_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_14_ctrl_serveStealReq_ready(_stealNet_io_connSS_14_ctrl_serveStealReq_ready),
		.io_connSS_14_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_14_ctrl_stealReq_ready(_stealNet_io_connSS_14_ctrl_stealReq_ready),
		.io_connSS_14_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connSS_14_data_availableTask_valid(_stealNet_io_connSS_14_data_availableTask_valid),
		.io_connSS_14_data_availableTask_bits(_stealNet_io_connSS_14_data_availableTask_bits),
		.io_connSS_14_data_qOutTask_ready(_stealNet_io_connSS_14_data_qOutTask_ready),
		.io_connSS_14_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connSS_14_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connSS_15_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_15_ctrl_serveStealReq_ready(_stealNet_io_connSS_15_ctrl_serveStealReq_ready),
		.io_connSS_15_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_15_ctrl_stealReq_ready(_stealNet_io_connSS_15_ctrl_stealReq_ready),
		.io_connSS_15_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connSS_15_data_availableTask_valid(_stealNet_io_connSS_15_data_availableTask_valid),
		.io_connSS_15_data_availableTask_bits(_stealNet_io_connSS_15_data_availableTask_bits),
		.io_connSS_15_data_qOutTask_ready(_stealNet_io_connSS_15_data_qOutTask_ready),
		.io_connSS_15_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connSS_15_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connSS_16_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_16_ctrl_serveStealReq_ready(_stealNet_io_connSS_16_ctrl_serveStealReq_ready),
		.io_connSS_16_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_16_ctrl_stealReq_ready(_stealNet_io_connSS_16_ctrl_stealReq_ready),
		.io_connSS_16_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connSS_16_data_availableTask_valid(_stealNet_io_connSS_16_data_availableTask_valid),
		.io_connSS_16_data_availableTask_bits(_stealNet_io_connSS_16_data_availableTask_bits),
		.io_connSS_16_data_qOutTask_ready(_stealNet_io_connSS_16_data_qOutTask_ready),
		.io_connSS_16_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connSS_16_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connSS_17_ctrl_serveStealReq_valid(_stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_17_ctrl_serveStealReq_ready(_stealNet_io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_17_ctrl_stealReq_valid(_stealServers_16_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_17_ctrl_stealReq_ready(_stealNet_io_connSS_17_ctrl_stealReq_ready),
		.io_connSS_17_data_availableTask_ready(_stealServers_16_io_connNetwork_data_availableTask_ready),
		.io_connSS_17_data_availableTask_valid(_stealNet_io_connSS_17_data_availableTask_valid),
		.io_connSS_17_data_availableTask_bits(_stealNet_io_connSS_17_data_availableTask_bits),
		.io_connSS_17_data_qOutTask_ready(_stealNet_io_connSS_17_data_qOutTask_ready),
		.io_connSS_17_data_qOutTask_valid(_stealServers_16_io_connNetwork_data_qOutTask_valid),
		.io_connSS_17_data_qOutTask_bits(_stealServers_16_io_connNetwork_data_qOutTask_bits),
		.io_connSS_18_ctrl_serveStealReq_valid(_stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_18_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_18_ctrl_stealReq_valid(_stealServers_17_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_18_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connSS_18_data_availableTask_ready(_stealServers_17_io_connNetwork_data_availableTask_ready),
		.io_connSS_18_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connSS_18_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connSS_18_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connSS_18_data_qOutTask_valid(_stealServers_17_io_connNetwork_data_qOutTask_valid),
		.io_connSS_18_data_qOutTask_bits(_stealServers_17_io_connNetwork_data_qOutTask_bits),
		.io_connSS_19_ctrl_serveStealReq_valid(_stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_19_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_19_ctrl_stealReq_valid(_stealServers_18_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_19_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connSS_19_data_availableTask_ready(_stealServers_18_io_connNetwork_data_availableTask_ready),
		.io_connSS_19_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connSS_19_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connSS_19_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connSS_19_data_qOutTask_valid(_stealServers_18_io_connNetwork_data_qOutTask_valid),
		.io_connSS_19_data_qOutTask_bits(_stealServers_18_io_connNetwork_data_qOutTask_bits),
		.io_connSS_20_ctrl_serveStealReq_valid(_stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_20_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_20_ctrl_stealReq_valid(_stealServers_19_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_20_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connSS_20_data_availableTask_ready(_stealServers_19_io_connNetwork_data_availableTask_ready),
		.io_connSS_20_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connSS_20_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connSS_20_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connSS_20_data_qOutTask_valid(_stealServers_19_io_connNetwork_data_qOutTask_valid),
		.io_connSS_20_data_qOutTask_bits(_stealServers_19_io_connNetwork_data_qOutTask_bits),
		.io_connSS_21_ctrl_serveStealReq_valid(_stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_21_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_21_ctrl_stealReq_valid(_stealServers_20_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_21_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connSS_21_data_availableTask_ready(_stealServers_20_io_connNetwork_data_availableTask_ready),
		.io_connSS_21_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connSS_21_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connSS_21_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connSS_21_data_qOutTask_valid(_stealServers_20_io_connNetwork_data_qOutTask_valid),
		.io_connSS_21_data_qOutTask_bits(_stealServers_20_io_connNetwork_data_qOutTask_bits),
		.io_connSS_22_ctrl_serveStealReq_valid(_stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_22_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_22_ctrl_stealReq_valid(_stealServers_21_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_22_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connSS_22_data_availableTask_ready(_stealServers_21_io_connNetwork_data_availableTask_ready),
		.io_connSS_22_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connSS_22_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connSS_22_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connSS_22_data_qOutTask_valid(_stealServers_21_io_connNetwork_data_qOutTask_valid),
		.io_connSS_22_data_qOutTask_bits(_stealServers_21_io_connNetwork_data_qOutTask_bits),
		.io_connSS_23_ctrl_serveStealReq_valid(_stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_23_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_23_ctrl_stealReq_valid(_stealServers_22_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_23_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connSS_23_data_availableTask_ready(_stealServers_22_io_connNetwork_data_availableTask_ready),
		.io_connSS_23_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connSS_23_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connSS_23_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connSS_23_data_qOutTask_valid(_stealServers_22_io_connNetwork_data_qOutTask_valid),
		.io_connSS_23_data_qOutTask_bits(_stealServers_22_io_connNetwork_data_qOutTask_bits),
		.io_connSS_24_ctrl_serveStealReq_valid(_stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_24_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_24_ctrl_stealReq_valid(_stealServers_23_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_24_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connSS_24_data_availableTask_ready(_stealServers_23_io_connNetwork_data_availableTask_ready),
		.io_connSS_24_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connSS_24_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connSS_24_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connSS_24_data_qOutTask_valid(_stealServers_23_io_connNetwork_data_qOutTask_valid),
		.io_connSS_24_data_qOutTask_bits(_stealServers_23_io_connNetwork_data_qOutTask_bits),
		.io_connSS_25_ctrl_serveStealReq_valid(_stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_25_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_25_ctrl_stealReq_valid(_stealServers_24_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_25_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connSS_25_data_availableTask_ready(_stealServers_24_io_connNetwork_data_availableTask_ready),
		.io_connSS_25_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connSS_25_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connSS_25_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connSS_25_data_qOutTask_valid(_stealServers_24_io_connNetwork_data_qOutTask_valid),
		.io_connSS_25_data_qOutTask_bits(_stealServers_24_io_connNetwork_data_qOutTask_bits),
		.io_connSS_26_ctrl_serveStealReq_valid(_stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_26_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_26_ctrl_stealReq_valid(_stealServers_25_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_26_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connSS_26_data_availableTask_ready(_stealServers_25_io_connNetwork_data_availableTask_ready),
		.io_connSS_26_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connSS_26_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connSS_26_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connSS_26_data_qOutTask_valid(_stealServers_25_io_connNetwork_data_qOutTask_valid),
		.io_connSS_26_data_qOutTask_bits(_stealServers_25_io_connNetwork_data_qOutTask_bits),
		.io_connSS_27_ctrl_serveStealReq_valid(_stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_27_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_27_ctrl_stealReq_valid(_stealServers_26_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_27_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connSS_27_data_availableTask_ready(_stealServers_26_io_connNetwork_data_availableTask_ready),
		.io_connSS_27_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connSS_27_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connSS_27_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connSS_27_data_qOutTask_valid(_stealServers_26_io_connNetwork_data_qOutTask_valid),
		.io_connSS_27_data_qOutTask_bits(_stealServers_26_io_connNetwork_data_qOutTask_bits),
		.io_connSS_28_ctrl_serveStealReq_valid(_stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_28_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_28_ctrl_stealReq_valid(_stealServers_27_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_28_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connSS_28_data_availableTask_ready(_stealServers_27_io_connNetwork_data_availableTask_ready),
		.io_connSS_28_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connSS_28_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connSS_28_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connSS_28_data_qOutTask_valid(_stealServers_27_io_connNetwork_data_qOutTask_valid),
		.io_connSS_28_data_qOutTask_bits(_stealServers_27_io_connNetwork_data_qOutTask_bits),
		.io_connSS_29_ctrl_serveStealReq_valid(_stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_29_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_29_ctrl_stealReq_valid(_stealServers_28_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_29_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connSS_29_data_availableTask_ready(_stealServers_28_io_connNetwork_data_availableTask_ready),
		.io_connSS_29_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connSS_29_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connSS_29_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connSS_29_data_qOutTask_valid(_stealServers_28_io_connNetwork_data_qOutTask_valid),
		.io_connSS_29_data_qOutTask_bits(_stealServers_28_io_connNetwork_data_qOutTask_bits),
		.io_connSS_30_ctrl_serveStealReq_valid(_stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_30_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_30_ctrl_stealReq_valid(_stealServers_29_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_30_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connSS_30_data_availableTask_ready(_stealServers_29_io_connNetwork_data_availableTask_ready),
		.io_connSS_30_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connSS_30_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connSS_30_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connSS_30_data_qOutTask_valid(_stealServers_29_io_connNetwork_data_qOutTask_valid),
		.io_connSS_30_data_qOutTask_bits(_stealServers_29_io_connNetwork_data_qOutTask_bits),
		.io_connSS_31_ctrl_serveStealReq_valid(_stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_31_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_31_ctrl_stealReq_valid(_stealServers_30_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_31_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connSS_31_data_availableTask_ready(_stealServers_30_io_connNetwork_data_availableTask_ready),
		.io_connSS_31_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connSS_31_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connSS_31_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connSS_31_data_qOutTask_valid(_stealServers_30_io_connNetwork_data_qOutTask_valid),
		.io_connSS_31_data_qOutTask_bits(_stealServers_30_io_connNetwork_data_qOutTask_bits),
		.io_connSS_32_ctrl_serveStealReq_valid(_stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_32_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_32_ctrl_stealReq_valid(_stealServers_31_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_32_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connSS_32_data_availableTask_ready(_stealServers_31_io_connNetwork_data_availableTask_ready),
		.io_connSS_32_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connSS_32_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connSS_32_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connSS_32_data_qOutTask_valid(_stealServers_31_io_connNetwork_data_qOutTask_valid),
		.io_connSS_32_data_qOutTask_bits(_stealServers_31_io_connNetwork_data_qOutTask_bits),
		.io_connSS_33_ctrl_serveStealReq_valid(io_connVSS_1_ctrl_serveStealReq_valid),
		.io_connSS_33_ctrl_serveStealReq_ready(io_connVSS_1_ctrl_serveStealReq_ready),
		.io_connSS_33_data_availableTask_ready(io_connVSS_1_data_availableTask_ready),
		.io_connSS_33_data_availableTask_valid(io_connVSS_1_data_availableTask_valid),
		.io_connSS_33_data_availableTask_bits(io_connVSS_1_data_availableTask_bits),
		.io_connSS_33_data_qOutTask_ready(io_connVSS_1_data_qOutTask_ready),
		.io_connSS_33_data_qOutTask_valid(io_connVSS_1_data_qOutTask_valid),
		.io_connSS_33_data_qOutTask_bits(io_connVSS_1_data_qOutTask_bits),
		.io_connSS_34_ctrl_serveStealReq_valid(_stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_34_ctrl_serveStealReq_ready(_stealNet_io_connSS_34_ctrl_serveStealReq_ready),
		.io_connSS_34_ctrl_stealReq_valid(_stealServers_32_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_34_ctrl_stealReq_ready(_stealNet_io_connSS_34_ctrl_stealReq_ready),
		.io_connSS_34_data_availableTask_ready(_stealServers_32_io_connNetwork_data_availableTask_ready),
		.io_connSS_34_data_availableTask_valid(_stealNet_io_connSS_34_data_availableTask_valid),
		.io_connSS_34_data_availableTask_bits(_stealNet_io_connSS_34_data_availableTask_bits),
		.io_connSS_34_data_qOutTask_ready(_stealNet_io_connSS_34_data_qOutTask_ready),
		.io_connSS_34_data_qOutTask_valid(_stealServers_32_io_connNetwork_data_qOutTask_valid),
		.io_connSS_34_data_qOutTask_bits(_stealServers_32_io_connNetwork_data_qOutTask_bits),
		.io_connSS_35_ctrl_serveStealReq_valid(_stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_35_ctrl_serveStealReq_ready(_stealNet_io_connSS_35_ctrl_serveStealReq_ready),
		.io_connSS_35_ctrl_stealReq_valid(_stealServers_33_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_35_ctrl_stealReq_ready(_stealNet_io_connSS_35_ctrl_stealReq_ready),
		.io_connSS_35_data_availableTask_ready(_stealServers_33_io_connNetwork_data_availableTask_ready),
		.io_connSS_35_data_availableTask_valid(_stealNet_io_connSS_35_data_availableTask_valid),
		.io_connSS_35_data_availableTask_bits(_stealNet_io_connSS_35_data_availableTask_bits),
		.io_connSS_35_data_qOutTask_ready(_stealNet_io_connSS_35_data_qOutTask_ready),
		.io_connSS_35_data_qOutTask_valid(_stealServers_33_io_connNetwork_data_qOutTask_valid),
		.io_connSS_35_data_qOutTask_bits(_stealServers_33_io_connNetwork_data_qOutTask_bits),
		.io_connSS_36_ctrl_serveStealReq_valid(_stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_36_ctrl_serveStealReq_ready(_stealNet_io_connSS_36_ctrl_serveStealReq_ready),
		.io_connSS_36_ctrl_stealReq_valid(_stealServers_34_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_36_ctrl_stealReq_ready(_stealNet_io_connSS_36_ctrl_stealReq_ready),
		.io_connSS_36_data_availableTask_ready(_stealServers_34_io_connNetwork_data_availableTask_ready),
		.io_connSS_36_data_availableTask_valid(_stealNet_io_connSS_36_data_availableTask_valid),
		.io_connSS_36_data_availableTask_bits(_stealNet_io_connSS_36_data_availableTask_bits),
		.io_connSS_36_data_qOutTask_ready(_stealNet_io_connSS_36_data_qOutTask_ready),
		.io_connSS_36_data_qOutTask_valid(_stealServers_34_io_connNetwork_data_qOutTask_valid),
		.io_connSS_36_data_qOutTask_bits(_stealServers_34_io_connNetwork_data_qOutTask_bits),
		.io_connSS_37_ctrl_serveStealReq_valid(_stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_37_ctrl_serveStealReq_ready(_stealNet_io_connSS_37_ctrl_serveStealReq_ready),
		.io_connSS_37_ctrl_stealReq_valid(_stealServers_35_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_37_ctrl_stealReq_ready(_stealNet_io_connSS_37_ctrl_stealReq_ready),
		.io_connSS_37_data_availableTask_ready(_stealServers_35_io_connNetwork_data_availableTask_ready),
		.io_connSS_37_data_availableTask_valid(_stealNet_io_connSS_37_data_availableTask_valid),
		.io_connSS_37_data_availableTask_bits(_stealNet_io_connSS_37_data_availableTask_bits),
		.io_connSS_37_data_qOutTask_ready(_stealNet_io_connSS_37_data_qOutTask_ready),
		.io_connSS_37_data_qOutTask_valid(_stealServers_35_io_connNetwork_data_qOutTask_valid),
		.io_connSS_37_data_qOutTask_bits(_stealServers_35_io_connNetwork_data_qOutTask_bits),
		.io_connSS_38_ctrl_serveStealReq_valid(_stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_38_ctrl_serveStealReq_ready(_stealNet_io_connSS_38_ctrl_serveStealReq_ready),
		.io_connSS_38_ctrl_stealReq_valid(_stealServers_36_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_38_ctrl_stealReq_ready(_stealNet_io_connSS_38_ctrl_stealReq_ready),
		.io_connSS_38_data_availableTask_ready(_stealServers_36_io_connNetwork_data_availableTask_ready),
		.io_connSS_38_data_availableTask_valid(_stealNet_io_connSS_38_data_availableTask_valid),
		.io_connSS_38_data_availableTask_bits(_stealNet_io_connSS_38_data_availableTask_bits),
		.io_connSS_38_data_qOutTask_ready(_stealNet_io_connSS_38_data_qOutTask_ready),
		.io_connSS_38_data_qOutTask_valid(_stealServers_36_io_connNetwork_data_qOutTask_valid),
		.io_connSS_38_data_qOutTask_bits(_stealServers_36_io_connNetwork_data_qOutTask_bits),
		.io_connSS_39_ctrl_serveStealReq_valid(_stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_39_ctrl_serveStealReq_ready(_stealNet_io_connSS_39_ctrl_serveStealReq_ready),
		.io_connSS_39_ctrl_stealReq_valid(_stealServers_37_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_39_ctrl_stealReq_ready(_stealNet_io_connSS_39_ctrl_stealReq_ready),
		.io_connSS_39_data_availableTask_ready(_stealServers_37_io_connNetwork_data_availableTask_ready),
		.io_connSS_39_data_availableTask_valid(_stealNet_io_connSS_39_data_availableTask_valid),
		.io_connSS_39_data_availableTask_bits(_stealNet_io_connSS_39_data_availableTask_bits),
		.io_connSS_39_data_qOutTask_ready(_stealNet_io_connSS_39_data_qOutTask_ready),
		.io_connSS_39_data_qOutTask_valid(_stealServers_37_io_connNetwork_data_qOutTask_valid),
		.io_connSS_39_data_qOutTask_bits(_stealServers_37_io_connNetwork_data_qOutTask_bits),
		.io_connSS_40_ctrl_serveStealReq_valid(_stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_40_ctrl_serveStealReq_ready(_stealNet_io_connSS_40_ctrl_serveStealReq_ready),
		.io_connSS_40_ctrl_stealReq_valid(_stealServers_38_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_40_ctrl_stealReq_ready(_stealNet_io_connSS_40_ctrl_stealReq_ready),
		.io_connSS_40_data_availableTask_ready(_stealServers_38_io_connNetwork_data_availableTask_ready),
		.io_connSS_40_data_availableTask_valid(_stealNet_io_connSS_40_data_availableTask_valid),
		.io_connSS_40_data_availableTask_bits(_stealNet_io_connSS_40_data_availableTask_bits),
		.io_connSS_40_data_qOutTask_ready(_stealNet_io_connSS_40_data_qOutTask_ready),
		.io_connSS_40_data_qOutTask_valid(_stealServers_38_io_connNetwork_data_qOutTask_valid),
		.io_connSS_40_data_qOutTask_bits(_stealServers_38_io_connNetwork_data_qOutTask_bits),
		.io_connSS_41_ctrl_serveStealReq_valid(_stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_41_ctrl_serveStealReq_ready(_stealNet_io_connSS_41_ctrl_serveStealReq_ready),
		.io_connSS_41_ctrl_stealReq_valid(_stealServers_39_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_41_ctrl_stealReq_ready(_stealNet_io_connSS_41_ctrl_stealReq_ready),
		.io_connSS_41_data_availableTask_ready(_stealServers_39_io_connNetwork_data_availableTask_ready),
		.io_connSS_41_data_availableTask_valid(_stealNet_io_connSS_41_data_availableTask_valid),
		.io_connSS_41_data_availableTask_bits(_stealNet_io_connSS_41_data_availableTask_bits),
		.io_connSS_41_data_qOutTask_ready(_stealNet_io_connSS_41_data_qOutTask_ready),
		.io_connSS_41_data_qOutTask_valid(_stealServers_39_io_connNetwork_data_qOutTask_valid),
		.io_connSS_41_data_qOutTask_bits(_stealServers_39_io_connNetwork_data_qOutTask_bits),
		.io_connSS_42_ctrl_serveStealReq_valid(_stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_42_ctrl_serveStealReq_ready(_stealNet_io_connSS_42_ctrl_serveStealReq_ready),
		.io_connSS_42_ctrl_stealReq_valid(_stealServers_40_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_42_ctrl_stealReq_ready(_stealNet_io_connSS_42_ctrl_stealReq_ready),
		.io_connSS_42_data_availableTask_ready(_stealServers_40_io_connNetwork_data_availableTask_ready),
		.io_connSS_42_data_availableTask_valid(_stealNet_io_connSS_42_data_availableTask_valid),
		.io_connSS_42_data_availableTask_bits(_stealNet_io_connSS_42_data_availableTask_bits),
		.io_connSS_42_data_qOutTask_ready(_stealNet_io_connSS_42_data_qOutTask_ready),
		.io_connSS_42_data_qOutTask_valid(_stealServers_40_io_connNetwork_data_qOutTask_valid),
		.io_connSS_42_data_qOutTask_bits(_stealServers_40_io_connNetwork_data_qOutTask_bits),
		.io_connSS_43_ctrl_serveStealReq_valid(_stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_43_ctrl_serveStealReq_ready(_stealNet_io_connSS_43_ctrl_serveStealReq_ready),
		.io_connSS_43_ctrl_stealReq_valid(_stealServers_41_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_43_ctrl_stealReq_ready(_stealNet_io_connSS_43_ctrl_stealReq_ready),
		.io_connSS_43_data_availableTask_ready(_stealServers_41_io_connNetwork_data_availableTask_ready),
		.io_connSS_43_data_availableTask_valid(_stealNet_io_connSS_43_data_availableTask_valid),
		.io_connSS_43_data_availableTask_bits(_stealNet_io_connSS_43_data_availableTask_bits),
		.io_connSS_43_data_qOutTask_ready(_stealNet_io_connSS_43_data_qOutTask_ready),
		.io_connSS_43_data_qOutTask_valid(_stealServers_41_io_connNetwork_data_qOutTask_valid),
		.io_connSS_43_data_qOutTask_bits(_stealServers_41_io_connNetwork_data_qOutTask_bits),
		.io_connSS_44_ctrl_serveStealReq_valid(_stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_44_ctrl_serveStealReq_ready(_stealNet_io_connSS_44_ctrl_serveStealReq_ready),
		.io_connSS_44_ctrl_stealReq_valid(_stealServers_42_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_44_ctrl_stealReq_ready(_stealNet_io_connSS_44_ctrl_stealReq_ready),
		.io_connSS_44_data_availableTask_ready(_stealServers_42_io_connNetwork_data_availableTask_ready),
		.io_connSS_44_data_availableTask_valid(_stealNet_io_connSS_44_data_availableTask_valid),
		.io_connSS_44_data_availableTask_bits(_stealNet_io_connSS_44_data_availableTask_bits),
		.io_connSS_44_data_qOutTask_ready(_stealNet_io_connSS_44_data_qOutTask_ready),
		.io_connSS_44_data_qOutTask_valid(_stealServers_42_io_connNetwork_data_qOutTask_valid),
		.io_connSS_44_data_qOutTask_bits(_stealServers_42_io_connNetwork_data_qOutTask_bits),
		.io_connSS_45_ctrl_serveStealReq_valid(_stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_45_ctrl_serveStealReq_ready(_stealNet_io_connSS_45_ctrl_serveStealReq_ready),
		.io_connSS_45_ctrl_stealReq_valid(_stealServers_43_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_45_ctrl_stealReq_ready(_stealNet_io_connSS_45_ctrl_stealReq_ready),
		.io_connSS_45_data_availableTask_ready(_stealServers_43_io_connNetwork_data_availableTask_ready),
		.io_connSS_45_data_availableTask_valid(_stealNet_io_connSS_45_data_availableTask_valid),
		.io_connSS_45_data_availableTask_bits(_stealNet_io_connSS_45_data_availableTask_bits),
		.io_connSS_45_data_qOutTask_ready(_stealNet_io_connSS_45_data_qOutTask_ready),
		.io_connSS_45_data_qOutTask_valid(_stealServers_43_io_connNetwork_data_qOutTask_valid),
		.io_connSS_45_data_qOutTask_bits(_stealServers_43_io_connNetwork_data_qOutTask_bits),
		.io_connSS_46_ctrl_serveStealReq_valid(_stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_46_ctrl_serveStealReq_ready(_stealNet_io_connSS_46_ctrl_serveStealReq_ready),
		.io_connSS_46_ctrl_stealReq_valid(_stealServers_44_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_46_ctrl_stealReq_ready(_stealNet_io_connSS_46_ctrl_stealReq_ready),
		.io_connSS_46_data_availableTask_ready(_stealServers_44_io_connNetwork_data_availableTask_ready),
		.io_connSS_46_data_availableTask_valid(_stealNet_io_connSS_46_data_availableTask_valid),
		.io_connSS_46_data_availableTask_bits(_stealNet_io_connSS_46_data_availableTask_bits),
		.io_connSS_46_data_qOutTask_ready(_stealNet_io_connSS_46_data_qOutTask_ready),
		.io_connSS_46_data_qOutTask_valid(_stealServers_44_io_connNetwork_data_qOutTask_valid),
		.io_connSS_46_data_qOutTask_bits(_stealServers_44_io_connNetwork_data_qOutTask_bits),
		.io_connSS_47_ctrl_serveStealReq_valid(_stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_47_ctrl_serveStealReq_ready(_stealNet_io_connSS_47_ctrl_serveStealReq_ready),
		.io_connSS_47_ctrl_stealReq_valid(_stealServers_45_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_47_ctrl_stealReq_ready(_stealNet_io_connSS_47_ctrl_stealReq_ready),
		.io_connSS_47_data_availableTask_ready(_stealServers_45_io_connNetwork_data_availableTask_ready),
		.io_connSS_47_data_availableTask_valid(_stealNet_io_connSS_47_data_availableTask_valid),
		.io_connSS_47_data_availableTask_bits(_stealNet_io_connSS_47_data_availableTask_bits),
		.io_connSS_47_data_qOutTask_ready(_stealNet_io_connSS_47_data_qOutTask_ready),
		.io_connSS_47_data_qOutTask_valid(_stealServers_45_io_connNetwork_data_qOutTask_valid),
		.io_connSS_47_data_qOutTask_bits(_stealServers_45_io_connNetwork_data_qOutTask_bits),
		.io_connSS_48_ctrl_serveStealReq_valid(_stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_48_ctrl_serveStealReq_ready(_stealNet_io_connSS_48_ctrl_serveStealReq_ready),
		.io_connSS_48_ctrl_stealReq_valid(_stealServers_46_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_48_ctrl_stealReq_ready(_stealNet_io_connSS_48_ctrl_stealReq_ready),
		.io_connSS_48_data_availableTask_ready(_stealServers_46_io_connNetwork_data_availableTask_ready),
		.io_connSS_48_data_availableTask_valid(_stealNet_io_connSS_48_data_availableTask_valid),
		.io_connSS_48_data_availableTask_bits(_stealNet_io_connSS_48_data_availableTask_bits),
		.io_connSS_48_data_qOutTask_ready(_stealNet_io_connSS_48_data_qOutTask_ready),
		.io_connSS_48_data_qOutTask_valid(_stealServers_46_io_connNetwork_data_qOutTask_valid),
		.io_connSS_48_data_qOutTask_bits(_stealServers_46_io_connNetwork_data_qOutTask_bits),
		.io_connSS_49_ctrl_serveStealReq_valid(_stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_49_ctrl_serveStealReq_ready(_stealNet_io_connSS_49_ctrl_serveStealReq_ready),
		.io_connSS_49_ctrl_stealReq_valid(_stealServers_47_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_49_ctrl_stealReq_ready(_stealNet_io_connSS_49_ctrl_stealReq_ready),
		.io_connSS_49_data_availableTask_ready(_stealServers_47_io_connNetwork_data_availableTask_ready),
		.io_connSS_49_data_availableTask_valid(_stealNet_io_connSS_49_data_availableTask_valid),
		.io_connSS_49_data_availableTask_bits(_stealNet_io_connSS_49_data_availableTask_bits),
		.io_connSS_49_data_qOutTask_ready(_stealNet_io_connSS_49_data_qOutTask_ready),
		.io_connSS_49_data_qOutTask_valid(_stealServers_47_io_connNetwork_data_qOutTask_valid),
		.io_connSS_49_data_qOutTask_bits(_stealServers_47_io_connNetwork_data_qOutTask_bits),
		.io_connSS_50_ctrl_serveStealReq_valid(_stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_50_ctrl_serveStealReq_ready(_stealNet_io_connSS_50_ctrl_serveStealReq_ready),
		.io_connSS_50_ctrl_stealReq_valid(_stealServers_48_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_50_ctrl_stealReq_ready(_stealNet_io_connSS_50_ctrl_stealReq_ready),
		.io_connSS_50_data_availableTask_ready(_stealServers_48_io_connNetwork_data_availableTask_ready),
		.io_connSS_50_data_availableTask_valid(_stealNet_io_connSS_50_data_availableTask_valid),
		.io_connSS_50_data_availableTask_bits(_stealNet_io_connSS_50_data_availableTask_bits),
		.io_connSS_50_data_qOutTask_ready(_stealNet_io_connSS_50_data_qOutTask_ready),
		.io_connSS_50_data_qOutTask_valid(_stealServers_48_io_connNetwork_data_qOutTask_valid),
		.io_connSS_50_data_qOutTask_bits(_stealServers_48_io_connNetwork_data_qOutTask_bits),
		.io_connSS_51_ctrl_serveStealReq_valid(_stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_51_ctrl_serveStealReq_ready(_stealNet_io_connSS_51_ctrl_serveStealReq_ready),
		.io_connSS_51_ctrl_stealReq_valid(_stealServers_49_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_51_ctrl_stealReq_ready(_stealNet_io_connSS_51_ctrl_stealReq_ready),
		.io_connSS_51_data_availableTask_ready(_stealServers_49_io_connNetwork_data_availableTask_ready),
		.io_connSS_51_data_availableTask_valid(_stealNet_io_connSS_51_data_availableTask_valid),
		.io_connSS_51_data_availableTask_bits(_stealNet_io_connSS_51_data_availableTask_bits),
		.io_connSS_51_data_qOutTask_ready(_stealNet_io_connSS_51_data_qOutTask_ready),
		.io_connSS_51_data_qOutTask_valid(_stealServers_49_io_connNetwork_data_qOutTask_valid),
		.io_connSS_51_data_qOutTask_bits(_stealServers_49_io_connNetwork_data_qOutTask_bits),
		.io_connSS_52_ctrl_serveStealReq_valid(_stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_52_ctrl_serveStealReq_ready(_stealNet_io_connSS_52_ctrl_serveStealReq_ready),
		.io_connSS_52_ctrl_stealReq_valid(_stealServers_50_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_52_ctrl_stealReq_ready(_stealNet_io_connSS_52_ctrl_stealReq_ready),
		.io_connSS_52_data_availableTask_ready(_stealServers_50_io_connNetwork_data_availableTask_ready),
		.io_connSS_52_data_availableTask_valid(_stealNet_io_connSS_52_data_availableTask_valid),
		.io_connSS_52_data_availableTask_bits(_stealNet_io_connSS_52_data_availableTask_bits),
		.io_connSS_52_data_qOutTask_ready(_stealNet_io_connSS_52_data_qOutTask_ready),
		.io_connSS_52_data_qOutTask_valid(_stealServers_50_io_connNetwork_data_qOutTask_valid),
		.io_connSS_52_data_qOutTask_bits(_stealServers_50_io_connNetwork_data_qOutTask_bits),
		.io_connSS_53_ctrl_serveStealReq_valid(_stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_53_ctrl_serveStealReq_ready(_stealNet_io_connSS_53_ctrl_serveStealReq_ready),
		.io_connSS_53_ctrl_stealReq_valid(_stealServers_51_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_53_ctrl_stealReq_ready(_stealNet_io_connSS_53_ctrl_stealReq_ready),
		.io_connSS_53_data_availableTask_ready(_stealServers_51_io_connNetwork_data_availableTask_ready),
		.io_connSS_53_data_availableTask_valid(_stealNet_io_connSS_53_data_availableTask_valid),
		.io_connSS_53_data_availableTask_bits(_stealNet_io_connSS_53_data_availableTask_bits),
		.io_connSS_53_data_qOutTask_ready(_stealNet_io_connSS_53_data_qOutTask_ready),
		.io_connSS_53_data_qOutTask_valid(_stealServers_51_io_connNetwork_data_qOutTask_valid),
		.io_connSS_53_data_qOutTask_bits(_stealServers_51_io_connNetwork_data_qOutTask_bits),
		.io_connSS_54_ctrl_serveStealReq_valid(_stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_54_ctrl_serveStealReq_ready(_stealNet_io_connSS_54_ctrl_serveStealReq_ready),
		.io_connSS_54_ctrl_stealReq_valid(_stealServers_52_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_54_ctrl_stealReq_ready(_stealNet_io_connSS_54_ctrl_stealReq_ready),
		.io_connSS_54_data_availableTask_ready(_stealServers_52_io_connNetwork_data_availableTask_ready),
		.io_connSS_54_data_availableTask_valid(_stealNet_io_connSS_54_data_availableTask_valid),
		.io_connSS_54_data_availableTask_bits(_stealNet_io_connSS_54_data_availableTask_bits),
		.io_connSS_54_data_qOutTask_ready(_stealNet_io_connSS_54_data_qOutTask_ready),
		.io_connSS_54_data_qOutTask_valid(_stealServers_52_io_connNetwork_data_qOutTask_valid),
		.io_connSS_54_data_qOutTask_bits(_stealServers_52_io_connNetwork_data_qOutTask_bits),
		.io_connSS_55_ctrl_serveStealReq_valid(_stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_55_ctrl_serveStealReq_ready(_stealNet_io_connSS_55_ctrl_serveStealReq_ready),
		.io_connSS_55_ctrl_stealReq_valid(_stealServers_53_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_55_ctrl_stealReq_ready(_stealNet_io_connSS_55_ctrl_stealReq_ready),
		.io_connSS_55_data_availableTask_ready(_stealServers_53_io_connNetwork_data_availableTask_ready),
		.io_connSS_55_data_availableTask_valid(_stealNet_io_connSS_55_data_availableTask_valid),
		.io_connSS_55_data_availableTask_bits(_stealNet_io_connSS_55_data_availableTask_bits),
		.io_connSS_55_data_qOutTask_ready(_stealNet_io_connSS_55_data_qOutTask_ready),
		.io_connSS_55_data_qOutTask_valid(_stealServers_53_io_connNetwork_data_qOutTask_valid),
		.io_connSS_55_data_qOutTask_bits(_stealServers_53_io_connNetwork_data_qOutTask_bits),
		.io_connSS_56_ctrl_serveStealReq_valid(_stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_56_ctrl_serveStealReq_ready(_stealNet_io_connSS_56_ctrl_serveStealReq_ready),
		.io_connSS_56_ctrl_stealReq_valid(_stealServers_54_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_56_ctrl_stealReq_ready(_stealNet_io_connSS_56_ctrl_stealReq_ready),
		.io_connSS_56_data_availableTask_ready(_stealServers_54_io_connNetwork_data_availableTask_ready),
		.io_connSS_56_data_availableTask_valid(_stealNet_io_connSS_56_data_availableTask_valid),
		.io_connSS_56_data_availableTask_bits(_stealNet_io_connSS_56_data_availableTask_bits),
		.io_connSS_56_data_qOutTask_ready(_stealNet_io_connSS_56_data_qOutTask_ready),
		.io_connSS_56_data_qOutTask_valid(_stealServers_54_io_connNetwork_data_qOutTask_valid),
		.io_connSS_56_data_qOutTask_bits(_stealServers_54_io_connNetwork_data_qOutTask_bits),
		.io_connSS_57_ctrl_serveStealReq_valid(_stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_57_ctrl_serveStealReq_ready(_stealNet_io_connSS_57_ctrl_serveStealReq_ready),
		.io_connSS_57_ctrl_stealReq_valid(_stealServers_55_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_57_ctrl_stealReq_ready(_stealNet_io_connSS_57_ctrl_stealReq_ready),
		.io_connSS_57_data_availableTask_ready(_stealServers_55_io_connNetwork_data_availableTask_ready),
		.io_connSS_57_data_availableTask_valid(_stealNet_io_connSS_57_data_availableTask_valid),
		.io_connSS_57_data_availableTask_bits(_stealNet_io_connSS_57_data_availableTask_bits),
		.io_connSS_57_data_qOutTask_ready(_stealNet_io_connSS_57_data_qOutTask_ready),
		.io_connSS_57_data_qOutTask_valid(_stealServers_55_io_connNetwork_data_qOutTask_valid),
		.io_connSS_57_data_qOutTask_bits(_stealServers_55_io_connNetwork_data_qOutTask_bits),
		.io_connSS_58_ctrl_serveStealReq_valid(_stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_58_ctrl_serveStealReq_ready(_stealNet_io_connSS_58_ctrl_serveStealReq_ready),
		.io_connSS_58_ctrl_stealReq_valid(_stealServers_56_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_58_ctrl_stealReq_ready(_stealNet_io_connSS_58_ctrl_stealReq_ready),
		.io_connSS_58_data_availableTask_ready(_stealServers_56_io_connNetwork_data_availableTask_ready),
		.io_connSS_58_data_availableTask_valid(_stealNet_io_connSS_58_data_availableTask_valid),
		.io_connSS_58_data_availableTask_bits(_stealNet_io_connSS_58_data_availableTask_bits),
		.io_connSS_58_data_qOutTask_ready(_stealNet_io_connSS_58_data_qOutTask_ready),
		.io_connSS_58_data_qOutTask_valid(_stealServers_56_io_connNetwork_data_qOutTask_valid),
		.io_connSS_58_data_qOutTask_bits(_stealServers_56_io_connNetwork_data_qOutTask_bits),
		.io_connSS_59_ctrl_serveStealReq_valid(_stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_59_ctrl_serveStealReq_ready(_stealNet_io_connSS_59_ctrl_serveStealReq_ready),
		.io_connSS_59_ctrl_stealReq_valid(_stealServers_57_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_59_ctrl_stealReq_ready(_stealNet_io_connSS_59_ctrl_stealReq_ready),
		.io_connSS_59_data_availableTask_ready(_stealServers_57_io_connNetwork_data_availableTask_ready),
		.io_connSS_59_data_availableTask_valid(_stealNet_io_connSS_59_data_availableTask_valid),
		.io_connSS_59_data_availableTask_bits(_stealNet_io_connSS_59_data_availableTask_bits),
		.io_connSS_59_data_qOutTask_ready(_stealNet_io_connSS_59_data_qOutTask_ready),
		.io_connSS_59_data_qOutTask_valid(_stealServers_57_io_connNetwork_data_qOutTask_valid),
		.io_connSS_59_data_qOutTask_bits(_stealServers_57_io_connNetwork_data_qOutTask_bits),
		.io_connSS_60_ctrl_serveStealReq_valid(_stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_60_ctrl_serveStealReq_ready(_stealNet_io_connSS_60_ctrl_serveStealReq_ready),
		.io_connSS_60_ctrl_stealReq_valid(_stealServers_58_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_60_ctrl_stealReq_ready(_stealNet_io_connSS_60_ctrl_stealReq_ready),
		.io_connSS_60_data_availableTask_ready(_stealServers_58_io_connNetwork_data_availableTask_ready),
		.io_connSS_60_data_availableTask_valid(_stealNet_io_connSS_60_data_availableTask_valid),
		.io_connSS_60_data_availableTask_bits(_stealNet_io_connSS_60_data_availableTask_bits),
		.io_connSS_60_data_qOutTask_ready(_stealNet_io_connSS_60_data_qOutTask_ready),
		.io_connSS_60_data_qOutTask_valid(_stealServers_58_io_connNetwork_data_qOutTask_valid),
		.io_connSS_60_data_qOutTask_bits(_stealServers_58_io_connNetwork_data_qOutTask_bits),
		.io_connSS_61_ctrl_serveStealReq_valid(_stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_61_ctrl_serveStealReq_ready(_stealNet_io_connSS_61_ctrl_serveStealReq_ready),
		.io_connSS_61_ctrl_stealReq_valid(_stealServers_59_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_61_ctrl_stealReq_ready(_stealNet_io_connSS_61_ctrl_stealReq_ready),
		.io_connSS_61_data_availableTask_ready(_stealServers_59_io_connNetwork_data_availableTask_ready),
		.io_connSS_61_data_availableTask_valid(_stealNet_io_connSS_61_data_availableTask_valid),
		.io_connSS_61_data_availableTask_bits(_stealNet_io_connSS_61_data_availableTask_bits),
		.io_connSS_61_data_qOutTask_ready(_stealNet_io_connSS_61_data_qOutTask_ready),
		.io_connSS_61_data_qOutTask_valid(_stealServers_59_io_connNetwork_data_qOutTask_valid),
		.io_connSS_61_data_qOutTask_bits(_stealServers_59_io_connNetwork_data_qOutTask_bits),
		.io_connSS_62_ctrl_serveStealReq_valid(_stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_62_ctrl_serveStealReq_ready(_stealNet_io_connSS_62_ctrl_serveStealReq_ready),
		.io_connSS_62_ctrl_stealReq_valid(_stealServers_60_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_62_ctrl_stealReq_ready(_stealNet_io_connSS_62_ctrl_stealReq_ready),
		.io_connSS_62_data_availableTask_ready(_stealServers_60_io_connNetwork_data_availableTask_ready),
		.io_connSS_62_data_availableTask_valid(_stealNet_io_connSS_62_data_availableTask_valid),
		.io_connSS_62_data_availableTask_bits(_stealNet_io_connSS_62_data_availableTask_bits),
		.io_connSS_62_data_qOutTask_ready(_stealNet_io_connSS_62_data_qOutTask_ready),
		.io_connSS_62_data_qOutTask_valid(_stealServers_60_io_connNetwork_data_qOutTask_valid),
		.io_connSS_62_data_qOutTask_bits(_stealServers_60_io_connNetwork_data_qOutTask_bits),
		.io_connSS_63_ctrl_serveStealReq_valid(_stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_63_ctrl_serveStealReq_ready(_stealNet_io_connSS_63_ctrl_serveStealReq_ready),
		.io_connSS_63_ctrl_stealReq_valid(_stealServers_61_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_63_ctrl_stealReq_ready(_stealNet_io_connSS_63_ctrl_stealReq_ready),
		.io_connSS_63_data_availableTask_ready(_stealServers_61_io_connNetwork_data_availableTask_ready),
		.io_connSS_63_data_availableTask_valid(_stealNet_io_connSS_63_data_availableTask_valid),
		.io_connSS_63_data_availableTask_bits(_stealNet_io_connSS_63_data_availableTask_bits),
		.io_connSS_63_data_qOutTask_ready(_stealNet_io_connSS_63_data_qOutTask_ready),
		.io_connSS_63_data_qOutTask_valid(_stealServers_61_io_connNetwork_data_qOutTask_valid),
		.io_connSS_63_data_qOutTask_bits(_stealServers_61_io_connNetwork_data_qOutTask_bits),
		.io_connSS_64_ctrl_serveStealReq_valid(_stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_64_ctrl_serveStealReq_ready(_stealNet_io_connSS_64_ctrl_serveStealReq_ready),
		.io_connSS_64_ctrl_stealReq_valid(_stealServers_62_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_64_ctrl_stealReq_ready(_stealNet_io_connSS_64_ctrl_stealReq_ready),
		.io_connSS_64_data_availableTask_ready(_stealServers_62_io_connNetwork_data_availableTask_ready),
		.io_connSS_64_data_availableTask_valid(_stealNet_io_connSS_64_data_availableTask_valid),
		.io_connSS_64_data_availableTask_bits(_stealNet_io_connSS_64_data_availableTask_bits),
		.io_connSS_64_data_qOutTask_ready(_stealNet_io_connSS_64_data_qOutTask_ready),
		.io_connSS_64_data_qOutTask_valid(_stealServers_62_io_connNetwork_data_qOutTask_valid),
		.io_connSS_64_data_qOutTask_bits(_stealServers_62_io_connNetwork_data_qOutTask_bits),
		.io_connSS_65_ctrl_serveStealReq_valid(_stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_65_ctrl_serveStealReq_ready(_stealNet_io_connSS_65_ctrl_serveStealReq_ready),
		.io_connSS_65_ctrl_stealReq_valid(_stealServers_63_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_65_ctrl_stealReq_ready(_stealNet_io_connSS_65_ctrl_stealReq_ready),
		.io_connSS_65_data_availableTask_ready(_stealServers_63_io_connNetwork_data_availableTask_ready),
		.io_connSS_65_data_availableTask_valid(_stealNet_io_connSS_65_data_availableTask_valid),
		.io_connSS_65_data_availableTask_bits(_stealNet_io_connSS_65_data_availableTask_bits),
		.io_connSS_65_data_qOutTask_ready(_stealNet_io_connSS_65_data_qOutTask_ready),
		.io_connSS_65_data_qOutTask_valid(_stealServers_63_io_connNetwork_data_qOutTask_valid),
		.io_connSS_65_data_qOutTask_bits(_stealServers_63_io_connNetwork_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(io_ntwDataUnitOccupancyVSS_0),
		.io_ntwDataUnitOccupancyVSS_1(io_ntwDataUnitOccupancyVSS_1)
	);
	SchedulerClient stealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_1_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_1_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_1_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_1_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_1_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_0_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_2_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_2_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_2_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_2_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_2_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_1_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_2(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_3_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_3_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_3_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_3_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_3_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_2_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_3(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_4_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_4_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_4_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_4_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_4_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_3_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_4(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_5_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_5_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_5_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_5_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_5_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_4_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_5(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_6_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_6_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_6_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_6_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_6_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_5_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_6(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_7_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_7_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_7_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_7_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_7_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_6_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_7(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_8_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_8_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_8_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_8_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_8_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_7_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_8(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_9_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_9_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_9_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_9_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_9_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_8_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_9(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_10_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_10_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_10_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_10_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_10_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_9_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_10(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_11_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_11_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_11_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_11_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_11_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_10_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_11(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_12_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_12_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_12_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_12_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_12_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_11_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_12(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_13_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_13_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_13_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_13_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_13_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_12_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_13(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_14_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_14_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_14_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_14_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_14_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_13_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_14(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_15_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_15_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_15_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_15_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_15_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_14_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_15(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_16_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_16_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_16_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_16_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_16_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_15_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_16(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_17_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_16_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_17_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_16_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_17_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_17_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_17_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_16_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_16_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_16_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_16_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_16_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_16_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_16_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_16_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_16_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_17(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_17_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_17_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_17_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_17_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_17_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_17_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_17_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_17_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_17_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_17_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_17_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_18(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_18_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_18_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_18_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_18_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_18_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_18_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_18_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_18_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_18_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_18_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_18_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_19(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_19_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_19_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_19_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_19_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_19_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_19_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_19_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_19_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_19_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_19_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_19_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_20(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_20_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_20_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_20_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_20_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_20_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_20_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_20_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_20_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_20_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_20_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_20_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_21(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_21_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_21_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_21_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_21_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_21_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_21_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_21_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_21_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_21_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_21_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_21_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_22(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_22_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_22_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_22_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_22_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_22_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_22_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_22_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_22_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_22_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_22_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_22_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_23(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_23_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_23_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_23_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_23_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_23_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_23_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_23_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_23_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_23_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_23_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_23_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_24(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_24_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_24_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_24_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_24_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_24_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_24_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_24_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_24_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_24_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_24_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_24_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_25(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_25_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_25_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_25_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_25_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_25_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_25_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_25_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_25_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_25_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_25_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_25_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_26(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_26_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_26_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_26_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_26_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_26_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_26_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_26_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_26_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_26_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_26_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_26_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_27(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_27_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_27_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_27_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_27_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_27_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_27_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_27_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_27_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_27_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_27_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_27_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_28(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_28_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_28_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_28_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_28_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_28_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_28_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_28_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_28_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_28_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_28_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_28_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_29(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_29_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_29_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_29_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_29_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_29_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_29_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_29_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_29_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_29_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_29_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_29_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_30(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_30_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_30_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_30_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_30_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_30_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_30_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_30_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_30_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_30_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_30_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_30_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_31(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_31_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_31_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_31_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_31_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_31_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_31_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_31_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_31_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_31_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_31_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_31_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_32(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_34_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_32_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_34_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_32_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_34_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_34_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_34_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_32_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_32_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_32_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_32_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_32_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_32_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_32_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_32_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_32_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_33(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_35_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_33_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_35_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_33_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_35_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_35_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_35_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_33_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_33_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_33_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_33_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_33_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_33_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_33_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_33_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_33_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_34(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_36_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_34_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_36_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_34_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_36_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_36_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_36_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_34_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_34_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_34_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_34_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_34_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_34_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_34_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_34_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_34_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_35(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_37_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_35_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_37_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_35_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_37_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_37_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_37_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_35_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_35_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_35_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_35_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_35_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_35_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_35_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_35_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_35_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_36(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_38_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_36_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_38_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_36_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_38_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_38_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_38_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_36_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_36_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_36_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_36_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_36_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_36_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_36_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_36_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_36_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_37(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_39_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_37_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_39_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_37_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_39_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_39_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_39_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_37_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_37_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_37_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_37_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_37_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_37_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_37_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_37_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_37_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_38(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_40_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_38_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_40_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_38_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_40_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_40_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_40_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_38_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_38_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_38_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_38_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_38_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_38_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_38_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_38_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_38_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_39(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_41_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_39_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_41_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_39_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_41_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_41_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_41_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_39_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_39_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_39_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_39_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_39_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_39_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_39_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_39_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_39_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_40(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_42_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_40_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_42_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_40_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_42_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_42_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_42_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_40_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_40_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_40_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_40_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_40_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_40_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_40_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_40_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_40_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_41(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_43_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_41_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_43_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_41_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_43_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_43_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_43_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_41_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_41_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_41_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_41_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_41_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_41_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_41_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_41_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_41_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_42(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_44_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_42_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_44_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_42_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_44_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_44_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_44_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_42_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_42_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_42_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_42_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_42_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_42_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_42_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_42_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_42_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_43(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_45_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_43_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_45_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_43_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_45_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_45_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_45_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_43_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_43_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_43_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_43_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_43_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_43_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_43_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_43_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_43_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_44(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_46_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_44_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_46_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_44_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_46_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_46_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_46_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_44_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_44_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_44_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_44_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_44_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_44_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_44_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_44_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_44_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_45(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_47_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_45_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_47_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_45_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_47_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_47_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_47_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_45_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_45_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_45_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_45_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_45_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_45_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_45_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_45_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_45_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_46(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_48_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_46_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_48_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_46_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_48_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_48_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_48_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_46_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_46_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_46_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_46_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_46_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_46_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_46_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_46_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_46_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_47(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_49_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_47_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_49_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_47_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_49_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_49_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_49_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_47_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_47_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_47_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_47_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_47_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_47_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_47_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_47_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_47_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_48(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_50_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_48_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_50_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_48_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_50_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_50_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_50_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_48_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_48_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_48_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_48_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_48_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_48_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_48_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_48_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_48_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_49(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_51_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_49_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_51_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_49_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_51_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_51_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_51_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_49_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_49_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_49_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_49_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_49_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_49_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_49_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_49_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_49_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_50(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_52_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_50_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_52_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_50_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_52_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_52_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_52_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_50_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_50_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_50_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_50_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_50_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_50_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_50_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_50_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_50_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_51(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_53_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_51_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_53_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_51_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_53_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_53_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_53_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_51_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_51_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_51_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_51_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_51_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_51_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_51_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_51_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_51_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_52(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_54_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_52_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_54_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_52_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_54_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_54_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_54_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_52_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_52_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_52_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_52_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_52_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_52_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_52_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_52_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_52_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_53(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_55_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_53_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_55_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_53_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_55_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_55_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_55_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_53_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_53_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_53_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_53_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_53_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_53_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_53_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_53_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_53_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_54(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_56_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_54_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_56_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_54_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_56_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_56_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_56_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_54_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_54_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_54_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_54_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_54_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_54_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_54_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_54_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_54_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_55(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_57_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_55_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_57_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_55_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_57_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_57_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_57_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_55_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_55_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_55_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_55_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_55_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_55_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_55_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_55_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_55_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_56(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_58_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_56_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_58_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_56_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_58_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_58_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_58_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_56_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_56_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_56_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_56_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_56_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_56_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_56_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_56_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_56_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_57(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_59_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_57_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_59_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_57_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_59_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_59_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_59_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_57_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_57_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_57_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_57_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_57_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_57_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_57_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_57_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_57_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_58(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_60_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_58_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_60_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_58_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_60_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_60_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_60_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_58_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_58_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_58_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_58_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_58_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_58_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_58_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_58_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_58_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_59(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_61_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_59_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_61_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_59_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_61_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_61_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_61_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_59_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_59_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_59_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_59_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_59_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_59_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_59_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_59_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_59_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_60(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_62_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_60_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_62_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_60_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_62_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_62_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_62_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_60_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_60_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_60_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_60_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_60_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_60_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_60_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_60_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_60_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_61(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_63_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_61_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_63_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_61_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_63_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_63_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_63_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_61_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_61_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_61_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_61_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_61_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_61_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_61_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_61_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_61_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_62(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_64_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_62_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_64_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_62_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_64_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_64_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_64_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_62_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_62_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_62_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_62_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_62_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_62_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_62_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_62_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_62_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_63(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_65_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_63_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_65_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_63_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_65_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_65_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_65_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_63_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_63_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_63_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_63_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_63_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_63_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_63_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_63_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_63_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_0(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_0_push_ready),
		.io_connVec_0_push_valid(io_connPE_0_push_valid),
		.io_connVec_0_push_bits(io_connPE_0_push_bits),
		.io_connVec_0_pop_ready(io_connPE_0_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_0_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_0_pop_bits),
		.io_connVec_1_currLength(_taskQueues_0_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_1(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_1_push_ready),
		.io_connVec_0_push_valid(io_connPE_1_push_valid),
		.io_connVec_0_push_bits(io_connPE_1_push_bits),
		.io_connVec_0_pop_ready(io_connPE_1_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_1_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_1_pop_bits),
		.io_connVec_1_currLength(_taskQueues_1_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_2(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_2_push_ready),
		.io_connVec_0_push_valid(io_connPE_2_push_valid),
		.io_connVec_0_push_bits(io_connPE_2_push_bits),
		.io_connVec_0_pop_ready(io_connPE_2_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_2_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_2_pop_bits),
		.io_connVec_1_currLength(_taskQueues_2_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_3(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_3_push_ready),
		.io_connVec_0_push_valid(io_connPE_3_push_valid),
		.io_connVec_0_push_bits(io_connPE_3_push_bits),
		.io_connVec_0_pop_ready(io_connPE_3_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_3_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_3_pop_bits),
		.io_connVec_1_currLength(_taskQueues_3_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_4(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_4_push_ready),
		.io_connVec_0_push_valid(io_connPE_4_push_valid),
		.io_connVec_0_push_bits(io_connPE_4_push_bits),
		.io_connVec_0_pop_ready(io_connPE_4_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_4_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_4_pop_bits),
		.io_connVec_1_currLength(_taskQueues_4_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_5(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_5_push_ready),
		.io_connVec_0_push_valid(io_connPE_5_push_valid),
		.io_connVec_0_push_bits(io_connPE_5_push_bits),
		.io_connVec_0_pop_ready(io_connPE_5_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_5_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_5_pop_bits),
		.io_connVec_1_currLength(_taskQueues_5_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_6(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_6_push_ready),
		.io_connVec_0_push_valid(io_connPE_6_push_valid),
		.io_connVec_0_push_bits(io_connPE_6_push_bits),
		.io_connVec_0_pop_ready(io_connPE_6_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_6_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_6_pop_bits),
		.io_connVec_1_currLength(_taskQueues_6_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_7(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_7_push_ready),
		.io_connVec_0_push_valid(io_connPE_7_push_valid),
		.io_connVec_0_push_bits(io_connPE_7_push_bits),
		.io_connVec_0_pop_ready(io_connPE_7_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_7_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_7_pop_bits),
		.io_connVec_1_currLength(_taskQueues_7_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_8(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_8_push_ready),
		.io_connVec_0_push_valid(io_connPE_8_push_valid),
		.io_connVec_0_push_bits(io_connPE_8_push_bits),
		.io_connVec_0_pop_ready(io_connPE_8_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_8_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_8_pop_bits),
		.io_connVec_1_currLength(_taskQueues_8_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_9(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_9_push_ready),
		.io_connVec_0_push_valid(io_connPE_9_push_valid),
		.io_connVec_0_push_bits(io_connPE_9_push_bits),
		.io_connVec_0_pop_ready(io_connPE_9_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_9_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_9_pop_bits),
		.io_connVec_1_currLength(_taskQueues_9_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_10(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_10_push_ready),
		.io_connVec_0_push_valid(io_connPE_10_push_valid),
		.io_connVec_0_push_bits(io_connPE_10_push_bits),
		.io_connVec_0_pop_ready(io_connPE_10_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_10_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_10_pop_bits),
		.io_connVec_1_currLength(_taskQueues_10_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_11(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_11_push_ready),
		.io_connVec_0_push_valid(io_connPE_11_push_valid),
		.io_connVec_0_push_bits(io_connPE_11_push_bits),
		.io_connVec_0_pop_ready(io_connPE_11_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_11_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_11_pop_bits),
		.io_connVec_1_currLength(_taskQueues_11_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_12(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_12_push_ready),
		.io_connVec_0_push_valid(io_connPE_12_push_valid),
		.io_connVec_0_push_bits(io_connPE_12_push_bits),
		.io_connVec_0_pop_ready(io_connPE_12_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_12_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_12_pop_bits),
		.io_connVec_1_currLength(_taskQueues_12_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_13(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_13_push_ready),
		.io_connVec_0_push_valid(io_connPE_13_push_valid),
		.io_connVec_0_push_bits(io_connPE_13_push_bits),
		.io_connVec_0_pop_ready(io_connPE_13_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_13_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_13_pop_bits),
		.io_connVec_1_currLength(_taskQueues_13_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_14(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_14_push_ready),
		.io_connVec_0_push_valid(io_connPE_14_push_valid),
		.io_connVec_0_push_bits(io_connPE_14_push_bits),
		.io_connVec_0_pop_ready(io_connPE_14_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_14_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_14_pop_bits),
		.io_connVec_1_currLength(_taskQueues_14_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_15(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_15_push_ready),
		.io_connVec_0_push_valid(io_connPE_15_push_valid),
		.io_connVec_0_push_bits(io_connPE_15_push_bits),
		.io_connVec_0_pop_ready(io_connPE_15_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_15_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_15_pop_bits),
		.io_connVec_1_currLength(_taskQueues_15_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_16(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_16_push_ready),
		.io_connVec_0_push_valid(io_connPE_16_push_valid),
		.io_connVec_0_push_bits(io_connPE_16_push_bits),
		.io_connVec_0_pop_ready(io_connPE_16_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_16_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_16_pop_bits),
		.io_connVec_1_currLength(_taskQueues_16_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_16_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_16_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_16_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_16_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_16_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_16_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_17(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_17_push_ready),
		.io_connVec_0_push_valid(io_connPE_17_push_valid),
		.io_connVec_0_push_bits(io_connPE_17_push_bits),
		.io_connVec_0_pop_ready(io_connPE_17_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_17_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_17_pop_bits),
		.io_connVec_1_currLength(_taskQueues_17_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_17_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_17_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_17_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_17_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_17_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_17_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_18(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_18_push_ready),
		.io_connVec_0_push_valid(io_connPE_18_push_valid),
		.io_connVec_0_push_bits(io_connPE_18_push_bits),
		.io_connVec_0_pop_ready(io_connPE_18_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_18_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_18_pop_bits),
		.io_connVec_1_currLength(_taskQueues_18_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_18_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_18_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_18_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_18_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_18_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_18_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_19(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_19_push_ready),
		.io_connVec_0_push_valid(io_connPE_19_push_valid),
		.io_connVec_0_push_bits(io_connPE_19_push_bits),
		.io_connVec_0_pop_ready(io_connPE_19_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_19_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_19_pop_bits),
		.io_connVec_1_currLength(_taskQueues_19_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_19_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_19_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_19_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_19_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_19_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_19_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_20(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_20_push_ready),
		.io_connVec_0_push_valid(io_connPE_20_push_valid),
		.io_connVec_0_push_bits(io_connPE_20_push_bits),
		.io_connVec_0_pop_ready(io_connPE_20_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_20_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_20_pop_bits),
		.io_connVec_1_currLength(_taskQueues_20_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_20_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_20_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_20_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_20_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_20_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_20_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_21(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_21_push_ready),
		.io_connVec_0_push_valid(io_connPE_21_push_valid),
		.io_connVec_0_push_bits(io_connPE_21_push_bits),
		.io_connVec_0_pop_ready(io_connPE_21_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_21_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_21_pop_bits),
		.io_connVec_1_currLength(_taskQueues_21_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_21_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_21_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_21_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_21_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_21_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_21_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_22(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_22_push_ready),
		.io_connVec_0_push_valid(io_connPE_22_push_valid),
		.io_connVec_0_push_bits(io_connPE_22_push_bits),
		.io_connVec_0_pop_ready(io_connPE_22_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_22_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_22_pop_bits),
		.io_connVec_1_currLength(_taskQueues_22_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_22_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_22_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_22_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_22_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_22_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_22_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_23(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_23_push_ready),
		.io_connVec_0_push_valid(io_connPE_23_push_valid),
		.io_connVec_0_push_bits(io_connPE_23_push_bits),
		.io_connVec_0_pop_ready(io_connPE_23_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_23_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_23_pop_bits),
		.io_connVec_1_currLength(_taskQueues_23_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_23_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_23_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_23_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_23_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_23_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_23_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_24(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_24_push_ready),
		.io_connVec_0_push_valid(io_connPE_24_push_valid),
		.io_connVec_0_push_bits(io_connPE_24_push_bits),
		.io_connVec_0_pop_ready(io_connPE_24_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_24_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_24_pop_bits),
		.io_connVec_1_currLength(_taskQueues_24_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_24_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_24_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_24_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_24_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_24_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_24_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_25(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_25_push_ready),
		.io_connVec_0_push_valid(io_connPE_25_push_valid),
		.io_connVec_0_push_bits(io_connPE_25_push_bits),
		.io_connVec_0_pop_ready(io_connPE_25_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_25_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_25_pop_bits),
		.io_connVec_1_currLength(_taskQueues_25_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_25_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_25_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_25_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_25_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_25_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_25_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_26(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_26_push_ready),
		.io_connVec_0_push_valid(io_connPE_26_push_valid),
		.io_connVec_0_push_bits(io_connPE_26_push_bits),
		.io_connVec_0_pop_ready(io_connPE_26_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_26_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_26_pop_bits),
		.io_connVec_1_currLength(_taskQueues_26_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_26_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_26_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_26_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_26_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_26_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_26_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_27(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_27_push_ready),
		.io_connVec_0_push_valid(io_connPE_27_push_valid),
		.io_connVec_0_push_bits(io_connPE_27_push_bits),
		.io_connVec_0_pop_ready(io_connPE_27_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_27_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_27_pop_bits),
		.io_connVec_1_currLength(_taskQueues_27_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_27_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_27_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_27_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_27_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_27_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_27_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_28(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_28_push_ready),
		.io_connVec_0_push_valid(io_connPE_28_push_valid),
		.io_connVec_0_push_bits(io_connPE_28_push_bits),
		.io_connVec_0_pop_ready(io_connPE_28_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_28_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_28_pop_bits),
		.io_connVec_1_currLength(_taskQueues_28_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_28_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_28_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_28_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_28_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_28_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_28_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_29(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_29_push_ready),
		.io_connVec_0_push_valid(io_connPE_29_push_valid),
		.io_connVec_0_push_bits(io_connPE_29_push_bits),
		.io_connVec_0_pop_ready(io_connPE_29_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_29_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_29_pop_bits),
		.io_connVec_1_currLength(_taskQueues_29_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_29_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_29_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_29_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_29_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_29_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_29_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_30(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_30_push_ready),
		.io_connVec_0_push_valid(io_connPE_30_push_valid),
		.io_connVec_0_push_bits(io_connPE_30_push_bits),
		.io_connVec_0_pop_ready(io_connPE_30_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_30_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_30_pop_bits),
		.io_connVec_1_currLength(_taskQueues_30_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_30_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_30_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_30_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_30_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_30_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_30_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_31(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_31_push_ready),
		.io_connVec_0_push_valid(io_connPE_31_push_valid),
		.io_connVec_0_push_bits(io_connPE_31_push_bits),
		.io_connVec_0_pop_ready(io_connPE_31_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_31_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_31_pop_bits),
		.io_connVec_1_currLength(_taskQueues_31_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_31_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_31_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_31_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_31_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_31_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_31_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_32(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_32_push_ready),
		.io_connVec_0_push_valid(io_connPE_32_push_valid),
		.io_connVec_0_push_bits(io_connPE_32_push_bits),
		.io_connVec_0_pop_ready(io_connPE_32_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_32_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_32_pop_bits),
		.io_connVec_1_currLength(_taskQueues_32_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_32_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_32_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_32_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_32_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_32_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_32_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_33(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_33_push_ready),
		.io_connVec_0_push_valid(io_connPE_33_push_valid),
		.io_connVec_0_push_bits(io_connPE_33_push_bits),
		.io_connVec_0_pop_ready(io_connPE_33_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_33_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_33_pop_bits),
		.io_connVec_1_currLength(_taskQueues_33_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_33_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_33_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_33_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_33_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_33_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_33_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_34(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_34_push_ready),
		.io_connVec_0_push_valid(io_connPE_34_push_valid),
		.io_connVec_0_push_bits(io_connPE_34_push_bits),
		.io_connVec_0_pop_ready(io_connPE_34_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_34_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_34_pop_bits),
		.io_connVec_1_currLength(_taskQueues_34_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_34_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_34_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_34_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_34_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_34_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_34_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_35(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_35_push_ready),
		.io_connVec_0_push_valid(io_connPE_35_push_valid),
		.io_connVec_0_push_bits(io_connPE_35_push_bits),
		.io_connVec_0_pop_ready(io_connPE_35_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_35_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_35_pop_bits),
		.io_connVec_1_currLength(_taskQueues_35_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_35_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_35_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_35_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_35_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_35_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_35_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_36(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_36_push_ready),
		.io_connVec_0_push_valid(io_connPE_36_push_valid),
		.io_connVec_0_push_bits(io_connPE_36_push_bits),
		.io_connVec_0_pop_ready(io_connPE_36_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_36_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_36_pop_bits),
		.io_connVec_1_currLength(_taskQueues_36_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_36_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_36_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_36_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_36_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_36_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_36_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_37(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_37_push_ready),
		.io_connVec_0_push_valid(io_connPE_37_push_valid),
		.io_connVec_0_push_bits(io_connPE_37_push_bits),
		.io_connVec_0_pop_ready(io_connPE_37_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_37_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_37_pop_bits),
		.io_connVec_1_currLength(_taskQueues_37_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_37_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_37_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_37_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_37_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_37_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_37_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_38(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_38_push_ready),
		.io_connVec_0_push_valid(io_connPE_38_push_valid),
		.io_connVec_0_push_bits(io_connPE_38_push_bits),
		.io_connVec_0_pop_ready(io_connPE_38_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_38_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_38_pop_bits),
		.io_connVec_1_currLength(_taskQueues_38_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_38_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_38_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_38_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_38_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_38_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_38_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_39(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_39_push_ready),
		.io_connVec_0_push_valid(io_connPE_39_push_valid),
		.io_connVec_0_push_bits(io_connPE_39_push_bits),
		.io_connVec_0_pop_ready(io_connPE_39_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_39_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_39_pop_bits),
		.io_connVec_1_currLength(_taskQueues_39_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_39_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_39_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_39_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_39_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_39_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_39_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_40(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_40_push_ready),
		.io_connVec_0_push_valid(io_connPE_40_push_valid),
		.io_connVec_0_push_bits(io_connPE_40_push_bits),
		.io_connVec_0_pop_ready(io_connPE_40_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_40_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_40_pop_bits),
		.io_connVec_1_currLength(_taskQueues_40_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_40_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_40_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_40_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_40_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_40_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_40_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_41(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_41_push_ready),
		.io_connVec_0_push_valid(io_connPE_41_push_valid),
		.io_connVec_0_push_bits(io_connPE_41_push_bits),
		.io_connVec_0_pop_ready(io_connPE_41_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_41_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_41_pop_bits),
		.io_connVec_1_currLength(_taskQueues_41_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_41_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_41_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_41_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_41_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_41_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_41_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_42(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_42_push_ready),
		.io_connVec_0_push_valid(io_connPE_42_push_valid),
		.io_connVec_0_push_bits(io_connPE_42_push_bits),
		.io_connVec_0_pop_ready(io_connPE_42_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_42_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_42_pop_bits),
		.io_connVec_1_currLength(_taskQueues_42_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_42_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_42_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_42_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_42_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_42_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_42_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_43(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_43_push_ready),
		.io_connVec_0_push_valid(io_connPE_43_push_valid),
		.io_connVec_0_push_bits(io_connPE_43_push_bits),
		.io_connVec_0_pop_ready(io_connPE_43_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_43_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_43_pop_bits),
		.io_connVec_1_currLength(_taskQueues_43_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_43_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_43_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_43_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_43_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_43_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_43_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_44(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_44_push_ready),
		.io_connVec_0_push_valid(io_connPE_44_push_valid),
		.io_connVec_0_push_bits(io_connPE_44_push_bits),
		.io_connVec_0_pop_ready(io_connPE_44_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_44_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_44_pop_bits),
		.io_connVec_1_currLength(_taskQueues_44_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_44_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_44_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_44_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_44_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_44_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_44_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_45(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_45_push_ready),
		.io_connVec_0_push_valid(io_connPE_45_push_valid),
		.io_connVec_0_push_bits(io_connPE_45_push_bits),
		.io_connVec_0_pop_ready(io_connPE_45_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_45_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_45_pop_bits),
		.io_connVec_1_currLength(_taskQueues_45_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_45_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_45_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_45_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_45_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_45_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_45_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_46(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_46_push_ready),
		.io_connVec_0_push_valid(io_connPE_46_push_valid),
		.io_connVec_0_push_bits(io_connPE_46_push_bits),
		.io_connVec_0_pop_ready(io_connPE_46_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_46_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_46_pop_bits),
		.io_connVec_1_currLength(_taskQueues_46_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_46_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_46_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_46_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_46_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_46_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_46_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_47(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_47_push_ready),
		.io_connVec_0_push_valid(io_connPE_47_push_valid),
		.io_connVec_0_push_bits(io_connPE_47_push_bits),
		.io_connVec_0_pop_ready(io_connPE_47_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_47_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_47_pop_bits),
		.io_connVec_1_currLength(_taskQueues_47_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_47_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_47_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_47_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_47_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_47_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_47_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_48(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_48_push_ready),
		.io_connVec_0_push_valid(io_connPE_48_push_valid),
		.io_connVec_0_push_bits(io_connPE_48_push_bits),
		.io_connVec_0_pop_ready(io_connPE_48_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_48_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_48_pop_bits),
		.io_connVec_1_currLength(_taskQueues_48_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_48_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_48_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_48_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_48_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_48_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_48_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_49(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_49_push_ready),
		.io_connVec_0_push_valid(io_connPE_49_push_valid),
		.io_connVec_0_push_bits(io_connPE_49_push_bits),
		.io_connVec_0_pop_ready(io_connPE_49_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_49_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_49_pop_bits),
		.io_connVec_1_currLength(_taskQueues_49_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_49_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_49_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_49_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_49_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_49_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_49_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_50(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_50_push_ready),
		.io_connVec_0_push_valid(io_connPE_50_push_valid),
		.io_connVec_0_push_bits(io_connPE_50_push_bits),
		.io_connVec_0_pop_ready(io_connPE_50_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_50_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_50_pop_bits),
		.io_connVec_1_currLength(_taskQueues_50_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_50_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_50_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_50_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_50_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_50_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_50_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_51(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_51_push_ready),
		.io_connVec_0_push_valid(io_connPE_51_push_valid),
		.io_connVec_0_push_bits(io_connPE_51_push_bits),
		.io_connVec_0_pop_ready(io_connPE_51_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_51_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_51_pop_bits),
		.io_connVec_1_currLength(_taskQueues_51_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_51_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_51_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_51_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_51_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_51_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_51_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_52(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_52_push_ready),
		.io_connVec_0_push_valid(io_connPE_52_push_valid),
		.io_connVec_0_push_bits(io_connPE_52_push_bits),
		.io_connVec_0_pop_ready(io_connPE_52_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_52_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_52_pop_bits),
		.io_connVec_1_currLength(_taskQueues_52_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_52_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_52_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_52_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_52_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_52_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_52_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_53(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_53_push_ready),
		.io_connVec_0_push_valid(io_connPE_53_push_valid),
		.io_connVec_0_push_bits(io_connPE_53_push_bits),
		.io_connVec_0_pop_ready(io_connPE_53_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_53_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_53_pop_bits),
		.io_connVec_1_currLength(_taskQueues_53_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_53_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_53_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_53_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_53_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_53_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_53_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_54(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_54_push_ready),
		.io_connVec_0_push_valid(io_connPE_54_push_valid),
		.io_connVec_0_push_bits(io_connPE_54_push_bits),
		.io_connVec_0_pop_ready(io_connPE_54_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_54_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_54_pop_bits),
		.io_connVec_1_currLength(_taskQueues_54_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_54_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_54_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_54_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_54_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_54_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_54_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_55(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_55_push_ready),
		.io_connVec_0_push_valid(io_connPE_55_push_valid),
		.io_connVec_0_push_bits(io_connPE_55_push_bits),
		.io_connVec_0_pop_ready(io_connPE_55_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_55_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_55_pop_bits),
		.io_connVec_1_currLength(_taskQueues_55_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_55_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_55_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_55_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_55_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_55_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_55_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_56(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_56_push_ready),
		.io_connVec_0_push_valid(io_connPE_56_push_valid),
		.io_connVec_0_push_bits(io_connPE_56_push_bits),
		.io_connVec_0_pop_ready(io_connPE_56_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_56_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_56_pop_bits),
		.io_connVec_1_currLength(_taskQueues_56_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_56_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_56_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_56_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_56_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_56_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_56_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_57(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_57_push_ready),
		.io_connVec_0_push_valid(io_connPE_57_push_valid),
		.io_connVec_0_push_bits(io_connPE_57_push_bits),
		.io_connVec_0_pop_ready(io_connPE_57_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_57_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_57_pop_bits),
		.io_connVec_1_currLength(_taskQueues_57_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_57_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_57_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_57_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_57_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_57_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_57_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_58(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_58_push_ready),
		.io_connVec_0_push_valid(io_connPE_58_push_valid),
		.io_connVec_0_push_bits(io_connPE_58_push_bits),
		.io_connVec_0_pop_ready(io_connPE_58_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_58_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_58_pop_bits),
		.io_connVec_1_currLength(_taskQueues_58_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_58_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_58_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_58_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_58_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_58_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_58_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_59(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_59_push_ready),
		.io_connVec_0_push_valid(io_connPE_59_push_valid),
		.io_connVec_0_push_bits(io_connPE_59_push_bits),
		.io_connVec_0_pop_ready(io_connPE_59_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_59_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_59_pop_bits),
		.io_connVec_1_currLength(_taskQueues_59_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_59_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_59_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_59_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_59_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_59_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_59_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_60(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_60_push_ready),
		.io_connVec_0_push_valid(io_connPE_60_push_valid),
		.io_connVec_0_push_bits(io_connPE_60_push_bits),
		.io_connVec_0_pop_ready(io_connPE_60_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_60_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_60_pop_bits),
		.io_connVec_1_currLength(_taskQueues_60_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_60_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_60_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_60_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_60_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_60_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_60_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_61(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_61_push_ready),
		.io_connVec_0_push_valid(io_connPE_61_push_valid),
		.io_connVec_0_push_bits(io_connPE_61_push_bits),
		.io_connVec_0_pop_ready(io_connPE_61_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_61_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_61_pop_bits),
		.io_connVec_1_currLength(_taskQueues_61_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_61_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_61_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_61_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_61_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_61_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_61_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_62(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_62_push_ready),
		.io_connVec_0_push_valid(io_connPE_62_push_valid),
		.io_connVec_0_push_bits(io_connPE_62_push_bits),
		.io_connVec_0_pop_ready(io_connPE_62_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_62_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_62_pop_bits),
		.io_connVec_1_currLength(_taskQueues_62_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_62_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_62_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_62_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_62_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_62_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_62_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_63(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_63_push_ready),
		.io_connVec_0_push_valid(io_connPE_63_push_valid),
		.io_connVec_0_push_bits(io_connPE_63_push_bits),
		.io_connVec_0_pop_ready(io_connPE_63_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_63_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_63_pop_bits),
		.io_connVec_1_currLength(_taskQueues_63_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_63_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_63_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_63_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_63_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_63_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_63_io_connVec_1_pop_bits)
	);
endmodule
module ram_2x9 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [8:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [8:0] W0_data;
	reg [8:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 9'bxxxxxxxxx);
endmodule
module Queue2_AddressChannel_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_prot,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_prot
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [5:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_prot;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [5:0] io_deq_bits_addr;
	output wire [2:0] io_deq_bits_prot;
	wire [8:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x9 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_prot, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[5:0];
	assign io_deq_bits_prot = _ram_ext_R0_data[8:6];
endmodule
module Queue1_AddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_prot,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [5:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_prot;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [5:0] io_deq_bits_addr;
	reg [8:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_prot, io_enq_bits_addr};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_addr = ram[5:0];
endmodule
module Queue1_ReadDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	reg [65:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {2'h0, io_enq_bits_data};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[63:0];
	assign io_deq_bits_resp = ram[65:64];
endmodule
module Queue1_WriteDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [7:0] io_enq_bits_strb;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [7:0] io_deq_bits_strb;
	reg [71:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_strb, io_enq_bits_data};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[63:0];
	assign io_deq_bits_strb = ram[71:64];
endmodule
module Queue1_WriteResponseChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_deq_ready,
	io_deq_valid
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_deq_ready;
	output wire io_deq_valid;
	reg full;
	always @(posedge clock)
		if (reset)
			full <= 1'h0;
		else begin : sv2v_autoblock_1
			reg do_enq;
			do_enq = ~full & io_enq_valid;
			if (~(do_enq == (io_deq_ready & full)))
				full <= do_enq;
		end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
endmodule
module ram_16x128 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [3:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [127:0] R0_data;
	input [3:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [127:0] W0_data;
	reg [127:0] Memory [0:15];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue16_UInt (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_bits,
	io_count
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [127:0] io_enq_bits;
	input io_deq_ready;
	output wire [127:0] io_deq_bits;
	output wire [4:0] io_count;
	reg [3:0] enq_ptr_value;
	reg [3:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 4'h0;
			deq_ptr_value <= 4'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~(ptr_match & ~maybe_full);
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 4'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 4'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_16x128 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_count = {maybe_full & ptr_match, enq_ptr_value - deq_ptr_value};
endmodule
module SchedulerServer (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_axi_mgmt_ar_ready,
	io_axi_mgmt_ar_valid,
	io_axi_mgmt_ar_bits_addr,
	io_axi_mgmt_ar_bits_prot,
	io_axi_mgmt_r_ready,
	io_axi_mgmt_r_valid,
	io_axi_mgmt_r_bits_data,
	io_axi_mgmt_r_bits_resp,
	io_axi_mgmt_aw_ready,
	io_axi_mgmt_aw_valid,
	io_axi_mgmt_aw_bits_addr,
	io_axi_mgmt_aw_bits_prot,
	io_axi_mgmt_w_ready,
	io_axi_mgmt_w_valid,
	io_axi_mgmt_w_bits_data,
	io_axi_mgmt_w_bits_strb,
	io_axi_mgmt_b_ready,
	io_axi_mgmt_b_valid,
	io_axi_mgmt_b_bits_resp,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_read_burst_len,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_write_burst_len,
	io_write_last,
	io_ntwDataUnitOccupancy
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [127:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [127:0] io_connNetwork_data_qOutTask_bits;
	output wire io_axi_mgmt_ar_ready;
	input io_axi_mgmt_ar_valid;
	input [5:0] io_axi_mgmt_ar_bits_addr;
	input [2:0] io_axi_mgmt_ar_bits_prot;
	input io_axi_mgmt_r_ready;
	output wire io_axi_mgmt_r_valid;
	output wire [63:0] io_axi_mgmt_r_bits_data;
	output wire [1:0] io_axi_mgmt_r_bits_resp;
	output wire io_axi_mgmt_aw_ready;
	input io_axi_mgmt_aw_valid;
	input [5:0] io_axi_mgmt_aw_bits_addr;
	input [2:0] io_axi_mgmt_aw_bits_prot;
	output wire io_axi_mgmt_w_ready;
	input io_axi_mgmt_w_valid;
	input [63:0] io_axi_mgmt_w_bits_data;
	input [7:0] io_axi_mgmt_w_bits_strb;
	input io_axi_mgmt_b_ready;
	output wire io_axi_mgmt_b_valid;
	output wire [1:0] io_axi_mgmt_b_bits_resp;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [127:0] io_read_data_bits;
	output wire [3:0] io_read_burst_len;
	input io_write_address_ready;
	output wire io_write_address_valid;
	output wire [63:0] io_write_address_bits;
	input io_write_data_ready;
	output wire io_write_data_valid;
	output wire [127:0] io_write_data_bits;
	output wire [3:0] io_write_burst_len;
	output wire io_write_last;
	input io_ntwDataUnitOccupancy;
	wire _taskQueueBuffer_io_enq_ready;
	wire [127:0] _taskQueueBuffer_io_deq_bits;
	wire [4:0] _taskQueueBuffer_io_count;
	wire _wrRespQueue__io_enq_ready;
	wire _wrRespQueue__io_deq_valid;
	wire _wrReqData__deq_q_io_enq_ready;
	wire _wrReqData__deq_q_io_deq_valid;
	wire [63:0] _wrReqData__deq_q_io_deq_bits_data;
	wire [7:0] _wrReqData__deq_q_io_deq_bits_strb;
	wire _wrReq__deq_q_io_enq_ready;
	wire _wrReq__deq_q_io_deq_valid;
	wire [5:0] _wrReq__deq_q_io_deq_bits_addr;
	wire _rdRespQueue__io_enq_ready;
	wire _rdRespQueue__io_deq_valid;
	wire [63:0] _rdRespQueue__io_deq_bits_data;
	wire [1:0] _rdRespQueue__io_deq_bits_resp;
	wire _rdReq__deq_q_io_enq_ready;
	wire _rdReq__deq_q_io_deq_valid;
	wire [5:0] _rdReq__deq_q_io_deq_bits_addr;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	wire rdReq = _rdReq__deq_q_io_deq_valid & _rdRespQueue__io_enq_ready;
	wire wrReq = (_wrReq__deq_q_io_deq_valid & _wrReqData__deq_q_io_deq_valid) & _wrRespQueue__io_enq_ready;
	reg [63:0] rAddr;
	reg [63:0] rPause;
	reg [63:0] procInterrupt;
	reg [63:0] maxLength;
	reg [3:0] stateReg;
	reg [63:0] currLen;
	reg [63:0] contentionCounter;
	reg networkCongested;
	reg [63:0] fifoTailReg;
	reg [63:0] fifoHeadReg;
	reg [4:0] memDataCounter;
	wire _GEN = stateReg == 4'h2;
	wire _GEN_0 = stateReg == 4'h4;
	wire _GEN_1 = stateReg == 4'h3;
	wire _GEN_2 = memDataCounter == 5'h01;
	wire _GEN_3 = _GEN | _GEN_0;
	wire _GEN_4 = stateReg == 4'h6;
	wire _GEN_5 = stateReg == 4'h5;
	wire _GEN_6 = (_GEN_0 | _GEN_1) | _GEN_4;
	wire _GEN_7 = _GEN | _GEN_6;
	wire _GEN_8 = stateReg == 4'h7;
	wire _GEN_9 = (_GEN | _GEN_0) | _GEN_1;
	wire _GEN_10 = _GEN_9 | ~_GEN_4;
	wire _GEN_11 = _GEN_4 | _GEN_5;
	wire [511:0] _GEN_12 = {64'hffffffffffffffff, currLen, procInterrupt, fifoHeadReg, fifoTailReg, maxLength, rAddr, rPause};
	always @(posedge clock)
		if (reset) begin
			rAddr <= 64'h0000000000000000;
			rPause <= 64'h0000000000000000;
			procInterrupt <= 64'h0000000000000000;
			maxLength <= 64'h0000000000000000;
			stateReg <= 4'h0;
			currLen <= 64'h0000000000000000;
			contentionCounter <= 64'h0000000000000000;
			networkCongested <= 1'h0;
			fifoTailReg <= 64'h0000000000000000;
			fifoHeadReg <= 64'h0000000000000000;
			memDataCounter <= 5'h00;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_13;
			reg _GEN_14;
			reg _GEN_15;
			reg [63:0] _GEN_16;
			reg _GEN_17;
			reg _GEN_18;
			reg _GEN_19;
			reg [63:0] _GEN_20;
			_GEN_19 = rPause == 64'h0000000000000000;
			_GEN_13 = stateReg == 4'h0;
			_GEN_14 = ((currLen == maxLength) & networkCongested) | (maxLength < (currLen + 64'h0000000000000010));
			_GEN_15 = io_write_data_ready & _GEN_2;
			_GEN_16 = maxLength - 64'h0000000000000001;
			_GEN_17 = _GEN_13 | _GEN_3;
			_GEN_18 = io_read_data_valid & _GEN_2;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h1))
				rAddr <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rAddr[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rAddr[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rAddr[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rAddr[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rAddr[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rAddr[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rAddr[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rAddr[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h0))
				rPause <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rPause[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rPause[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rPause[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rPause[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rPause[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rPause[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rPause[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rPause[7:0])};
			else if (_GEN_13 & (|procInterrupt | _GEN_14))
				rPause <= 64'hffffffffffffffff;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h5))
				procInterrupt <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : procInterrupt[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : procInterrupt[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : procInterrupt[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : procInterrupt[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : procInterrupt[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : procInterrupt[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : procInterrupt[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : procInterrupt[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h2))
				maxLength <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : maxLength[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : maxLength[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : maxLength[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : maxLength[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : maxLength[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : maxLength[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : maxLength[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : maxLength[7:0])};
			_GEN_20 = {stateReg, stateReg, stateReg, stateReg, stateReg, (_GEN_19 ? 4'h0 : 4'ha), (_GEN_19 ? 4'h0 : 4'h9), (io_connNetwork_ctrl_serveStealReq_ready ? 4'h7 : (networkCongested | (|procInterrupt) ? 4'h0 : stateReg)), (io_connNetwork_data_qOutTask_ready | networkCongested ? 4'h0 : 4'h7), (io_read_address_ready ? 4'h5 : stateReg), (_GEN_18 ? 4'h8 : stateReg), (io_write_address_ready ? 4'h3 : stateReg), (_GEN_15 ? 4'h0 : stateReg), ((_taskQueueBuffer_io_count == 5'h0f) & io_connNetwork_data_availableTask_valid ? 4'h4 : (io_connNetwork_data_availableTask_valid & networkCongested ? 4'h2 : (networkCongested ? stateReg : 4'h0))), stateReg, (|procInterrupt ? 4'ha : (_GEN_14 ? 4'h9 : (networkCongested & (_taskQueueBuffer_io_count == 5'h10) ? 4'h4 : (networkCongested ? 4'h2 : ((~networkCongested & |currLen) & ~(|_taskQueueBuffer_io_count) ? 4'h6 : (~networkCongested & |_taskQueueBuffer_io_count ? 4'h7 : stateReg))))))};
			stateReg <= _GEN_20[stateReg * 4+:4];
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h6))
				currLen <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : currLen[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : currLen[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : currLen[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : currLen[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : currLen[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : currLen[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : currLen[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : currLen[7:0])};
			else if (~_GEN_17) begin
				if (_GEN_1) begin
					if (_GEN_15)
						currLen <= currLen + 64'h0000000000000001;
					else if (io_write_data_ready)
						currLen <= currLen + 64'h0000000000000001;
				end
				else if (_GEN_4 | ~_GEN_5)
					;
				else if (_GEN_18)
					currLen <= currLen - 64'h0000000000000001;
				else if (io_read_data_valid)
					currLen <= currLen - 64'h0000000000000001;
			end
			if ((~io_connNetwork_ctrl_serveStealReq_ready & io_ntwDataUnitOccupancy) & (contentionCounter != 64'h0000000000000040))
				contentionCounter <= contentionCounter + 64'h0000000000000001;
			else if ((io_connNetwork_ctrl_serveStealReq_ready & |contentionCounter) & ~io_ntwDataUnitOccupancy)
				contentionCounter <= contentionCounter - 64'h0000000000000001;
			networkCongested <= (contentionCounter > 64'h0000000000000035) | ((contentionCounter > 64'h0000000000000033) & networkCongested);
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h3))
				fifoTailReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoTailReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoTailReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoTailReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoTailReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoTailReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoTailReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoTailReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoTailReg[7:0])};
			else if (_GEN_17 | ~_GEN_1)
				;
			else begin : sv2v_autoblock_2
				reg _GEN_21;
				_GEN_21 = fifoTailReg < _GEN_16;
				if (_GEN_15) begin
					if (_GEN_21)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
				else if (io_write_data_ready) begin
					if (_GEN_21)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
			end
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h4))
				fifoHeadReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoHeadReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoHeadReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoHeadReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoHeadReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoHeadReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoHeadReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoHeadReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoHeadReg[7:0])};
			else if ((_GEN_13 | _GEN_7) | ~_GEN_5)
				;
			else begin : sv2v_autoblock_3
				reg _GEN_22;
				_GEN_22 = fifoHeadReg < _GEN_16;
				if (_GEN_18) begin
					if (_GEN_22)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
				else if (io_read_data_valid) begin
					if (_GEN_22)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
			end
			if (~(_GEN_13 | _GEN)) begin
				if (_GEN_0) begin
					if (io_write_address_ready)
						memDataCounter <= 5'h10;
				end
				else if (_GEN_1) begin
					if (_GEN_15 | ~io_write_data_ready)
						;
					else
						memDataCounter <= memDataCounter - 5'h01;
				end
				else if (_GEN_4) begin
					if (io_read_address_ready)
						memDataCounter <= (currLen < 64'h0000000000000010 ? currLen[4:0] : 5'h10);
				end
				else if ((~_GEN_5 | _GEN_18) | ~io_read_data_valid)
					;
				else
					memDataCounter <= memDataCounter - 5'h01;
			end
		end
	Queue2_AddressChannel_2 s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_ar_ready),
		.io_enq_valid(io_axi_mgmt_ar_valid),
		.io_enq_bits_addr(io_axi_mgmt_ar_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_ar_bits_prot),
		.io_deq_ready(_rdReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_rdRespQueue__io_deq_valid),
		.io_enq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_enq_bits_resp(_rdRespQueue__io_deq_bits_resp),
		.io_deq_ready(io_axi_mgmt_r_ready),
		.io_deq_valid(io_axi_mgmt_r_valid),
		.io_deq_bits_data(io_axi_mgmt_r_bits_data),
		.io_deq_bits_resp(io_axi_mgmt_r_bits_resp)
	);
	Queue2_AddressChannel_2 s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_aw_ready),
		.io_enq_valid(io_axi_mgmt_aw_valid),
		.io_enq_bits_addr(io_axi_mgmt_aw_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_aw_bits_prot),
		.io_deq_ready(_wrReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_w_ready),
		.io_enq_valid(io_axi_mgmt_w_valid),
		.io_enq_bits_data(io_axi_mgmt_w_bits_data),
		.io_enq_bits_strb(io_axi_mgmt_w_bits_strb),
		.io_deq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_wrRespQueue__io_deq_valid),
		.io_enq_bits_resp(2'h0),
		.io_deq_ready(io_axi_mgmt_b_ready),
		.io_deq_valid(io_axi_mgmt_b_valid),
		.io_deq_bits_resp(io_axi_mgmt_b_bits_resp)
	);
	Queue1_AddressChannel rdReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_deq_ready(rdReq),
		.io_deq_valid(_rdReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_rdReq__deq_q_io_deq_bits_addr)
	);
	Queue1_ReadDataChannel rdRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdRespQueue__io_enq_ready),
		.io_enq_valid(rdReq),
		.io_enq_bits_data(_GEN_12[_rdReq__deq_q_io_deq_bits_addr[5:3] * 64+:64]),
		.io_deq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_deq_valid(_rdRespQueue__io_deq_valid),
		.io_deq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_deq_bits_resp(_rdRespQueue__io_deq_bits_resp)
	);
	Queue1_AddressChannel wrReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_wrReq__deq_q_io_deq_bits_addr)
	);
	Queue1_WriteDataChannel wrReqData__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_enq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_enq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReqData__deq_q_io_deq_valid),
		.io_deq_bits_data(_wrReqData__deq_q_io_deq_bits_data),
		.io_deq_bits_strb(_wrReqData__deq_q_io_deq_bits_strb)
	);
	Queue1_WriteResponseChannel wrRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrRespQueue__io_enq_ready),
		.io_enq_valid(wrReq),
		.io_deq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_deq_valid(_wrRespQueue__io_deq_valid)
	);
	Queue16_UInt taskQueueBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_taskQueueBuffer_io_enq_ready),
		.io_enq_valid((_GEN ? io_connNetwork_data_availableTask_valid : (~_GEN_6 & _GEN_5) & io_read_data_valid)),
		.io_enq_bits((_GEN ? io_connNetwork_data_availableTask_bits : (_GEN_6 | ~_GEN_5 ? 128'h00000000000000000000000000000000 : io_read_data_bits))),
		.io_deq_ready(~_GEN_3 & (_GEN_1 ? io_write_data_ready : (~_GEN_11 & _GEN_8) & io_connNetwork_data_qOutTask_ready)),
		.io_deq_bits(_taskQueueBuffer_io_deq_bits),
		.io_count(_taskQueueBuffer_io_count)
	);
	assign io_connNetwork_ctrl_serveStealReq_valid = ~(((((_GEN | _GEN_0) | _GEN_1) | _GEN_4) | _GEN_5) | _GEN_8) & (stateReg == 4'h8);
	assign io_connNetwork_data_availableTask_ready = _GEN & _taskQueueBuffer_io_enq_ready;
	assign io_connNetwork_data_qOutTask_valid = ~(((_GEN | _GEN_0) | _GEN_1) | _GEN_11) & _GEN_8;
	assign io_connNetwork_data_qOutTask_bits = _taskQueueBuffer_io_deq_bits;
	assign io_read_address_valid = ~_GEN_9 & _GEN_4;
	assign io_read_address_bits = (_GEN_10 ? 64'h0000000000000000 : {fifoHeadReg[59:0], 4'h0} + rAddr);
	assign io_read_data_ready = ~_GEN_7 & _GEN_5;
	assign io_read_burst_len = (_GEN_10 ? 4'h0 : (currLen < 64'h0000000000000010 ? currLen[3:0] - 4'h1 : 4'hf));
	assign io_write_address_valid = ~_GEN & _GEN_0;
	assign io_write_address_bits = (_GEN | ~_GEN_0 ? 64'h0000000000000000 : {fifoTailReg[59:0], 4'h0} + rAddr);
	assign io_write_data_valid = ~_GEN_3 & _GEN_1;
	assign io_write_data_bits = _taskQueueBuffer_io_deq_bits;
	assign io_write_burst_len = (_GEN ? 4'h0 : {4 {_GEN_0}});
	assign io_write_last = (~_GEN_3 & _GEN_1) & _GEN_2;
endmodule
module RVtoAXIBridge (
	clock,
	reset,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_writeBurst_len,
	io_writeBurst_last,
	io_readBurst_len,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_ar_bits_len,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data,
	axi_aw_ready,
	axi_aw_valid,
	axi_aw_bits_addr,
	axi_aw_bits_len,
	axi_w_ready,
	axi_w_valid,
	axi_w_bits_data,
	axi_w_bits_last,
	axi_b_valid
);
	input clock;
	input reset;
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [127:0] io_read_data_bits;
	output wire io_write_address_ready;
	input io_write_address_valid;
	input [63:0] io_write_address_bits;
	output wire io_write_data_ready;
	input io_write_data_valid;
	input [127:0] io_write_data_bits;
	input [3:0] io_writeBurst_len;
	input io_writeBurst_last;
	input [3:0] io_readBurst_len;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire [7:0] axi_ar_bits_len;
	output wire axi_r_ready;
	input axi_r_valid;
	input [127:0] axi_r_bits_data;
	input axi_aw_ready;
	output wire axi_aw_valid;
	output wire [63:0] axi_aw_bits_addr;
	output wire [7:0] axi_aw_bits_len;
	input axi_w_ready;
	output wire axi_w_valid;
	output wire [127:0] axi_w_bits_data;
	output wire axi_w_bits_last;
	input axi_b_valid;
	reg writeHandshakeDetector;
	wire axi_w_valid_0 = (io_write_data_valid & axi_w_ready) & ~writeHandshakeDetector;
	always @(posedge clock)
		if (reset)
			writeHandshakeDetector <= 1'h0;
		else if (axi_w_valid_0)
			writeHandshakeDetector <= io_writeBurst_last | writeHandshakeDetector;
		else
			writeHandshakeDetector <= ~axi_b_valid & writeHandshakeDetector;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign io_write_address_ready = axi_aw_ready;
	assign io_write_data_ready = axi_w_ready & ~writeHandshakeDetector;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_ar_bits_len = {4'h0, io_readBurst_len};
	assign axi_r_ready = io_read_data_ready;
	assign axi_aw_valid = io_write_address_valid;
	assign axi_aw_bits_addr = io_write_address_bits;
	assign axi_aw_bits_len = {4'h0, io_writeBurst_len};
	assign axi_w_valid = axi_w_valid_0;
	assign axi_w_bits_data = io_write_data_bits;
	assign axi_w_bits_last = io_writeBurst_last;
endmodule
module Queue1_ReadAddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	reg [93:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, 1'h0};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_id = ram[0];
	assign io_deq_bits_addr = ram[64:1];
	assign io_deq_bits_len = ram[72:65];
	assign io_deq_bits_size = ram[75:73];
	assign io_deq_bits_burst = ram[77:76];
	assign io_deq_bits_lock = ram[78];
	assign io_deq_bits_cache = ram[82:79];
	assign io_deq_bits_prot = ram[85:83];
	assign io_deq_bits_qos = ram[89:86];
	assign io_deq_bits_region = ram[93:90];
endmodule
module Queue1_ReadDataChannel_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits_id;
	input [127:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [127:0] io_deq_bits_data;
	reg [131:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_last, io_enq_bits_resp, io_enq_bits_data, io_enq_bits_id};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[128:1];
endmodule
module Queue1_WriteAddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	reg [93:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, 1'h0};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_id = ram[0];
	assign io_deq_bits_addr = ram[64:1];
	assign io_deq_bits_len = ram[72:65];
	assign io_deq_bits_size = ram[75:73];
	assign io_deq_bits_burst = ram[77:76];
	assign io_deq_bits_lock = ram[78];
	assign io_deq_bits_cache = ram[82:79];
	assign io_deq_bits_prot = ram[85:83];
	assign io_deq_bits_qos = ram[89:86];
	assign io_deq_bits_region = ram[93:90];
endmodule
module Queue1_WriteDataChannel_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [127:0] io_enq_bits_data;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [127:0] io_deq_bits_data;
	output wire [15:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	reg [144:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_last, 16'hffff, io_enq_bits_data};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[127:0];
	assign io_deq_bits_strb = ram[143:128];
	assign io_deq_bits_last = ram[144];
endmodule
module Queue1_WriteResponseChannel_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_deq_valid
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	output wire io_deq_valid;
	reg full;
	always @(posedge clock)
		if (reset)
			full <= 1'h0;
		else begin : sv2v_autoblock_1
			reg do_enq;
			do_enq = ~full & io_enq_valid;
			if (~(do_enq == full))
				full <= do_enq;
		end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
endmodule
module ram_2x95 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [94:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [94:0] W0_data;
	reg [94:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 95'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadAddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_id;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [94:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x95 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[1:0];
	assign io_deq_bits_addr = _ram_ext_R0_data[65:2];
	assign io_deq_bits_len = _ram_ext_R0_data[73:66];
	assign io_deq_bits_size = _ram_ext_R0_data[76:74];
	assign io_deq_bits_burst = _ram_ext_R0_data[78:77];
	assign io_deq_bits_lock = _ram_ext_R0_data[79];
	assign io_deq_bits_cache = _ram_ext_R0_data[83:80];
	assign io_deq_bits_prot = _ram_ext_R0_data[86:84];
	assign io_deq_bits_qos = _ram_ext_R0_data[90:87];
	assign io_deq_bits_region = _ram_ext_R0_data[94:91];
endmodule
module ram_2x133 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [132:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [132:0] W0_data;
	reg [132:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 133'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel_3 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_data,
	io_deq_bits_resp,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_id;
	input [127:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_id;
	output wire [127:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	output wire io_deq_bits_last;
	wire [132:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x133 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_resp, io_enq_bits_data, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[1:0];
	assign io_deq_bits_data = _ram_ext_R0_data[129:2];
	assign io_deq_bits_resp = _ram_ext_R0_data[131:130];
	assign io_deq_bits_last = _ram_ext_R0_data[132];
endmodule
module Queue2_WriteAddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_id;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [94:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x95 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[1:0];
	assign io_deq_bits_addr = _ram_ext_R0_data[65:2];
	assign io_deq_bits_len = _ram_ext_R0_data[73:66];
	assign io_deq_bits_size = _ram_ext_R0_data[76:74];
	assign io_deq_bits_burst = _ram_ext_R0_data[78:77];
	assign io_deq_bits_lock = _ram_ext_R0_data[79];
	assign io_deq_bits_cache = _ram_ext_R0_data[83:80];
	assign io_deq_bits_prot = _ram_ext_R0_data[86:84];
	assign io_deq_bits_qos = _ram_ext_R0_data[90:87];
	assign io_deq_bits_region = _ram_ext_R0_data[94:91];
endmodule
module ram_2x145 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [144:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [144:0] W0_data;
	reg [144:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 145'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteDataChannel_3 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [127:0] io_enq_bits_data;
	input [15:0] io_enq_bits_strb;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [127:0] io_deq_bits_data;
	output wire [15:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	wire [144:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x145 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_strb, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[127:0];
	assign io_deq_bits_strb = _ram_ext_R0_data[143:128];
	assign io_deq_bits_last = _ram_ext_R0_data[144];
endmodule
module Queue2_WriteResponseChannel_3 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_id;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_id;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x2 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_id),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_id)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module elasticArbiter (
	clock,
	reset,
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_id,
	io_sources_0_bits_addr,
	io_sources_0_bits_len,
	io_sources_0_bits_size,
	io_sources_0_bits_burst,
	io_sources_0_bits_lock,
	io_sources_0_bits_cache,
	io_sources_0_bits_prot,
	io_sources_0_bits_qos,
	io_sources_0_bits_region,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_id,
	io_sources_1_bits_addr,
	io_sources_1_bits_len,
	io_sources_1_bits_size,
	io_sources_1_bits_burst,
	io_sources_1_bits_lock,
	io_sources_1_bits_cache,
	io_sources_1_bits_prot,
	io_sources_1_bits_qos,
	io_sources_1_bits_region,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_id,
	io_sink_bits_addr,
	io_sink_bits_len,
	io_sink_bits_size,
	io_sink_bits_burst,
	io_sink_bits_lock,
	io_sink_bits_cache,
	io_sink_bits_prot,
	io_sink_bits_qos,
	io_sink_bits_region,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	input clock;
	input reset;
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [1:0] io_sources_0_bits_id;
	input [63:0] io_sources_0_bits_addr;
	input [7:0] io_sources_0_bits_len;
	input [2:0] io_sources_0_bits_size;
	input [1:0] io_sources_0_bits_burst;
	input io_sources_0_bits_lock;
	input [3:0] io_sources_0_bits_cache;
	input [2:0] io_sources_0_bits_prot;
	input [3:0] io_sources_0_bits_qos;
	input [3:0] io_sources_0_bits_region;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [1:0] io_sources_1_bits_id;
	input [63:0] io_sources_1_bits_addr;
	input [7:0] io_sources_1_bits_len;
	input [2:0] io_sources_1_bits_size;
	input [1:0] io_sources_1_bits_burst;
	input io_sources_1_bits_lock;
	input [3:0] io_sources_1_bits_cache;
	input [2:0] io_sources_1_bits_prot;
	input [3:0] io_sources_1_bits_qos;
	input [3:0] io_sources_1_bits_region;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [1:0] io_sink_bits_id;
	output wire [63:0] io_sink_bits_addr;
	output wire [7:0] io_sink_bits_len;
	output wire [2:0] io_sink_bits_size;
	output wire [1:0] io_sink_bits_burst;
	output wire io_sink_bits_lock;
	output wire [3:0] io_sink_bits_cache;
	output wire [2:0] io_sink_bits_prot;
	output wire [3:0] io_sink_bits_qos;
	output wire [3:0] io_sink_bits_region;
	input io_select_ready;
	output wire io_select_valid;
	output wire io_select_bits;
	wire sourceReady;
	reg chooser_lastChoice;
	wire _GEN = (chooser_lastChoice ? io_sources_0_valid : io_sources_1_valid);
	wire io_select_bits_0 = (_GEN ? ~chooser_lastChoice : ~io_sources_0_valid);
	wire _GEN_0 = (io_select_bits_0 ? io_sources_1_valid : io_sources_0_valid);
	reg sinkSent;
	reg selectSent;
	assign sourceReady = (sinkSent | io_sink_ready) & (selectSent | io_select_ready);
	always @(posedge clock)
		if (reset) begin
			chooser_lastChoice <= 1'h0;
			sinkSent <= 1'h0;
			selectSent <= 1'h0;
		end
		else begin
			if (_GEN_0 & sourceReady) begin
				if (_GEN)
					chooser_lastChoice <= ~chooser_lastChoice;
				else
					chooser_lastChoice <= ~io_sources_0_valid;
			end
			sinkSent <= ((io_sink_ready | sinkSent) & _GEN_0) & ~sourceReady;
			selectSent <= ((io_select_ready | selectSent) & _GEN_0) & ~sourceReady;
		end
	assign io_sources_0_ready = sourceReady & ~io_select_bits_0;
	assign io_sources_1_ready = sourceReady & io_select_bits_0;
	assign io_sink_valid = _GEN_0 & ~sinkSent;
	assign io_sink_bits_id = (io_select_bits_0 ? io_sources_1_bits_id : io_sources_0_bits_id);
	assign io_sink_bits_addr = (io_select_bits_0 ? io_sources_1_bits_addr : io_sources_0_bits_addr);
	assign io_sink_bits_len = (io_select_bits_0 ? io_sources_1_bits_len : io_sources_0_bits_len);
	assign io_sink_bits_size = (io_select_bits_0 ? io_sources_1_bits_size : io_sources_0_bits_size);
	assign io_sink_bits_burst = (io_select_bits_0 ? io_sources_1_bits_burst : io_sources_0_bits_burst);
	assign io_sink_bits_lock = (io_select_bits_0 ? io_sources_1_bits_lock : io_sources_0_bits_lock);
	assign io_sink_bits_cache = (io_select_bits_0 ? io_sources_1_bits_cache : io_sources_0_bits_cache);
	assign io_sink_bits_prot = (io_select_bits_0 ? io_sources_1_bits_prot : io_sources_0_bits_prot);
	assign io_sink_bits_qos = (io_select_bits_0 ? io_sources_1_bits_qos : io_sources_0_bits_qos);
	assign io_sink_bits_region = (io_select_bits_0 ? io_sources_1_bits_region : io_sources_0_bits_region);
	assign io_select_valid = _GEN_0 & ~selectSent;
	assign io_select_bits = io_select_bits_0;
endmodule
module elasticDemux_3 (
	io_source_ready,
	io_source_valid,
	io_source_bits_id,
	io_source_bits_data,
	io_source_bits_resp,
	io_source_bits_last,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_id,
	io_sinks_0_bits_data,
	io_sinks_0_bits_resp,
	io_sinks_0_bits_last,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_id,
	io_sinks_1_bits_data,
	io_sinks_1_bits_resp,
	io_sinks_1_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [1:0] io_source_bits_id;
	input [127:0] io_source_bits_data;
	input [1:0] io_source_bits_resp;
	input io_source_bits_last;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [1:0] io_sinks_0_bits_id;
	output wire [127:0] io_sinks_0_bits_data;
	output wire [1:0] io_sinks_0_bits_resp;
	output wire io_sinks_0_bits_last;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [1:0] io_sinks_1_bits_id;
	output wire [127:0] io_sinks_1_bits_data;
	output wire [1:0] io_sinks_1_bits_resp;
	output wire io_sinks_1_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire fire = valid & (io_select_bits ? io_sinks_1_ready : io_sinks_0_ready);
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & ~io_select_bits;
	assign io_sinks_0_bits_id = io_source_bits_id;
	assign io_sinks_0_bits_data = io_source_bits_data;
	assign io_sinks_0_bits_resp = io_source_bits_resp;
	assign io_sinks_0_bits_last = io_source_bits_last;
	assign io_sinks_1_valid = valid & io_select_bits;
	assign io_sinks_1_bits_id = io_source_bits_id;
	assign io_sinks_1_bits_data = io_source_bits_data;
	assign io_sinks_1_bits_resp = io_source_bits_resp;
	assign io_sinks_1_bits_last = io_source_bits_last;
	assign io_select_ready = fire;
endmodule
module ram_32x1 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [4:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire R0_data;
	input [4:0] W0_addr;
	input W0_en;
	input W0_clk;
	input W0_data;
	reg Memory [0:31];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 1'bx);
endmodule
module Queue32_UInt1 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits;
	wire io_enq_ready_0;
	wire _ram_ext_R0_data;
	reg [4:0] enq_ptr_value;
	reg [4:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire io_deq_valid_0 = io_enq_valid | ~empty;
	wire do_deq = (~empty & io_deq_ready) & io_deq_valid_0;
	wire do_enq = (~(empty & io_deq_ready) & io_enq_ready_0) & io_enq_valid;
	assign io_enq_ready_0 = io_deq_ready | ~(ptr_match & maybe_full);
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 5'h00;
			deq_ptr_value <= 5'h00;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 5'h01;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 5'h01;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_32x1 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = io_enq_ready_0;
	assign io_deq_valid = io_deq_valid_0;
	assign io_deq_bits = (empty ? io_enq_bits : _ram_ext_R0_data);
endmodule
module elasticMux_2 (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_data,
	io_sources_0_bits_strb,
	io_sources_0_bits_last,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_data,
	io_sources_1_bits_strb,
	io_sources_1_bits_last,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_data,
	io_sink_bits_strb,
	io_sink_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [127:0] io_sources_0_bits_data;
	input [15:0] io_sources_0_bits_strb;
	input io_sources_0_bits_last;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [127:0] io_sources_1_bits_data;
	input [15:0] io_sources_1_bits_strb;
	input io_sources_1_bits_last;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [127:0] io_sink_bits_data;
	output wire [15:0] io_sink_bits_strb;
	output wire io_sink_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input io_select_bits;
	wire io_sink_bits_last_0 = (io_select_bits ? io_sources_1_bits_last : io_sources_0_bits_last);
	wire valid = io_select_valid & (io_select_bits ? io_sources_1_valid : io_sources_0_valid);
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & ~io_select_bits;
	assign io_sources_1_ready = fire & io_select_bits;
	assign io_sink_valid = valid;
	assign io_sink_bits_data = (io_select_bits ? io_sources_1_bits_data : io_sources_0_bits_data);
	assign io_sink_bits_strb = (io_select_bits ? io_sources_1_bits_strb : io_sources_0_bits_strb);
	assign io_sink_bits_last = io_sink_bits_last_0;
	assign io_select_ready = fire & io_sink_bits_last_0;
endmodule
module elasticDemux_4 (
	io_source_ready,
	io_source_valid,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire io_select_ready;
	input io_select_valid;
	input io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire fire = valid & (io_select_bits ? io_sinks_1_ready : io_sinks_0_ready);
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & ~io_select_bits;
	assign io_sinks_1_valid = valid & io_select_bits;
	assign io_select_ready = fire;
endmodule
module axi4FullMux (
	clock,
	reset,
	s_axi_0_ar_ready,
	s_axi_0_ar_valid,
	s_axi_0_ar_bits_addr,
	s_axi_0_ar_bits_len,
	s_axi_0_ar_bits_size,
	s_axi_0_ar_bits_burst,
	s_axi_0_ar_bits_lock,
	s_axi_0_ar_bits_cache,
	s_axi_0_ar_bits_prot,
	s_axi_0_ar_bits_qos,
	s_axi_0_ar_bits_region,
	s_axi_0_r_ready,
	s_axi_0_r_valid,
	s_axi_0_r_bits_data,
	s_axi_0_aw_ready,
	s_axi_0_aw_valid,
	s_axi_0_aw_bits_addr,
	s_axi_0_aw_bits_len,
	s_axi_0_aw_bits_size,
	s_axi_0_aw_bits_burst,
	s_axi_0_aw_bits_lock,
	s_axi_0_aw_bits_cache,
	s_axi_0_aw_bits_prot,
	s_axi_0_aw_bits_qos,
	s_axi_0_aw_bits_region,
	s_axi_0_w_ready,
	s_axi_0_w_valid,
	s_axi_0_w_bits_data,
	s_axi_0_w_bits_last,
	s_axi_0_b_valid,
	s_axi_1_ar_ready,
	s_axi_1_ar_valid,
	s_axi_1_ar_bits_addr,
	s_axi_1_ar_bits_len,
	s_axi_1_ar_bits_size,
	s_axi_1_ar_bits_burst,
	s_axi_1_ar_bits_lock,
	s_axi_1_ar_bits_cache,
	s_axi_1_ar_bits_prot,
	s_axi_1_ar_bits_qos,
	s_axi_1_ar_bits_region,
	s_axi_1_r_ready,
	s_axi_1_r_valid,
	s_axi_1_r_bits_data,
	s_axi_1_aw_ready,
	s_axi_1_aw_valid,
	s_axi_1_aw_bits_addr,
	s_axi_1_aw_bits_len,
	s_axi_1_aw_bits_size,
	s_axi_1_aw_bits_burst,
	s_axi_1_aw_bits_lock,
	s_axi_1_aw_bits_cache,
	s_axi_1_aw_bits_prot,
	s_axi_1_aw_bits_qos,
	s_axi_1_aw_bits_region,
	s_axi_1_w_ready,
	s_axi_1_w_valid,
	s_axi_1_w_bits_data,
	s_axi_1_w_bits_last,
	s_axi_1_b_valid,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_id,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_id,
	m_axi_r_bits_data,
	m_axi_r_bits_resp,
	m_axi_r_bits_last,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_id,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_strb,
	m_axi_w_bits_last,
	m_axi_b_ready,
	m_axi_b_valid,
	m_axi_b_bits_id,
	m_axi_b_bits_resp
);
	input clock;
	input reset;
	output wire s_axi_0_ar_ready;
	input s_axi_0_ar_valid;
	input [63:0] s_axi_0_ar_bits_addr;
	input [7:0] s_axi_0_ar_bits_len;
	input [2:0] s_axi_0_ar_bits_size;
	input [1:0] s_axi_0_ar_bits_burst;
	input s_axi_0_ar_bits_lock;
	input [3:0] s_axi_0_ar_bits_cache;
	input [2:0] s_axi_0_ar_bits_prot;
	input [3:0] s_axi_0_ar_bits_qos;
	input [3:0] s_axi_0_ar_bits_region;
	input s_axi_0_r_ready;
	output wire s_axi_0_r_valid;
	output wire [127:0] s_axi_0_r_bits_data;
	output wire s_axi_0_aw_ready;
	input s_axi_0_aw_valid;
	input [63:0] s_axi_0_aw_bits_addr;
	input [7:0] s_axi_0_aw_bits_len;
	input [2:0] s_axi_0_aw_bits_size;
	input [1:0] s_axi_0_aw_bits_burst;
	input s_axi_0_aw_bits_lock;
	input [3:0] s_axi_0_aw_bits_cache;
	input [2:0] s_axi_0_aw_bits_prot;
	input [3:0] s_axi_0_aw_bits_qos;
	input [3:0] s_axi_0_aw_bits_region;
	output wire s_axi_0_w_ready;
	input s_axi_0_w_valid;
	input [127:0] s_axi_0_w_bits_data;
	input s_axi_0_w_bits_last;
	output wire s_axi_0_b_valid;
	output wire s_axi_1_ar_ready;
	input s_axi_1_ar_valid;
	input [63:0] s_axi_1_ar_bits_addr;
	input [7:0] s_axi_1_ar_bits_len;
	input [2:0] s_axi_1_ar_bits_size;
	input [1:0] s_axi_1_ar_bits_burst;
	input s_axi_1_ar_bits_lock;
	input [3:0] s_axi_1_ar_bits_cache;
	input [2:0] s_axi_1_ar_bits_prot;
	input [3:0] s_axi_1_ar_bits_qos;
	input [3:0] s_axi_1_ar_bits_region;
	input s_axi_1_r_ready;
	output wire s_axi_1_r_valid;
	output wire [127:0] s_axi_1_r_bits_data;
	output wire s_axi_1_aw_ready;
	input s_axi_1_aw_valid;
	input [63:0] s_axi_1_aw_bits_addr;
	input [7:0] s_axi_1_aw_bits_len;
	input [2:0] s_axi_1_aw_bits_size;
	input [1:0] s_axi_1_aw_bits_burst;
	input s_axi_1_aw_bits_lock;
	input [3:0] s_axi_1_aw_bits_cache;
	input [2:0] s_axi_1_aw_bits_prot;
	input [3:0] s_axi_1_aw_bits_qos;
	input [3:0] s_axi_1_aw_bits_region;
	output wire s_axi_1_w_ready;
	input s_axi_1_w_valid;
	input [127:0] s_axi_1_w_bits_data;
	input s_axi_1_w_bits_last;
	output wire s_axi_1_b_valid;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [1:0] m_axi_ar_bits_id;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [1:0] m_axi_r_bits_id;
	input [127:0] m_axi_r_bits_data;
	input [1:0] m_axi_r_bits_resp;
	input m_axi_r_bits_last;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [1:0] m_axi_aw_bits_id;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [127:0] m_axi_w_bits_data;
	output wire [15:0] m_axi_w_bits_strb;
	output wire m_axi_w_bits_last;
	output wire m_axi_b_ready;
	input m_axi_b_valid;
	input [1:0] m_axi_b_bits_id;
	input [1:0] m_axi_b_bits_resp;
	wire _write_demux_io_source_ready;
	wire _write_demux_io_sinks_0_valid;
	wire _write_demux_io_sinks_1_valid;
	wire _write_demux_io_select_ready;
	wire _write_mux_io_sources_0_ready;
	wire _write_mux_io_sources_1_ready;
	wire _write_mux_io_sink_valid;
	wire [127:0] _write_mux_io_sink_bits_data;
	wire [15:0] _write_mux_io_sink_bits_strb;
	wire _write_mux_io_sink_bits_last;
	wire _write_mux_io_select_ready;
	wire _write_arbiter_io_sources_0_ready;
	wire _write_arbiter_io_sources_1_ready;
	wire _write_arbiter_io_sink_valid;
	wire [1:0] _write_arbiter_io_sink_bits_id;
	wire [63:0] _write_arbiter_io_sink_bits_addr;
	wire [7:0] _write_arbiter_io_sink_bits_len;
	wire [2:0] _write_arbiter_io_sink_bits_size;
	wire [1:0] _write_arbiter_io_sink_bits_burst;
	wire _write_arbiter_io_sink_bits_lock;
	wire [3:0] _write_arbiter_io_sink_bits_cache;
	wire [2:0] _write_arbiter_io_sink_bits_prot;
	wire [3:0] _write_arbiter_io_sink_bits_qos;
	wire [3:0] _write_arbiter_io_sink_bits_region;
	wire _write_arbiter_io_select_valid;
	wire _write_arbiter_io_select_bits;
	wire _write_portQueue_io_enq_ready;
	wire _write_portQueue_io_deq_valid;
	wire _write_portQueue_io_deq_bits;
	wire _read_demux_io_source_ready;
	wire _read_demux_io_sinks_0_valid;
	wire [1:0] _read_demux_io_sinks_0_bits_id;
	wire [127:0] _read_demux_io_sinks_0_bits_data;
	wire [1:0] _read_demux_io_sinks_0_bits_resp;
	wire _read_demux_io_sinks_0_bits_last;
	wire _read_demux_io_sinks_1_valid;
	wire [1:0] _read_demux_io_sinks_1_bits_id;
	wire [127:0] _read_demux_io_sinks_1_bits_data;
	wire [1:0] _read_demux_io_sinks_1_bits_resp;
	wire _read_demux_io_sinks_1_bits_last;
	wire _read_demux_io_select_ready;
	wire _read_arbiter_io_sources_0_ready;
	wire _read_arbiter_io_sources_1_ready;
	wire _read_arbiter_io_sink_valid;
	wire [1:0] _read_arbiter_io_sink_bits_id;
	wire [63:0] _read_arbiter_io_sink_bits_addr;
	wire [7:0] _read_arbiter_io_sink_bits_len;
	wire [2:0] _read_arbiter_io_sink_bits_size;
	wire [1:0] _read_arbiter_io_sink_bits_burst;
	wire _read_arbiter_io_sink_bits_lock;
	wire [3:0] _read_arbiter_io_sink_bits_cache;
	wire [2:0] _read_arbiter_io_sink_bits_prot;
	wire [3:0] _read_arbiter_io_sink_bits_qos;
	wire [3:0] _read_arbiter_io_sink_bits_region;
	wire _m_axi__sinkBuffer_1_io_deq_valid;
	wire [1:0] _m_axi__sinkBuffer_1_io_deq_bits_id;
	wire _m_axi__sourceBuffer_2_io_enq_ready;
	wire _m_axi__sourceBuffer_1_io_enq_ready;
	wire _m_axi__sinkBuffer_io_deq_valid;
	wire [1:0] _m_axi__sinkBuffer_io_deq_bits_id;
	wire [127:0] _m_axi__sinkBuffer_io_deq_bits_data;
	wire [1:0] _m_axi__sinkBuffer_io_deq_bits_resp;
	wire _m_axi__sinkBuffer_io_deq_bits_last;
	wire _m_axi__sourceBuffer_io_enq_ready;
	wire _s_axi__buffered_sinkBuffer_3_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_valid;
	wire [127:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_data;
	wire [15:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_2_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_1_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_valid;
	wire [127:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_data;
	wire [15:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_region;
	reg read_eagerFork_regs_0;
	reg read_eagerFork_regs_1;
	wire read_eagerFork_m_axi__r_ready_qual1_0 = _read_demux_io_source_ready | read_eagerFork_regs_0;
	wire read_eagerFork_m_axi__r_ready_qual1_1 = _read_demux_io_select_ready | read_eagerFork_regs_1;
	wire m_axi__r_ready = read_eagerFork_m_axi__r_ready_qual1_0 & read_eagerFork_m_axi__r_ready_qual1_1;
	reg write_eagerFork_regs_0;
	reg write_eagerFork_regs_1;
	wire write_eagerFork_m_axi__b_ready_qual1_0 = _write_demux_io_source_ready | write_eagerFork_regs_0;
	wire write_eagerFork_m_axi__b_ready_qual1_1 = _write_demux_io_select_ready | write_eagerFork_regs_1;
	wire m_axi__b_ready = write_eagerFork_m_axi__b_ready_qual1_0 & write_eagerFork_m_axi__b_ready_qual1_1;
	always @(posedge clock)
		if (reset) begin
			read_eagerFork_regs_0 <= 1'h0;
			read_eagerFork_regs_1 <= 1'h0;
			write_eagerFork_regs_0 <= 1'h0;
			write_eagerFork_regs_1 <= 1'h0;
		end
		else begin
			read_eagerFork_regs_0 <= (read_eagerFork_m_axi__r_ready_qual1_0 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			read_eagerFork_regs_1 <= (read_eagerFork_m_axi__r_ready_qual1_1 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			write_eagerFork_regs_0 <= (write_eagerFork_m_axi__b_ready_qual1_0 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
			write_eagerFork_regs_1 <= (write_eagerFork_m_axi__b_ready_qual1_1 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
		end
	Queue1_ReadAddressChannel s_axi__buffered_sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_ar_ready),
		.io_enq_valid(s_axi_0_ar_valid),
		.io_enq_bits_addr(s_axi_0_ar_bits_addr),
		.io_enq_bits_len(s_axi_0_ar_bits_len),
		.io_enq_bits_size(s_axi_0_ar_bits_size),
		.io_enq_bits_burst(s_axi_0_ar_bits_burst),
		.io_enq_bits_lock(s_axi_0_ar_bits_lock),
		.io_enq_bits_cache(s_axi_0_ar_bits_cache),
		.io_enq_bits_prot(s_axi_0_ar_bits_prot),
		.io_enq_bits_qos(s_axi_0_ar_bits_qos),
		.io_enq_bits_region(s_axi_0_ar_bits_region),
		.io_deq_ready(_read_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region)
	);
	Queue1_ReadDataChannel_2 s_axi__buffered_sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_0_valid),
		.io_enq_bits_id(_read_demux_io_sinks_0_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_deq_ready(s_axi_0_r_ready),
		.io_deq_valid(s_axi_0_r_valid),
		.io_deq_bits_data(s_axi_0_r_bits_data)
	);
	Queue1_WriteAddressChannel s_axi__buffered_sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_aw_ready),
		.io_enq_valid(s_axi_0_aw_valid),
		.io_enq_bits_addr(s_axi_0_aw_bits_addr),
		.io_enq_bits_len(s_axi_0_aw_bits_len),
		.io_enq_bits_size(s_axi_0_aw_bits_size),
		.io_enq_bits_burst(s_axi_0_aw_bits_burst),
		.io_enq_bits_lock(s_axi_0_aw_bits_lock),
		.io_enq_bits_cache(s_axi_0_aw_bits_cache),
		.io_enq_bits_prot(s_axi_0_aw_bits_prot),
		.io_enq_bits_qos(s_axi_0_aw_bits_qos),
		.io_enq_bits_region(s_axi_0_aw_bits_region),
		.io_deq_ready(_write_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_1_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region)
	);
	Queue1_WriteDataChannel_2 s_axi__buffered_sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_w_ready),
		.io_enq_valid(s_axi_0_w_valid),
		.io_enq_bits_data(s_axi_0_w_bits_data),
		.io_enq_bits_last(s_axi_0_w_bits_last),
		.io_deq_ready(_write_mux_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last)
	);
	Queue1_WriteResponseChannel_2 s_axi__buffered_sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_0_valid),
		.io_deq_valid(s_axi_0_b_valid)
	);
	Queue1_ReadAddressChannel s_axi__buffered_sourceBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_ar_ready),
		.io_enq_valid(s_axi_1_ar_valid),
		.io_enq_bits_addr(s_axi_1_ar_bits_addr),
		.io_enq_bits_len(s_axi_1_ar_bits_len),
		.io_enq_bits_size(s_axi_1_ar_bits_size),
		.io_enq_bits_burst(s_axi_1_ar_bits_burst),
		.io_enq_bits_lock(s_axi_1_ar_bits_lock),
		.io_enq_bits_cache(s_axi_1_ar_bits_cache),
		.io_enq_bits_prot(s_axi_1_ar_bits_prot),
		.io_enq_bits_qos(s_axi_1_ar_bits_qos),
		.io_enq_bits_region(s_axi_1_ar_bits_region),
		.io_deq_ready(_read_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_3_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region)
	);
	Queue1_ReadDataChannel_2 s_axi__buffered_sinkBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_1_valid),
		.io_enq_bits_id(_read_demux_io_sinks_1_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_deq_ready(s_axi_1_r_ready),
		.io_deq_valid(s_axi_1_r_valid),
		.io_deq_bits_data(s_axi_1_r_bits_data)
	);
	Queue1_WriteAddressChannel s_axi__buffered_sourceBuffer_4(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_aw_ready),
		.io_enq_valid(s_axi_1_aw_valid),
		.io_enq_bits_addr(s_axi_1_aw_bits_addr),
		.io_enq_bits_len(s_axi_1_aw_bits_len),
		.io_enq_bits_size(s_axi_1_aw_bits_size),
		.io_enq_bits_burst(s_axi_1_aw_bits_burst),
		.io_enq_bits_lock(s_axi_1_aw_bits_lock),
		.io_enq_bits_cache(s_axi_1_aw_bits_cache),
		.io_enq_bits_prot(s_axi_1_aw_bits_prot),
		.io_enq_bits_qos(s_axi_1_aw_bits_qos),
		.io_enq_bits_region(s_axi_1_aw_bits_region),
		.io_deq_ready(_write_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_4_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region)
	);
	Queue1_WriteDataChannel_2 s_axi__buffered_sourceBuffer_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_w_ready),
		.io_enq_valid(s_axi_1_w_valid),
		.io_enq_bits_data(s_axi_1_w_bits_data),
		.io_enq_bits_last(s_axi_1_w_bits_last),
		.io_deq_ready(_write_mux_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last)
	);
	Queue1_WriteResponseChannel_2 s_axi__buffered_sinkBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_1_valid),
		.io_deq_valid(s_axi_1_b_valid)
	);
	Queue2_ReadAddressChannel m_axi__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_enq_valid(_read_arbiter_io_sink_valid),
		.io_enq_bits_id(_read_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_read_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_read_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_read_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_id(m_axi_ar_bits_id),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	Queue2_ReadDataChannel_3 m_axi__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_r_ready),
		.io_enq_valid(m_axi_r_valid),
		.io_enq_bits_id(m_axi_r_bits_id),
		.io_enq_bits_data(m_axi_r_bits_data),
		.io_enq_bits_resp(m_axi_r_bits_resp),
		.io_enq_bits_last(m_axi_r_bits_last),
		.io_deq_ready(m_axi__r_ready),
		.io_deq_valid(_m_axi__sinkBuffer_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_deq_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_deq_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_deq_bits_last(_m_axi__sinkBuffer_io_deq_bits_last)
	);
	Queue2_WriteAddressChannel m_axi__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_sink_valid),
		.io_enq_bits_id(_write_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_write_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_write_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_write_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_id(m_axi_aw_bits_id),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_WriteDataChannel_3 m_axi__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_enq_valid(_write_mux_io_sink_valid),
		.io_enq_bits_data(_write_mux_io_sink_bits_data),
		.io_enq_bits_strb(_write_mux_io_sink_bits_strb),
		.io_enq_bits_last(_write_mux_io_sink_bits_last),
		.io_deq_ready(m_axi_w_ready),
		.io_deq_valid(m_axi_w_valid),
		.io_deq_bits_data(m_axi_w_bits_data),
		.io_deq_bits_strb(m_axi_w_bits_strb),
		.io_deq_bits_last(m_axi_w_bits_last)
	);
	Queue2_WriteResponseChannel_3 m_axi__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_b_ready),
		.io_enq_valid(m_axi_b_valid),
		.io_enq_bits_id(m_axi_b_bits_id),
		.io_enq_bits_resp(m_axi_b_bits_resp),
		.io_deq_ready(m_axi__b_ready),
		.io_deq_valid(_m_axi__sinkBuffer_1_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_1_io_deq_bits_id)
	);
	elasticArbiter read_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_read_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_sources_0_bits_id({1'h0, _s_axi__buffered_sourceBuffer_io_deq_bits_id}),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region),
		.io_sources_1_ready(_read_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_sources_1_bits_id({1'h1, _s_axi__buffered_sourceBuffer_3_io_deq_bits_id}),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_sink_valid(_read_arbiter_io_sink_valid),
		.io_sink_bits_id(_read_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_read_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_read_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_read_arbiter_io_sink_bits_region),
		.io_select_ready(1'h1),
		.io_select_valid(),
		.io_select_bits()
	);
	elasticDemux_3 read_demux(
		.io_source_ready(_read_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_0),
		.io_source_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_source_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_source_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_source_bits_last(_m_axi__sinkBuffer_io_deq_bits_last),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_sinks_0_valid(_read_demux_io_sinks_0_valid),
		.io_sinks_0_bits_id(_read_demux_io_sinks_0_bits_id),
		.io_sinks_0_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_sinks_0_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_sinks_0_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_sinks_1_valid(_read_demux_io_sinks_1_valid),
		.io_sinks_1_bits_id(_read_demux_io_sinks_1_bits_id),
		.io_sinks_1_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_sinks_1_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_sinks_1_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_select_ready(_read_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_io_deq_bits_id[1])
	);
	Queue32_UInt1 write_portQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueue_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_select_valid),
		.io_enq_bits(_write_arbiter_io_select_bits),
		.io_deq_ready(_write_mux_io_select_ready),
		.io_deq_valid(_write_portQueue_io_deq_valid),
		.io_deq_bits(_write_portQueue_io_deq_bits)
	);
	elasticArbiter write_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_write_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_sources_0_bits_id({1'h0, _s_axi__buffered_sourceBuffer_1_io_deq_bits_id}),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region),
		.io_sources_1_ready(_write_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_sources_1_bits_id({1'h1, _s_axi__buffered_sourceBuffer_4_io_deq_bits_id}),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_sink_valid(_write_arbiter_io_sink_valid),
		.io_sink_bits_id(_write_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_write_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_write_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_write_arbiter_io_sink_bits_region),
		.io_select_ready(_write_portQueue_io_enq_ready),
		.io_select_valid(_write_arbiter_io_select_valid),
		.io_select_bits(_write_arbiter_io_select_bits)
	);
	elasticMux_2 write_mux(
		.io_sources_0_ready(_write_mux_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_sources_0_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_sources_0_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_sources_0_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last),
		.io_sources_1_ready(_write_mux_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_sources_1_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_sources_1_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_sources_1_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last),
		.io_sink_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_sink_valid(_write_mux_io_sink_valid),
		.io_sink_bits_data(_write_mux_io_sink_bits_data),
		.io_sink_bits_strb(_write_mux_io_sink_bits_strb),
		.io_sink_bits_last(_write_mux_io_sink_bits_last),
		.io_select_ready(_write_mux_io_select_ready),
		.io_select_valid(_write_portQueue_io_deq_valid),
		.io_select_bits(_write_portQueue_io_deq_bits)
	);
	elasticDemux_4 write_demux(
		.io_source_ready(_write_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_0),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_sinks_0_valid(_write_demux_io_sinks_0_valid),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_sinks_1_valid(_write_demux_io_sinks_1_valid),
		.io_select_ready(_write_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_1_io_deq_bits_id[1])
	);
endmodule
module Counter (
	clock,
	reset,
	io_incEn,
	io_decEn,
	io_empty,
	io_full
);
	input clock;
	input reset;
	input io_incEn;
	input io_decEn;
	output wire io_empty;
	output wire io_full;
	reg [1:0] rCounter;
	always @(posedge clock)
		if (reset)
			rCounter <= 2'h0;
		else if (~(io_incEn & io_decEn)) begin
			if (io_incEn)
				rCounter <= rCounter + 2'h1;
			else if (io_decEn)
				rCounter <= rCounter - 2'h1;
		end
	assign io_empty = rCounter == 2'h0;
	assign io_full = &rCounter;
endmodule
module ram_2x93 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [92:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [92:0] W0_data;
	reg [92:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 93'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteAddressChannel_1 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [92:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_deq == do_enq))
				maybe_full <= do_enq;
		end
	ram_2x93 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({16'h0000, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[63:0];
	assign io_deq_bits_len = _ram_ext_R0_data[71:64];
	assign io_deq_bits_size = _ram_ext_R0_data[74:72];
	assign io_deq_bits_burst = _ram_ext_R0_data[76:75];
	assign io_deq_bits_lock = _ram_ext_R0_data[77];
	assign io_deq_bits_cache = _ram_ext_R0_data[81:78];
	assign io_deq_bits_prot = _ram_ext_R0_data[84:82];
	assign io_deq_bits_qos = _ram_ext_R0_data[88:85];
	assign io_deq_bits_region = _ram_ext_R0_data[92:89];
endmodule
module Queue2_ReadAddressChannel_1 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [92:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x93 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({18'h00001, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[63:0];
	assign io_deq_bits_len = _ram_ext_R0_data[71:64];
	assign io_deq_bits_size = _ram_ext_R0_data[74:72];
	assign io_deq_bits_burst = _ram_ext_R0_data[76:75];
	assign io_deq_bits_lock = _ram_ext_R0_data[77];
	assign io_deq_bits_cache = _ram_ext_R0_data[81:78];
	assign io_deq_bits_prot = _ram_ext_R0_data[84:82];
	assign io_deq_bits_qos = _ram_ext_R0_data[88:85];
	assign io_deq_bits_region = _ram_ext_R0_data[92:89];
endmodule
module AxiWriteBuffer (
	clock,
	reset,
	s_axi_ar_ready,
	s_axi_ar_valid,
	s_axi_ar_bits_addr,
	s_axi_ar_bits_len,
	s_axi_r_ready,
	s_axi_r_valid,
	s_axi_r_bits_data,
	s_axi_aw_ready,
	s_axi_aw_valid,
	s_axi_aw_bits_addr,
	s_axi_aw_bits_len,
	s_axi_w_ready,
	s_axi_w_valid,
	s_axi_w_bits_data,
	s_axi_w_bits_last,
	s_axi_b_valid,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_data,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_last,
	m_axi_b_valid
);
	input clock;
	input reset;
	output wire s_axi_ar_ready;
	input s_axi_ar_valid;
	input [63:0] s_axi_ar_bits_addr;
	input [7:0] s_axi_ar_bits_len;
	input s_axi_r_ready;
	output wire s_axi_r_valid;
	output wire [127:0] s_axi_r_bits_data;
	output wire s_axi_aw_ready;
	input s_axi_aw_valid;
	input [63:0] s_axi_aw_bits_addr;
	input [7:0] s_axi_aw_bits_len;
	output wire s_axi_w_ready;
	input s_axi_w_valid;
	input [127:0] s_axi_w_bits_data;
	input s_axi_w_bits_last;
	output wire s_axi_b_valid;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [127:0] m_axi_r_bits_data;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [127:0] m_axi_w_bits_data;
	output wire m_axi_w_bits_last;
	input m_axi_b_valid;
	wire s_axi_aw_ready_0;
	wire _sinkBuffered__sinkBuffer_1_io_enq_ready;
	wire _sinkBuffered__sinkBuffer_io_enq_ready;
	wire _counter_io_empty;
	wire _counter_io_full;
	wire _counter_io_incEn_T = s_axi_aw_ready_0 & s_axi_aw_valid;
	assign s_axi_aw_ready_0 = (_sinkBuffered__sinkBuffer_io_enq_ready & s_axi_aw_valid) & ~_counter_io_full;
	wire s_axi_ar_ready_0 = ((_sinkBuffered__sinkBuffer_1_io_enq_ready & s_axi_ar_valid) & _counter_io_empty) & ~_counter_io_incEn_T;
	Counter counter(
		.clock(clock),
		.reset(reset),
		.io_incEn(_counter_io_incEn_T),
		.io_decEn(m_axi_b_valid),
		.io_empty(_counter_io_empty),
		.io_full(_counter_io_full)
	);
	Queue2_WriteAddressChannel_1 sinkBuffered__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_io_enq_ready),
		.io_enq_valid(s_axi_aw_ready_0),
		.io_enq_bits_addr(s_axi_aw_bits_addr),
		.io_enq_bits_len(s_axi_aw_bits_len),
		.io_enq_bits_size(3'h4),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_ReadAddressChannel_1 sinkBuffered__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(s_axi_ar_ready_0),
		.io_enq_bits_addr(s_axi_ar_bits_addr),
		.io_enq_bits_len(s_axi_ar_bits_len),
		.io_enq_bits_size(3'h4),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	assign s_axi_ar_ready = s_axi_ar_ready_0;
	assign s_axi_r_valid = m_axi_r_valid;
	assign s_axi_r_bits_data = m_axi_r_bits_data;
	assign s_axi_aw_ready = s_axi_aw_ready_0;
	assign s_axi_w_ready = m_axi_w_ready;
	assign s_axi_b_valid = m_axi_b_valid;
	assign m_axi_r_ready = s_axi_r_ready;
	assign m_axi_w_valid = s_axi_w_valid;
	assign m_axi_w_bits_data = s_axi_w_bits_data;
	assign m_axi_w_bits_last = s_axi_w_bits_last;
endmodule
module AxisDataWidthConverter (
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [127:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [127:0] io_dataOut_TDATA;
	assign io_dataIn_TREADY = io_dataOut_TREADY;
	assign io_dataOut_TVALID = io_dataIn_TVALID;
	assign io_dataOut_TDATA = io_dataIn_TDATA;
endmodule
module Scheduler (
	clock,
	reset,
	io_export_taskOut_0_TREADY,
	io_export_taskOut_0_TVALID,
	io_export_taskOut_0_TDATA,
	io_export_taskOut_1_TREADY,
	io_export_taskOut_1_TVALID,
	io_export_taskOut_1_TDATA,
	io_export_taskOut_2_TREADY,
	io_export_taskOut_2_TVALID,
	io_export_taskOut_2_TDATA,
	io_export_taskOut_3_TREADY,
	io_export_taskOut_3_TVALID,
	io_export_taskOut_3_TDATA,
	io_export_taskOut_4_TREADY,
	io_export_taskOut_4_TVALID,
	io_export_taskOut_4_TDATA,
	io_export_taskOut_5_TREADY,
	io_export_taskOut_5_TVALID,
	io_export_taskOut_5_TDATA,
	io_export_taskOut_6_TREADY,
	io_export_taskOut_6_TVALID,
	io_export_taskOut_6_TDATA,
	io_export_taskOut_7_TREADY,
	io_export_taskOut_7_TVALID,
	io_export_taskOut_7_TDATA,
	io_export_taskOut_8_TREADY,
	io_export_taskOut_8_TVALID,
	io_export_taskOut_8_TDATA,
	io_export_taskOut_9_TREADY,
	io_export_taskOut_9_TVALID,
	io_export_taskOut_9_TDATA,
	io_export_taskOut_10_TREADY,
	io_export_taskOut_10_TVALID,
	io_export_taskOut_10_TDATA,
	io_export_taskOut_11_TREADY,
	io_export_taskOut_11_TVALID,
	io_export_taskOut_11_TDATA,
	io_export_taskOut_12_TREADY,
	io_export_taskOut_12_TVALID,
	io_export_taskOut_12_TDATA,
	io_export_taskOut_13_TREADY,
	io_export_taskOut_13_TVALID,
	io_export_taskOut_13_TDATA,
	io_export_taskOut_14_TREADY,
	io_export_taskOut_14_TVALID,
	io_export_taskOut_14_TDATA,
	io_export_taskOut_15_TREADY,
	io_export_taskOut_15_TVALID,
	io_export_taskOut_15_TDATA,
	io_export_taskOut_16_TREADY,
	io_export_taskOut_16_TVALID,
	io_export_taskOut_16_TDATA,
	io_export_taskOut_17_TREADY,
	io_export_taskOut_17_TVALID,
	io_export_taskOut_17_TDATA,
	io_export_taskOut_18_TREADY,
	io_export_taskOut_18_TVALID,
	io_export_taskOut_18_TDATA,
	io_export_taskOut_19_TREADY,
	io_export_taskOut_19_TVALID,
	io_export_taskOut_19_TDATA,
	io_export_taskOut_20_TREADY,
	io_export_taskOut_20_TVALID,
	io_export_taskOut_20_TDATA,
	io_export_taskOut_21_TREADY,
	io_export_taskOut_21_TVALID,
	io_export_taskOut_21_TDATA,
	io_export_taskOut_22_TREADY,
	io_export_taskOut_22_TVALID,
	io_export_taskOut_22_TDATA,
	io_export_taskOut_23_TREADY,
	io_export_taskOut_23_TVALID,
	io_export_taskOut_23_TDATA,
	io_export_taskOut_24_TREADY,
	io_export_taskOut_24_TVALID,
	io_export_taskOut_24_TDATA,
	io_export_taskOut_25_TREADY,
	io_export_taskOut_25_TVALID,
	io_export_taskOut_25_TDATA,
	io_export_taskOut_26_TREADY,
	io_export_taskOut_26_TVALID,
	io_export_taskOut_26_TDATA,
	io_export_taskOut_27_TREADY,
	io_export_taskOut_27_TVALID,
	io_export_taskOut_27_TDATA,
	io_export_taskOut_28_TREADY,
	io_export_taskOut_28_TVALID,
	io_export_taskOut_28_TDATA,
	io_export_taskOut_29_TREADY,
	io_export_taskOut_29_TVALID,
	io_export_taskOut_29_TDATA,
	io_export_taskOut_30_TREADY,
	io_export_taskOut_30_TVALID,
	io_export_taskOut_30_TDATA,
	io_export_taskOut_31_TREADY,
	io_export_taskOut_31_TVALID,
	io_export_taskOut_31_TDATA,
	io_export_taskOut_32_TREADY,
	io_export_taskOut_32_TVALID,
	io_export_taskOut_32_TDATA,
	io_export_taskOut_33_TREADY,
	io_export_taskOut_33_TVALID,
	io_export_taskOut_33_TDATA,
	io_export_taskOut_34_TREADY,
	io_export_taskOut_34_TVALID,
	io_export_taskOut_34_TDATA,
	io_export_taskOut_35_TREADY,
	io_export_taskOut_35_TVALID,
	io_export_taskOut_35_TDATA,
	io_export_taskOut_36_TREADY,
	io_export_taskOut_36_TVALID,
	io_export_taskOut_36_TDATA,
	io_export_taskOut_37_TREADY,
	io_export_taskOut_37_TVALID,
	io_export_taskOut_37_TDATA,
	io_export_taskOut_38_TREADY,
	io_export_taskOut_38_TVALID,
	io_export_taskOut_38_TDATA,
	io_export_taskOut_39_TREADY,
	io_export_taskOut_39_TVALID,
	io_export_taskOut_39_TDATA,
	io_export_taskOut_40_TREADY,
	io_export_taskOut_40_TVALID,
	io_export_taskOut_40_TDATA,
	io_export_taskOut_41_TREADY,
	io_export_taskOut_41_TVALID,
	io_export_taskOut_41_TDATA,
	io_export_taskOut_42_TREADY,
	io_export_taskOut_42_TVALID,
	io_export_taskOut_42_TDATA,
	io_export_taskOut_43_TREADY,
	io_export_taskOut_43_TVALID,
	io_export_taskOut_43_TDATA,
	io_export_taskOut_44_TREADY,
	io_export_taskOut_44_TVALID,
	io_export_taskOut_44_TDATA,
	io_export_taskOut_45_TREADY,
	io_export_taskOut_45_TVALID,
	io_export_taskOut_45_TDATA,
	io_export_taskOut_46_TREADY,
	io_export_taskOut_46_TVALID,
	io_export_taskOut_46_TDATA,
	io_export_taskOut_47_TREADY,
	io_export_taskOut_47_TVALID,
	io_export_taskOut_47_TDATA,
	io_export_taskOut_48_TREADY,
	io_export_taskOut_48_TVALID,
	io_export_taskOut_48_TDATA,
	io_export_taskOut_49_TREADY,
	io_export_taskOut_49_TVALID,
	io_export_taskOut_49_TDATA,
	io_export_taskOut_50_TREADY,
	io_export_taskOut_50_TVALID,
	io_export_taskOut_50_TDATA,
	io_export_taskOut_51_TREADY,
	io_export_taskOut_51_TVALID,
	io_export_taskOut_51_TDATA,
	io_export_taskOut_52_TREADY,
	io_export_taskOut_52_TVALID,
	io_export_taskOut_52_TDATA,
	io_export_taskOut_53_TREADY,
	io_export_taskOut_53_TVALID,
	io_export_taskOut_53_TDATA,
	io_export_taskOut_54_TREADY,
	io_export_taskOut_54_TVALID,
	io_export_taskOut_54_TDATA,
	io_export_taskOut_55_TREADY,
	io_export_taskOut_55_TVALID,
	io_export_taskOut_55_TDATA,
	io_export_taskOut_56_TREADY,
	io_export_taskOut_56_TVALID,
	io_export_taskOut_56_TDATA,
	io_export_taskOut_57_TREADY,
	io_export_taskOut_57_TVALID,
	io_export_taskOut_57_TDATA,
	io_export_taskOut_58_TREADY,
	io_export_taskOut_58_TVALID,
	io_export_taskOut_58_TDATA,
	io_export_taskOut_59_TREADY,
	io_export_taskOut_59_TVALID,
	io_export_taskOut_59_TDATA,
	io_export_taskOut_60_TREADY,
	io_export_taskOut_60_TVALID,
	io_export_taskOut_60_TDATA,
	io_export_taskOut_61_TREADY,
	io_export_taskOut_61_TVALID,
	io_export_taskOut_61_TDATA,
	io_export_taskOut_62_TREADY,
	io_export_taskOut_62_TVALID,
	io_export_taskOut_62_TDATA,
	io_export_taskOut_63_TREADY,
	io_export_taskOut_63_TVALID,
	io_export_taskOut_63_TDATA,
	io_export_taskIn_0_TREADY,
	io_export_taskIn_0_TVALID,
	io_export_taskIn_0_TDATA,
	io_export_taskIn_1_TREADY,
	io_export_taskIn_1_TVALID,
	io_export_taskIn_1_TDATA,
	io_export_taskIn_2_TREADY,
	io_export_taskIn_2_TVALID,
	io_export_taskIn_2_TDATA,
	io_export_taskIn_3_TREADY,
	io_export_taskIn_3_TVALID,
	io_export_taskIn_3_TDATA,
	io_export_taskIn_4_TREADY,
	io_export_taskIn_4_TVALID,
	io_export_taskIn_4_TDATA,
	io_export_taskIn_5_TREADY,
	io_export_taskIn_5_TVALID,
	io_export_taskIn_5_TDATA,
	io_export_taskIn_6_TREADY,
	io_export_taskIn_6_TVALID,
	io_export_taskIn_6_TDATA,
	io_export_taskIn_7_TREADY,
	io_export_taskIn_7_TVALID,
	io_export_taskIn_7_TDATA,
	io_export_taskIn_8_TREADY,
	io_export_taskIn_8_TVALID,
	io_export_taskIn_8_TDATA,
	io_export_taskIn_9_TREADY,
	io_export_taskIn_9_TVALID,
	io_export_taskIn_9_TDATA,
	io_export_taskIn_10_TREADY,
	io_export_taskIn_10_TVALID,
	io_export_taskIn_10_TDATA,
	io_export_taskIn_11_TREADY,
	io_export_taskIn_11_TVALID,
	io_export_taskIn_11_TDATA,
	io_export_taskIn_12_TREADY,
	io_export_taskIn_12_TVALID,
	io_export_taskIn_12_TDATA,
	io_export_taskIn_13_TREADY,
	io_export_taskIn_13_TVALID,
	io_export_taskIn_13_TDATA,
	io_export_taskIn_14_TREADY,
	io_export_taskIn_14_TVALID,
	io_export_taskIn_14_TDATA,
	io_export_taskIn_15_TREADY,
	io_export_taskIn_15_TVALID,
	io_export_taskIn_15_TDATA,
	io_export_taskIn_16_TREADY,
	io_export_taskIn_16_TVALID,
	io_export_taskIn_16_TDATA,
	io_export_taskIn_17_TREADY,
	io_export_taskIn_17_TVALID,
	io_export_taskIn_17_TDATA,
	io_export_taskIn_18_TREADY,
	io_export_taskIn_18_TVALID,
	io_export_taskIn_18_TDATA,
	io_export_taskIn_19_TREADY,
	io_export_taskIn_19_TVALID,
	io_export_taskIn_19_TDATA,
	io_export_taskIn_20_TREADY,
	io_export_taskIn_20_TVALID,
	io_export_taskIn_20_TDATA,
	io_export_taskIn_21_TREADY,
	io_export_taskIn_21_TVALID,
	io_export_taskIn_21_TDATA,
	io_export_taskIn_22_TREADY,
	io_export_taskIn_22_TVALID,
	io_export_taskIn_22_TDATA,
	io_export_taskIn_23_TREADY,
	io_export_taskIn_23_TVALID,
	io_export_taskIn_23_TDATA,
	io_export_taskIn_24_TREADY,
	io_export_taskIn_24_TVALID,
	io_export_taskIn_24_TDATA,
	io_export_taskIn_25_TREADY,
	io_export_taskIn_25_TVALID,
	io_export_taskIn_25_TDATA,
	io_export_taskIn_26_TREADY,
	io_export_taskIn_26_TVALID,
	io_export_taskIn_26_TDATA,
	io_export_taskIn_27_TREADY,
	io_export_taskIn_27_TVALID,
	io_export_taskIn_27_TDATA,
	io_export_taskIn_28_TREADY,
	io_export_taskIn_28_TVALID,
	io_export_taskIn_28_TDATA,
	io_export_taskIn_29_TREADY,
	io_export_taskIn_29_TVALID,
	io_export_taskIn_29_TDATA,
	io_export_taskIn_30_TREADY,
	io_export_taskIn_30_TVALID,
	io_export_taskIn_30_TDATA,
	io_export_taskIn_31_TREADY,
	io_export_taskIn_31_TVALID,
	io_export_taskIn_31_TDATA,
	io_export_taskIn_32_TREADY,
	io_export_taskIn_32_TVALID,
	io_export_taskIn_32_TDATA,
	io_export_taskIn_33_TREADY,
	io_export_taskIn_33_TVALID,
	io_export_taskIn_33_TDATA,
	io_export_taskIn_34_TREADY,
	io_export_taskIn_34_TVALID,
	io_export_taskIn_34_TDATA,
	io_export_taskIn_35_TREADY,
	io_export_taskIn_35_TVALID,
	io_export_taskIn_35_TDATA,
	io_export_taskIn_36_TREADY,
	io_export_taskIn_36_TVALID,
	io_export_taskIn_36_TDATA,
	io_export_taskIn_37_TREADY,
	io_export_taskIn_37_TVALID,
	io_export_taskIn_37_TDATA,
	io_export_taskIn_38_TREADY,
	io_export_taskIn_38_TVALID,
	io_export_taskIn_38_TDATA,
	io_export_taskIn_39_TREADY,
	io_export_taskIn_39_TVALID,
	io_export_taskIn_39_TDATA,
	io_export_taskIn_40_TREADY,
	io_export_taskIn_40_TVALID,
	io_export_taskIn_40_TDATA,
	io_export_taskIn_41_TREADY,
	io_export_taskIn_41_TVALID,
	io_export_taskIn_41_TDATA,
	io_export_taskIn_42_TREADY,
	io_export_taskIn_42_TVALID,
	io_export_taskIn_42_TDATA,
	io_export_taskIn_43_TREADY,
	io_export_taskIn_43_TVALID,
	io_export_taskIn_43_TDATA,
	io_export_taskIn_44_TREADY,
	io_export_taskIn_44_TVALID,
	io_export_taskIn_44_TDATA,
	io_export_taskIn_45_TREADY,
	io_export_taskIn_45_TVALID,
	io_export_taskIn_45_TDATA,
	io_export_taskIn_46_TREADY,
	io_export_taskIn_46_TVALID,
	io_export_taskIn_46_TDATA,
	io_export_taskIn_47_TREADY,
	io_export_taskIn_47_TVALID,
	io_export_taskIn_47_TDATA,
	io_export_taskIn_48_TREADY,
	io_export_taskIn_48_TVALID,
	io_export_taskIn_48_TDATA,
	io_export_taskIn_49_TREADY,
	io_export_taskIn_49_TVALID,
	io_export_taskIn_49_TDATA,
	io_export_taskIn_50_TREADY,
	io_export_taskIn_50_TVALID,
	io_export_taskIn_50_TDATA,
	io_export_taskIn_51_TREADY,
	io_export_taskIn_51_TVALID,
	io_export_taskIn_51_TDATA,
	io_export_taskIn_52_TREADY,
	io_export_taskIn_52_TVALID,
	io_export_taskIn_52_TDATA,
	io_export_taskIn_53_TREADY,
	io_export_taskIn_53_TVALID,
	io_export_taskIn_53_TDATA,
	io_export_taskIn_54_TREADY,
	io_export_taskIn_54_TVALID,
	io_export_taskIn_54_TDATA,
	io_export_taskIn_55_TREADY,
	io_export_taskIn_55_TVALID,
	io_export_taskIn_55_TDATA,
	io_export_taskIn_56_TREADY,
	io_export_taskIn_56_TVALID,
	io_export_taskIn_56_TDATA,
	io_export_taskIn_57_TREADY,
	io_export_taskIn_57_TVALID,
	io_export_taskIn_57_TDATA,
	io_export_taskIn_58_TREADY,
	io_export_taskIn_58_TVALID,
	io_export_taskIn_58_TDATA,
	io_export_taskIn_59_TREADY,
	io_export_taskIn_59_TVALID,
	io_export_taskIn_59_TDATA,
	io_export_taskIn_60_TREADY,
	io_export_taskIn_60_TVALID,
	io_export_taskIn_60_TDATA,
	io_export_taskIn_61_TREADY,
	io_export_taskIn_61_TVALID,
	io_export_taskIn_61_TDATA,
	io_export_taskIn_62_TREADY,
	io_export_taskIn_62_TVALID,
	io_export_taskIn_62_TDATA,
	io_export_taskIn_63_TREADY,
	io_export_taskIn_63_TVALID,
	io_export_taskIn_63_TDATA,
	io_internal_vss_axi_full_0_ar_ready,
	io_internal_vss_axi_full_0_ar_valid,
	io_internal_vss_axi_full_0_ar_bits_id,
	io_internal_vss_axi_full_0_ar_bits_addr,
	io_internal_vss_axi_full_0_ar_bits_len,
	io_internal_vss_axi_full_0_ar_bits_size,
	io_internal_vss_axi_full_0_ar_bits_burst,
	io_internal_vss_axi_full_0_ar_bits_lock,
	io_internal_vss_axi_full_0_ar_bits_cache,
	io_internal_vss_axi_full_0_ar_bits_prot,
	io_internal_vss_axi_full_0_ar_bits_qos,
	io_internal_vss_axi_full_0_ar_bits_region,
	io_internal_vss_axi_full_0_r_ready,
	io_internal_vss_axi_full_0_r_valid,
	io_internal_vss_axi_full_0_r_bits_id,
	io_internal_vss_axi_full_0_r_bits_data,
	io_internal_vss_axi_full_0_r_bits_resp,
	io_internal_vss_axi_full_0_r_bits_last,
	io_internal_vss_axi_full_0_aw_ready,
	io_internal_vss_axi_full_0_aw_valid,
	io_internal_vss_axi_full_0_aw_bits_id,
	io_internal_vss_axi_full_0_aw_bits_addr,
	io_internal_vss_axi_full_0_aw_bits_len,
	io_internal_vss_axi_full_0_aw_bits_size,
	io_internal_vss_axi_full_0_aw_bits_burst,
	io_internal_vss_axi_full_0_aw_bits_lock,
	io_internal_vss_axi_full_0_aw_bits_cache,
	io_internal_vss_axi_full_0_aw_bits_prot,
	io_internal_vss_axi_full_0_aw_bits_qos,
	io_internal_vss_axi_full_0_aw_bits_region,
	io_internal_vss_axi_full_0_w_ready,
	io_internal_vss_axi_full_0_w_valid,
	io_internal_vss_axi_full_0_w_bits_data,
	io_internal_vss_axi_full_0_w_bits_strb,
	io_internal_vss_axi_full_0_w_bits_last,
	io_internal_vss_axi_full_0_b_ready,
	io_internal_vss_axi_full_0_b_valid,
	io_internal_vss_axi_full_0_b_bits_id,
	io_internal_vss_axi_full_0_b_bits_resp,
	io_internal_axi_mgmt_vss_0_ar_ready,
	io_internal_axi_mgmt_vss_0_ar_valid,
	io_internal_axi_mgmt_vss_0_ar_bits_addr,
	io_internal_axi_mgmt_vss_0_ar_bits_prot,
	io_internal_axi_mgmt_vss_0_r_ready,
	io_internal_axi_mgmt_vss_0_r_valid,
	io_internal_axi_mgmt_vss_0_r_bits_data,
	io_internal_axi_mgmt_vss_0_r_bits_resp,
	io_internal_axi_mgmt_vss_0_aw_ready,
	io_internal_axi_mgmt_vss_0_aw_valid,
	io_internal_axi_mgmt_vss_0_aw_bits_addr,
	io_internal_axi_mgmt_vss_0_aw_bits_prot,
	io_internal_axi_mgmt_vss_0_w_ready,
	io_internal_axi_mgmt_vss_0_w_valid,
	io_internal_axi_mgmt_vss_0_w_bits_data,
	io_internal_axi_mgmt_vss_0_w_bits_strb,
	io_internal_axi_mgmt_vss_0_b_ready,
	io_internal_axi_mgmt_vss_0_b_valid,
	io_internal_axi_mgmt_vss_0_b_bits_resp,
	io_internal_axi_mgmt_vss_1_ar_ready,
	io_internal_axi_mgmt_vss_1_ar_valid,
	io_internal_axi_mgmt_vss_1_ar_bits_addr,
	io_internal_axi_mgmt_vss_1_ar_bits_prot,
	io_internal_axi_mgmt_vss_1_r_ready,
	io_internal_axi_mgmt_vss_1_r_valid,
	io_internal_axi_mgmt_vss_1_r_bits_data,
	io_internal_axi_mgmt_vss_1_r_bits_resp,
	io_internal_axi_mgmt_vss_1_aw_ready,
	io_internal_axi_mgmt_vss_1_aw_valid,
	io_internal_axi_mgmt_vss_1_aw_bits_addr,
	io_internal_axi_mgmt_vss_1_aw_bits_prot,
	io_internal_axi_mgmt_vss_1_w_ready,
	io_internal_axi_mgmt_vss_1_w_valid,
	io_internal_axi_mgmt_vss_1_w_bits_data,
	io_internal_axi_mgmt_vss_1_w_bits_strb,
	io_internal_axi_mgmt_vss_1_b_ready,
	io_internal_axi_mgmt_vss_1_b_valid,
	io_internal_axi_mgmt_vss_1_b_bits_resp
);
	input clock;
	input reset;
	input io_export_taskOut_0_TREADY;
	output wire io_export_taskOut_0_TVALID;
	output wire [127:0] io_export_taskOut_0_TDATA;
	input io_export_taskOut_1_TREADY;
	output wire io_export_taskOut_1_TVALID;
	output wire [127:0] io_export_taskOut_1_TDATA;
	input io_export_taskOut_2_TREADY;
	output wire io_export_taskOut_2_TVALID;
	output wire [127:0] io_export_taskOut_2_TDATA;
	input io_export_taskOut_3_TREADY;
	output wire io_export_taskOut_3_TVALID;
	output wire [127:0] io_export_taskOut_3_TDATA;
	input io_export_taskOut_4_TREADY;
	output wire io_export_taskOut_4_TVALID;
	output wire [127:0] io_export_taskOut_4_TDATA;
	input io_export_taskOut_5_TREADY;
	output wire io_export_taskOut_5_TVALID;
	output wire [127:0] io_export_taskOut_5_TDATA;
	input io_export_taskOut_6_TREADY;
	output wire io_export_taskOut_6_TVALID;
	output wire [127:0] io_export_taskOut_6_TDATA;
	input io_export_taskOut_7_TREADY;
	output wire io_export_taskOut_7_TVALID;
	output wire [127:0] io_export_taskOut_7_TDATA;
	input io_export_taskOut_8_TREADY;
	output wire io_export_taskOut_8_TVALID;
	output wire [127:0] io_export_taskOut_8_TDATA;
	input io_export_taskOut_9_TREADY;
	output wire io_export_taskOut_9_TVALID;
	output wire [127:0] io_export_taskOut_9_TDATA;
	input io_export_taskOut_10_TREADY;
	output wire io_export_taskOut_10_TVALID;
	output wire [127:0] io_export_taskOut_10_TDATA;
	input io_export_taskOut_11_TREADY;
	output wire io_export_taskOut_11_TVALID;
	output wire [127:0] io_export_taskOut_11_TDATA;
	input io_export_taskOut_12_TREADY;
	output wire io_export_taskOut_12_TVALID;
	output wire [127:0] io_export_taskOut_12_TDATA;
	input io_export_taskOut_13_TREADY;
	output wire io_export_taskOut_13_TVALID;
	output wire [127:0] io_export_taskOut_13_TDATA;
	input io_export_taskOut_14_TREADY;
	output wire io_export_taskOut_14_TVALID;
	output wire [127:0] io_export_taskOut_14_TDATA;
	input io_export_taskOut_15_TREADY;
	output wire io_export_taskOut_15_TVALID;
	output wire [127:0] io_export_taskOut_15_TDATA;
	input io_export_taskOut_16_TREADY;
	output wire io_export_taskOut_16_TVALID;
	output wire [127:0] io_export_taskOut_16_TDATA;
	input io_export_taskOut_17_TREADY;
	output wire io_export_taskOut_17_TVALID;
	output wire [127:0] io_export_taskOut_17_TDATA;
	input io_export_taskOut_18_TREADY;
	output wire io_export_taskOut_18_TVALID;
	output wire [127:0] io_export_taskOut_18_TDATA;
	input io_export_taskOut_19_TREADY;
	output wire io_export_taskOut_19_TVALID;
	output wire [127:0] io_export_taskOut_19_TDATA;
	input io_export_taskOut_20_TREADY;
	output wire io_export_taskOut_20_TVALID;
	output wire [127:0] io_export_taskOut_20_TDATA;
	input io_export_taskOut_21_TREADY;
	output wire io_export_taskOut_21_TVALID;
	output wire [127:0] io_export_taskOut_21_TDATA;
	input io_export_taskOut_22_TREADY;
	output wire io_export_taskOut_22_TVALID;
	output wire [127:0] io_export_taskOut_22_TDATA;
	input io_export_taskOut_23_TREADY;
	output wire io_export_taskOut_23_TVALID;
	output wire [127:0] io_export_taskOut_23_TDATA;
	input io_export_taskOut_24_TREADY;
	output wire io_export_taskOut_24_TVALID;
	output wire [127:0] io_export_taskOut_24_TDATA;
	input io_export_taskOut_25_TREADY;
	output wire io_export_taskOut_25_TVALID;
	output wire [127:0] io_export_taskOut_25_TDATA;
	input io_export_taskOut_26_TREADY;
	output wire io_export_taskOut_26_TVALID;
	output wire [127:0] io_export_taskOut_26_TDATA;
	input io_export_taskOut_27_TREADY;
	output wire io_export_taskOut_27_TVALID;
	output wire [127:0] io_export_taskOut_27_TDATA;
	input io_export_taskOut_28_TREADY;
	output wire io_export_taskOut_28_TVALID;
	output wire [127:0] io_export_taskOut_28_TDATA;
	input io_export_taskOut_29_TREADY;
	output wire io_export_taskOut_29_TVALID;
	output wire [127:0] io_export_taskOut_29_TDATA;
	input io_export_taskOut_30_TREADY;
	output wire io_export_taskOut_30_TVALID;
	output wire [127:0] io_export_taskOut_30_TDATA;
	input io_export_taskOut_31_TREADY;
	output wire io_export_taskOut_31_TVALID;
	output wire [127:0] io_export_taskOut_31_TDATA;
	input io_export_taskOut_32_TREADY;
	output wire io_export_taskOut_32_TVALID;
	output wire [127:0] io_export_taskOut_32_TDATA;
	input io_export_taskOut_33_TREADY;
	output wire io_export_taskOut_33_TVALID;
	output wire [127:0] io_export_taskOut_33_TDATA;
	input io_export_taskOut_34_TREADY;
	output wire io_export_taskOut_34_TVALID;
	output wire [127:0] io_export_taskOut_34_TDATA;
	input io_export_taskOut_35_TREADY;
	output wire io_export_taskOut_35_TVALID;
	output wire [127:0] io_export_taskOut_35_TDATA;
	input io_export_taskOut_36_TREADY;
	output wire io_export_taskOut_36_TVALID;
	output wire [127:0] io_export_taskOut_36_TDATA;
	input io_export_taskOut_37_TREADY;
	output wire io_export_taskOut_37_TVALID;
	output wire [127:0] io_export_taskOut_37_TDATA;
	input io_export_taskOut_38_TREADY;
	output wire io_export_taskOut_38_TVALID;
	output wire [127:0] io_export_taskOut_38_TDATA;
	input io_export_taskOut_39_TREADY;
	output wire io_export_taskOut_39_TVALID;
	output wire [127:0] io_export_taskOut_39_TDATA;
	input io_export_taskOut_40_TREADY;
	output wire io_export_taskOut_40_TVALID;
	output wire [127:0] io_export_taskOut_40_TDATA;
	input io_export_taskOut_41_TREADY;
	output wire io_export_taskOut_41_TVALID;
	output wire [127:0] io_export_taskOut_41_TDATA;
	input io_export_taskOut_42_TREADY;
	output wire io_export_taskOut_42_TVALID;
	output wire [127:0] io_export_taskOut_42_TDATA;
	input io_export_taskOut_43_TREADY;
	output wire io_export_taskOut_43_TVALID;
	output wire [127:0] io_export_taskOut_43_TDATA;
	input io_export_taskOut_44_TREADY;
	output wire io_export_taskOut_44_TVALID;
	output wire [127:0] io_export_taskOut_44_TDATA;
	input io_export_taskOut_45_TREADY;
	output wire io_export_taskOut_45_TVALID;
	output wire [127:0] io_export_taskOut_45_TDATA;
	input io_export_taskOut_46_TREADY;
	output wire io_export_taskOut_46_TVALID;
	output wire [127:0] io_export_taskOut_46_TDATA;
	input io_export_taskOut_47_TREADY;
	output wire io_export_taskOut_47_TVALID;
	output wire [127:0] io_export_taskOut_47_TDATA;
	input io_export_taskOut_48_TREADY;
	output wire io_export_taskOut_48_TVALID;
	output wire [127:0] io_export_taskOut_48_TDATA;
	input io_export_taskOut_49_TREADY;
	output wire io_export_taskOut_49_TVALID;
	output wire [127:0] io_export_taskOut_49_TDATA;
	input io_export_taskOut_50_TREADY;
	output wire io_export_taskOut_50_TVALID;
	output wire [127:0] io_export_taskOut_50_TDATA;
	input io_export_taskOut_51_TREADY;
	output wire io_export_taskOut_51_TVALID;
	output wire [127:0] io_export_taskOut_51_TDATA;
	input io_export_taskOut_52_TREADY;
	output wire io_export_taskOut_52_TVALID;
	output wire [127:0] io_export_taskOut_52_TDATA;
	input io_export_taskOut_53_TREADY;
	output wire io_export_taskOut_53_TVALID;
	output wire [127:0] io_export_taskOut_53_TDATA;
	input io_export_taskOut_54_TREADY;
	output wire io_export_taskOut_54_TVALID;
	output wire [127:0] io_export_taskOut_54_TDATA;
	input io_export_taskOut_55_TREADY;
	output wire io_export_taskOut_55_TVALID;
	output wire [127:0] io_export_taskOut_55_TDATA;
	input io_export_taskOut_56_TREADY;
	output wire io_export_taskOut_56_TVALID;
	output wire [127:0] io_export_taskOut_56_TDATA;
	input io_export_taskOut_57_TREADY;
	output wire io_export_taskOut_57_TVALID;
	output wire [127:0] io_export_taskOut_57_TDATA;
	input io_export_taskOut_58_TREADY;
	output wire io_export_taskOut_58_TVALID;
	output wire [127:0] io_export_taskOut_58_TDATA;
	input io_export_taskOut_59_TREADY;
	output wire io_export_taskOut_59_TVALID;
	output wire [127:0] io_export_taskOut_59_TDATA;
	input io_export_taskOut_60_TREADY;
	output wire io_export_taskOut_60_TVALID;
	output wire [127:0] io_export_taskOut_60_TDATA;
	input io_export_taskOut_61_TREADY;
	output wire io_export_taskOut_61_TVALID;
	output wire [127:0] io_export_taskOut_61_TDATA;
	input io_export_taskOut_62_TREADY;
	output wire io_export_taskOut_62_TVALID;
	output wire [127:0] io_export_taskOut_62_TDATA;
	input io_export_taskOut_63_TREADY;
	output wire io_export_taskOut_63_TVALID;
	output wire [127:0] io_export_taskOut_63_TDATA;
	output wire io_export_taskIn_0_TREADY;
	input io_export_taskIn_0_TVALID;
	input [127:0] io_export_taskIn_0_TDATA;
	output wire io_export_taskIn_1_TREADY;
	input io_export_taskIn_1_TVALID;
	input [127:0] io_export_taskIn_1_TDATA;
	output wire io_export_taskIn_2_TREADY;
	input io_export_taskIn_2_TVALID;
	input [127:0] io_export_taskIn_2_TDATA;
	output wire io_export_taskIn_3_TREADY;
	input io_export_taskIn_3_TVALID;
	input [127:0] io_export_taskIn_3_TDATA;
	output wire io_export_taskIn_4_TREADY;
	input io_export_taskIn_4_TVALID;
	input [127:0] io_export_taskIn_4_TDATA;
	output wire io_export_taskIn_5_TREADY;
	input io_export_taskIn_5_TVALID;
	input [127:0] io_export_taskIn_5_TDATA;
	output wire io_export_taskIn_6_TREADY;
	input io_export_taskIn_6_TVALID;
	input [127:0] io_export_taskIn_6_TDATA;
	output wire io_export_taskIn_7_TREADY;
	input io_export_taskIn_7_TVALID;
	input [127:0] io_export_taskIn_7_TDATA;
	output wire io_export_taskIn_8_TREADY;
	input io_export_taskIn_8_TVALID;
	input [127:0] io_export_taskIn_8_TDATA;
	output wire io_export_taskIn_9_TREADY;
	input io_export_taskIn_9_TVALID;
	input [127:0] io_export_taskIn_9_TDATA;
	output wire io_export_taskIn_10_TREADY;
	input io_export_taskIn_10_TVALID;
	input [127:0] io_export_taskIn_10_TDATA;
	output wire io_export_taskIn_11_TREADY;
	input io_export_taskIn_11_TVALID;
	input [127:0] io_export_taskIn_11_TDATA;
	output wire io_export_taskIn_12_TREADY;
	input io_export_taskIn_12_TVALID;
	input [127:0] io_export_taskIn_12_TDATA;
	output wire io_export_taskIn_13_TREADY;
	input io_export_taskIn_13_TVALID;
	input [127:0] io_export_taskIn_13_TDATA;
	output wire io_export_taskIn_14_TREADY;
	input io_export_taskIn_14_TVALID;
	input [127:0] io_export_taskIn_14_TDATA;
	output wire io_export_taskIn_15_TREADY;
	input io_export_taskIn_15_TVALID;
	input [127:0] io_export_taskIn_15_TDATA;
	output wire io_export_taskIn_16_TREADY;
	input io_export_taskIn_16_TVALID;
	input [127:0] io_export_taskIn_16_TDATA;
	output wire io_export_taskIn_17_TREADY;
	input io_export_taskIn_17_TVALID;
	input [127:0] io_export_taskIn_17_TDATA;
	output wire io_export_taskIn_18_TREADY;
	input io_export_taskIn_18_TVALID;
	input [127:0] io_export_taskIn_18_TDATA;
	output wire io_export_taskIn_19_TREADY;
	input io_export_taskIn_19_TVALID;
	input [127:0] io_export_taskIn_19_TDATA;
	output wire io_export_taskIn_20_TREADY;
	input io_export_taskIn_20_TVALID;
	input [127:0] io_export_taskIn_20_TDATA;
	output wire io_export_taskIn_21_TREADY;
	input io_export_taskIn_21_TVALID;
	input [127:0] io_export_taskIn_21_TDATA;
	output wire io_export_taskIn_22_TREADY;
	input io_export_taskIn_22_TVALID;
	input [127:0] io_export_taskIn_22_TDATA;
	output wire io_export_taskIn_23_TREADY;
	input io_export_taskIn_23_TVALID;
	input [127:0] io_export_taskIn_23_TDATA;
	output wire io_export_taskIn_24_TREADY;
	input io_export_taskIn_24_TVALID;
	input [127:0] io_export_taskIn_24_TDATA;
	output wire io_export_taskIn_25_TREADY;
	input io_export_taskIn_25_TVALID;
	input [127:0] io_export_taskIn_25_TDATA;
	output wire io_export_taskIn_26_TREADY;
	input io_export_taskIn_26_TVALID;
	input [127:0] io_export_taskIn_26_TDATA;
	output wire io_export_taskIn_27_TREADY;
	input io_export_taskIn_27_TVALID;
	input [127:0] io_export_taskIn_27_TDATA;
	output wire io_export_taskIn_28_TREADY;
	input io_export_taskIn_28_TVALID;
	input [127:0] io_export_taskIn_28_TDATA;
	output wire io_export_taskIn_29_TREADY;
	input io_export_taskIn_29_TVALID;
	input [127:0] io_export_taskIn_29_TDATA;
	output wire io_export_taskIn_30_TREADY;
	input io_export_taskIn_30_TVALID;
	input [127:0] io_export_taskIn_30_TDATA;
	output wire io_export_taskIn_31_TREADY;
	input io_export_taskIn_31_TVALID;
	input [127:0] io_export_taskIn_31_TDATA;
	output wire io_export_taskIn_32_TREADY;
	input io_export_taskIn_32_TVALID;
	input [127:0] io_export_taskIn_32_TDATA;
	output wire io_export_taskIn_33_TREADY;
	input io_export_taskIn_33_TVALID;
	input [127:0] io_export_taskIn_33_TDATA;
	output wire io_export_taskIn_34_TREADY;
	input io_export_taskIn_34_TVALID;
	input [127:0] io_export_taskIn_34_TDATA;
	output wire io_export_taskIn_35_TREADY;
	input io_export_taskIn_35_TVALID;
	input [127:0] io_export_taskIn_35_TDATA;
	output wire io_export_taskIn_36_TREADY;
	input io_export_taskIn_36_TVALID;
	input [127:0] io_export_taskIn_36_TDATA;
	output wire io_export_taskIn_37_TREADY;
	input io_export_taskIn_37_TVALID;
	input [127:0] io_export_taskIn_37_TDATA;
	output wire io_export_taskIn_38_TREADY;
	input io_export_taskIn_38_TVALID;
	input [127:0] io_export_taskIn_38_TDATA;
	output wire io_export_taskIn_39_TREADY;
	input io_export_taskIn_39_TVALID;
	input [127:0] io_export_taskIn_39_TDATA;
	output wire io_export_taskIn_40_TREADY;
	input io_export_taskIn_40_TVALID;
	input [127:0] io_export_taskIn_40_TDATA;
	output wire io_export_taskIn_41_TREADY;
	input io_export_taskIn_41_TVALID;
	input [127:0] io_export_taskIn_41_TDATA;
	output wire io_export_taskIn_42_TREADY;
	input io_export_taskIn_42_TVALID;
	input [127:0] io_export_taskIn_42_TDATA;
	output wire io_export_taskIn_43_TREADY;
	input io_export_taskIn_43_TVALID;
	input [127:0] io_export_taskIn_43_TDATA;
	output wire io_export_taskIn_44_TREADY;
	input io_export_taskIn_44_TVALID;
	input [127:0] io_export_taskIn_44_TDATA;
	output wire io_export_taskIn_45_TREADY;
	input io_export_taskIn_45_TVALID;
	input [127:0] io_export_taskIn_45_TDATA;
	output wire io_export_taskIn_46_TREADY;
	input io_export_taskIn_46_TVALID;
	input [127:0] io_export_taskIn_46_TDATA;
	output wire io_export_taskIn_47_TREADY;
	input io_export_taskIn_47_TVALID;
	input [127:0] io_export_taskIn_47_TDATA;
	output wire io_export_taskIn_48_TREADY;
	input io_export_taskIn_48_TVALID;
	input [127:0] io_export_taskIn_48_TDATA;
	output wire io_export_taskIn_49_TREADY;
	input io_export_taskIn_49_TVALID;
	input [127:0] io_export_taskIn_49_TDATA;
	output wire io_export_taskIn_50_TREADY;
	input io_export_taskIn_50_TVALID;
	input [127:0] io_export_taskIn_50_TDATA;
	output wire io_export_taskIn_51_TREADY;
	input io_export_taskIn_51_TVALID;
	input [127:0] io_export_taskIn_51_TDATA;
	output wire io_export_taskIn_52_TREADY;
	input io_export_taskIn_52_TVALID;
	input [127:0] io_export_taskIn_52_TDATA;
	output wire io_export_taskIn_53_TREADY;
	input io_export_taskIn_53_TVALID;
	input [127:0] io_export_taskIn_53_TDATA;
	output wire io_export_taskIn_54_TREADY;
	input io_export_taskIn_54_TVALID;
	input [127:0] io_export_taskIn_54_TDATA;
	output wire io_export_taskIn_55_TREADY;
	input io_export_taskIn_55_TVALID;
	input [127:0] io_export_taskIn_55_TDATA;
	output wire io_export_taskIn_56_TREADY;
	input io_export_taskIn_56_TVALID;
	input [127:0] io_export_taskIn_56_TDATA;
	output wire io_export_taskIn_57_TREADY;
	input io_export_taskIn_57_TVALID;
	input [127:0] io_export_taskIn_57_TDATA;
	output wire io_export_taskIn_58_TREADY;
	input io_export_taskIn_58_TVALID;
	input [127:0] io_export_taskIn_58_TDATA;
	output wire io_export_taskIn_59_TREADY;
	input io_export_taskIn_59_TVALID;
	input [127:0] io_export_taskIn_59_TDATA;
	output wire io_export_taskIn_60_TREADY;
	input io_export_taskIn_60_TVALID;
	input [127:0] io_export_taskIn_60_TDATA;
	output wire io_export_taskIn_61_TREADY;
	input io_export_taskIn_61_TVALID;
	input [127:0] io_export_taskIn_61_TDATA;
	output wire io_export_taskIn_62_TREADY;
	input io_export_taskIn_62_TVALID;
	input [127:0] io_export_taskIn_62_TDATA;
	output wire io_export_taskIn_63_TREADY;
	input io_export_taskIn_63_TVALID;
	input [127:0] io_export_taskIn_63_TDATA;
	input io_internal_vss_axi_full_0_ar_ready;
	output wire io_internal_vss_axi_full_0_ar_valid;
	output wire [1:0] io_internal_vss_axi_full_0_ar_bits_id;
	output wire [63:0] io_internal_vss_axi_full_0_ar_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_ar_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_ar_bits_burst;
	output wire io_internal_vss_axi_full_0_ar_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_region;
	output wire io_internal_vss_axi_full_0_r_ready;
	input io_internal_vss_axi_full_0_r_valid;
	input [1:0] io_internal_vss_axi_full_0_r_bits_id;
	input [127:0] io_internal_vss_axi_full_0_r_bits_data;
	input [1:0] io_internal_vss_axi_full_0_r_bits_resp;
	input io_internal_vss_axi_full_0_r_bits_last;
	input io_internal_vss_axi_full_0_aw_ready;
	output wire io_internal_vss_axi_full_0_aw_valid;
	output wire [1:0] io_internal_vss_axi_full_0_aw_bits_id;
	output wire [63:0] io_internal_vss_axi_full_0_aw_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_aw_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_aw_bits_burst;
	output wire io_internal_vss_axi_full_0_aw_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_region;
	input io_internal_vss_axi_full_0_w_ready;
	output wire io_internal_vss_axi_full_0_w_valid;
	output wire [127:0] io_internal_vss_axi_full_0_w_bits_data;
	output wire [15:0] io_internal_vss_axi_full_0_w_bits_strb;
	output wire io_internal_vss_axi_full_0_w_bits_last;
	output wire io_internal_vss_axi_full_0_b_ready;
	input io_internal_vss_axi_full_0_b_valid;
	input [1:0] io_internal_vss_axi_full_0_b_bits_id;
	input [1:0] io_internal_vss_axi_full_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vss_0_ar_ready;
	input io_internal_axi_mgmt_vss_0_ar_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_ar_bits_prot;
	input io_internal_axi_mgmt_vss_0_r_ready;
	output wire io_internal_axi_mgmt_vss_0_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vss_0_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vss_0_r_bits_resp;
	output wire io_internal_axi_mgmt_vss_0_aw_ready;
	input io_internal_axi_mgmt_vss_0_aw_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_aw_bits_prot;
	output wire io_internal_axi_mgmt_vss_0_w_ready;
	input io_internal_axi_mgmt_vss_0_w_valid;
	input [63:0] io_internal_axi_mgmt_vss_0_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vss_0_w_bits_strb;
	input io_internal_axi_mgmt_vss_0_b_ready;
	output wire io_internal_axi_mgmt_vss_0_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vss_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vss_1_ar_ready;
	input io_internal_axi_mgmt_vss_1_ar_valid;
	input [5:0] io_internal_axi_mgmt_vss_1_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_1_ar_bits_prot;
	input io_internal_axi_mgmt_vss_1_r_ready;
	output wire io_internal_axi_mgmt_vss_1_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vss_1_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vss_1_r_bits_resp;
	output wire io_internal_axi_mgmt_vss_1_aw_ready;
	input io_internal_axi_mgmt_vss_1_aw_valid;
	input [5:0] io_internal_axi_mgmt_vss_1_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_1_aw_bits_prot;
	output wire io_internal_axi_mgmt_vss_1_w_ready;
	input io_internal_axi_mgmt_vss_1_w_valid;
	input [63:0] io_internal_axi_mgmt_vss_1_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vss_1_w_bits_strb;
	input io_internal_axi_mgmt_vss_1_b_ready;
	output wire io_internal_axi_mgmt_vss_1_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vss_1_b_bits_resp;
	wire _axis_stream_converters_in_63_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_63_io_dataOut_TDATA;
	wire _axis_stream_converters_in_62_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_62_io_dataOut_TDATA;
	wire _axis_stream_converters_in_61_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_61_io_dataOut_TDATA;
	wire _axis_stream_converters_in_60_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_60_io_dataOut_TDATA;
	wire _axis_stream_converters_in_59_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_59_io_dataOut_TDATA;
	wire _axis_stream_converters_in_58_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_58_io_dataOut_TDATA;
	wire _axis_stream_converters_in_57_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_57_io_dataOut_TDATA;
	wire _axis_stream_converters_in_56_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_56_io_dataOut_TDATA;
	wire _axis_stream_converters_in_55_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_55_io_dataOut_TDATA;
	wire _axis_stream_converters_in_54_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_54_io_dataOut_TDATA;
	wire _axis_stream_converters_in_53_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_53_io_dataOut_TDATA;
	wire _axis_stream_converters_in_52_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_52_io_dataOut_TDATA;
	wire _axis_stream_converters_in_51_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_51_io_dataOut_TDATA;
	wire _axis_stream_converters_in_50_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_50_io_dataOut_TDATA;
	wire _axis_stream_converters_in_49_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_49_io_dataOut_TDATA;
	wire _axis_stream_converters_in_48_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_48_io_dataOut_TDATA;
	wire _axis_stream_converters_in_47_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_47_io_dataOut_TDATA;
	wire _axis_stream_converters_in_46_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_46_io_dataOut_TDATA;
	wire _axis_stream_converters_in_45_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_45_io_dataOut_TDATA;
	wire _axis_stream_converters_in_44_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_44_io_dataOut_TDATA;
	wire _axis_stream_converters_in_43_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_43_io_dataOut_TDATA;
	wire _axis_stream_converters_in_42_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_42_io_dataOut_TDATA;
	wire _axis_stream_converters_in_41_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_41_io_dataOut_TDATA;
	wire _axis_stream_converters_in_40_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_40_io_dataOut_TDATA;
	wire _axis_stream_converters_in_39_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_39_io_dataOut_TDATA;
	wire _axis_stream_converters_in_38_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_38_io_dataOut_TDATA;
	wire _axis_stream_converters_in_37_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_37_io_dataOut_TDATA;
	wire _axis_stream_converters_in_36_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_36_io_dataOut_TDATA;
	wire _axis_stream_converters_in_35_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_35_io_dataOut_TDATA;
	wire _axis_stream_converters_in_34_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_34_io_dataOut_TDATA;
	wire _axis_stream_converters_in_33_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_33_io_dataOut_TDATA;
	wire _axis_stream_converters_in_32_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_32_io_dataOut_TDATA;
	wire _axis_stream_converters_in_31_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_31_io_dataOut_TDATA;
	wire _axis_stream_converters_in_30_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_30_io_dataOut_TDATA;
	wire _axis_stream_converters_in_29_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_29_io_dataOut_TDATA;
	wire _axis_stream_converters_in_28_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_28_io_dataOut_TDATA;
	wire _axis_stream_converters_in_27_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_27_io_dataOut_TDATA;
	wire _axis_stream_converters_in_26_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_26_io_dataOut_TDATA;
	wire _axis_stream_converters_in_25_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_25_io_dataOut_TDATA;
	wire _axis_stream_converters_in_24_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_24_io_dataOut_TDATA;
	wire _axis_stream_converters_in_23_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_23_io_dataOut_TDATA;
	wire _axis_stream_converters_in_22_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_22_io_dataOut_TDATA;
	wire _axis_stream_converters_in_21_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_21_io_dataOut_TDATA;
	wire _axis_stream_converters_in_20_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_20_io_dataOut_TDATA;
	wire _axis_stream_converters_in_19_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_19_io_dataOut_TDATA;
	wire _axis_stream_converters_in_18_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_18_io_dataOut_TDATA;
	wire _axis_stream_converters_in_17_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_17_io_dataOut_TDATA;
	wire _axis_stream_converters_in_16_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_16_io_dataOut_TDATA;
	wire _axis_stream_converters_in_15_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_15_io_dataOut_TDATA;
	wire _axis_stream_converters_in_14_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_14_io_dataOut_TDATA;
	wire _axis_stream_converters_in_13_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_13_io_dataOut_TDATA;
	wire _axis_stream_converters_in_12_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_12_io_dataOut_TDATA;
	wire _axis_stream_converters_in_11_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_11_io_dataOut_TDATA;
	wire _axis_stream_converters_in_10_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_10_io_dataOut_TDATA;
	wire _axis_stream_converters_in_9_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_9_io_dataOut_TDATA;
	wire _axis_stream_converters_in_8_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_8_io_dataOut_TDATA;
	wire _axis_stream_converters_in_7_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_7_io_dataOut_TDATA;
	wire _axis_stream_converters_in_6_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_6_io_dataOut_TDATA;
	wire _axis_stream_converters_in_5_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_5_io_dataOut_TDATA;
	wire _axis_stream_converters_in_4_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_4_io_dataOut_TDATA;
	wire _axis_stream_converters_in_3_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_3_io_dataOut_TDATA;
	wire _axis_stream_converters_in_2_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_2_io_dataOut_TDATA;
	wire _axis_stream_converters_in_1_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_1_io_dataOut_TDATA;
	wire _axis_stream_converters_in_0_io_dataOut_TVALID;
	wire [127:0] _axis_stream_converters_in_0_io_dataOut_TDATA;
	wire _axis_stream_converters_out_63_io_dataIn_TREADY;
	wire _axis_stream_converters_out_62_io_dataIn_TREADY;
	wire _axis_stream_converters_out_61_io_dataIn_TREADY;
	wire _axis_stream_converters_out_60_io_dataIn_TREADY;
	wire _axis_stream_converters_out_59_io_dataIn_TREADY;
	wire _axis_stream_converters_out_58_io_dataIn_TREADY;
	wire _axis_stream_converters_out_57_io_dataIn_TREADY;
	wire _axis_stream_converters_out_56_io_dataIn_TREADY;
	wire _axis_stream_converters_out_55_io_dataIn_TREADY;
	wire _axis_stream_converters_out_54_io_dataIn_TREADY;
	wire _axis_stream_converters_out_53_io_dataIn_TREADY;
	wire _axis_stream_converters_out_52_io_dataIn_TREADY;
	wire _axis_stream_converters_out_51_io_dataIn_TREADY;
	wire _axis_stream_converters_out_50_io_dataIn_TREADY;
	wire _axis_stream_converters_out_49_io_dataIn_TREADY;
	wire _axis_stream_converters_out_48_io_dataIn_TREADY;
	wire _axis_stream_converters_out_47_io_dataIn_TREADY;
	wire _axis_stream_converters_out_46_io_dataIn_TREADY;
	wire _axis_stream_converters_out_45_io_dataIn_TREADY;
	wire _axis_stream_converters_out_44_io_dataIn_TREADY;
	wire _axis_stream_converters_out_43_io_dataIn_TREADY;
	wire _axis_stream_converters_out_42_io_dataIn_TREADY;
	wire _axis_stream_converters_out_41_io_dataIn_TREADY;
	wire _axis_stream_converters_out_40_io_dataIn_TREADY;
	wire _axis_stream_converters_out_39_io_dataIn_TREADY;
	wire _axis_stream_converters_out_38_io_dataIn_TREADY;
	wire _axis_stream_converters_out_37_io_dataIn_TREADY;
	wire _axis_stream_converters_out_36_io_dataIn_TREADY;
	wire _axis_stream_converters_out_35_io_dataIn_TREADY;
	wire _axis_stream_converters_out_34_io_dataIn_TREADY;
	wire _axis_stream_converters_out_33_io_dataIn_TREADY;
	wire _axis_stream_converters_out_32_io_dataIn_TREADY;
	wire _axis_stream_converters_out_31_io_dataIn_TREADY;
	wire _axis_stream_converters_out_30_io_dataIn_TREADY;
	wire _axis_stream_converters_out_29_io_dataIn_TREADY;
	wire _axis_stream_converters_out_28_io_dataIn_TREADY;
	wire _axis_stream_converters_out_27_io_dataIn_TREADY;
	wire _axis_stream_converters_out_26_io_dataIn_TREADY;
	wire _axis_stream_converters_out_25_io_dataIn_TREADY;
	wire _axis_stream_converters_out_24_io_dataIn_TREADY;
	wire _axis_stream_converters_out_23_io_dataIn_TREADY;
	wire _axis_stream_converters_out_22_io_dataIn_TREADY;
	wire _axis_stream_converters_out_21_io_dataIn_TREADY;
	wire _axis_stream_converters_out_20_io_dataIn_TREADY;
	wire _axis_stream_converters_out_19_io_dataIn_TREADY;
	wire _axis_stream_converters_out_18_io_dataIn_TREADY;
	wire _axis_stream_converters_out_17_io_dataIn_TREADY;
	wire _axis_stream_converters_out_16_io_dataIn_TREADY;
	wire _axis_stream_converters_out_15_io_dataIn_TREADY;
	wire _axis_stream_converters_out_14_io_dataIn_TREADY;
	wire _axis_stream_converters_out_13_io_dataIn_TREADY;
	wire _axis_stream_converters_out_12_io_dataIn_TREADY;
	wire _axis_stream_converters_out_11_io_dataIn_TREADY;
	wire _axis_stream_converters_out_10_io_dataIn_TREADY;
	wire _axis_stream_converters_out_9_io_dataIn_TREADY;
	wire _axis_stream_converters_out_8_io_dataIn_TREADY;
	wire _axis_stream_converters_out_7_io_dataIn_TREADY;
	wire _axis_stream_converters_out_6_io_dataIn_TREADY;
	wire _axis_stream_converters_out_5_io_dataIn_TREADY;
	wire _axis_stream_converters_out_4_io_dataIn_TREADY;
	wire _axis_stream_converters_out_3_io_dataIn_TREADY;
	wire _axis_stream_converters_out_2_io_dataIn_TREADY;
	wire _axis_stream_converters_out_1_io_dataIn_TREADY;
	wire _axis_stream_converters_out_0_io_dataIn_TREADY;
	wire _module_1_s_axi_ar_ready;
	wire _module_1_s_axi_r_valid;
	wire [127:0] _module_1_s_axi_r_bits_data;
	wire _module_1_s_axi_aw_ready;
	wire _module_1_s_axi_w_ready;
	wire _module_1_s_axi_b_valid;
	wire _module_1_m_axi_ar_valid;
	wire [63:0] _module_1_m_axi_ar_bits_addr;
	wire [7:0] _module_1_m_axi_ar_bits_len;
	wire [2:0] _module_1_m_axi_ar_bits_size;
	wire [1:0] _module_1_m_axi_ar_bits_burst;
	wire _module_1_m_axi_ar_bits_lock;
	wire [3:0] _module_1_m_axi_ar_bits_cache;
	wire [2:0] _module_1_m_axi_ar_bits_prot;
	wire [3:0] _module_1_m_axi_ar_bits_qos;
	wire [3:0] _module_1_m_axi_ar_bits_region;
	wire _module_1_m_axi_r_ready;
	wire _module_1_m_axi_aw_valid;
	wire [63:0] _module_1_m_axi_aw_bits_addr;
	wire [7:0] _module_1_m_axi_aw_bits_len;
	wire [2:0] _module_1_m_axi_aw_bits_size;
	wire [1:0] _module_1_m_axi_aw_bits_burst;
	wire _module_1_m_axi_aw_bits_lock;
	wire [3:0] _module_1_m_axi_aw_bits_cache;
	wire [2:0] _module_1_m_axi_aw_bits_prot;
	wire [3:0] _module_1_m_axi_aw_bits_qos;
	wire [3:0] _module_1_m_axi_aw_bits_region;
	wire _module_1_m_axi_w_valid;
	wire [127:0] _module_1_m_axi_w_bits_data;
	wire _module_1_m_axi_w_bits_last;
	wire _module_s_axi_ar_ready;
	wire _module_s_axi_r_valid;
	wire [127:0] _module_s_axi_r_bits_data;
	wire _module_s_axi_aw_ready;
	wire _module_s_axi_w_ready;
	wire _module_s_axi_b_valid;
	wire _module_m_axi_ar_valid;
	wire [63:0] _module_m_axi_ar_bits_addr;
	wire [7:0] _module_m_axi_ar_bits_len;
	wire [2:0] _module_m_axi_ar_bits_size;
	wire [1:0] _module_m_axi_ar_bits_burst;
	wire _module_m_axi_ar_bits_lock;
	wire [3:0] _module_m_axi_ar_bits_cache;
	wire [2:0] _module_m_axi_ar_bits_prot;
	wire [3:0] _module_m_axi_ar_bits_qos;
	wire [3:0] _module_m_axi_ar_bits_region;
	wire _module_m_axi_r_ready;
	wire _module_m_axi_aw_valid;
	wire [63:0] _module_m_axi_aw_bits_addr;
	wire [7:0] _module_m_axi_aw_bits_len;
	wire [2:0] _module_m_axi_aw_bits_size;
	wire [1:0] _module_m_axi_aw_bits_burst;
	wire _module_m_axi_aw_bits_lock;
	wire [3:0] _module_m_axi_aw_bits_cache;
	wire [2:0] _module_m_axi_aw_bits_prot;
	wire [3:0] _module_m_axi_aw_bits_qos;
	wire [3:0] _module_m_axi_aw_bits_region;
	wire _module_m_axi_w_valid;
	wire [127:0] _module_m_axi_w_bits_data;
	wire _module_m_axi_w_bits_last;
	wire _mux_s_axi_0_ar_ready;
	wire _mux_s_axi_0_r_valid;
	wire [127:0] _mux_s_axi_0_r_bits_data;
	wire _mux_s_axi_0_aw_ready;
	wire _mux_s_axi_0_w_ready;
	wire _mux_s_axi_0_b_valid;
	wire _mux_s_axi_1_ar_ready;
	wire _mux_s_axi_1_r_valid;
	wire [127:0] _mux_s_axi_1_r_bits_data;
	wire _mux_s_axi_1_aw_ready;
	wire _mux_s_axi_1_w_ready;
	wire _mux_s_axi_1_b_valid;
	wire _vssRvm_1_io_read_address_ready;
	wire _vssRvm_1_io_read_data_valid;
	wire [127:0] _vssRvm_1_io_read_data_bits;
	wire _vssRvm_1_io_write_address_ready;
	wire _vssRvm_1_io_write_data_ready;
	wire _vssRvm_1_axi_ar_valid;
	wire [63:0] _vssRvm_1_axi_ar_bits_addr;
	wire [7:0] _vssRvm_1_axi_ar_bits_len;
	wire _vssRvm_1_axi_r_ready;
	wire _vssRvm_1_axi_aw_valid;
	wire [63:0] _vssRvm_1_axi_aw_bits_addr;
	wire [7:0] _vssRvm_1_axi_aw_bits_len;
	wire _vssRvm_1_axi_w_valid;
	wire [127:0] _vssRvm_1_axi_w_bits_data;
	wire _vssRvm_1_axi_w_bits_last;
	wire _vssRvm_0_io_read_address_ready;
	wire _vssRvm_0_io_read_data_valid;
	wire [127:0] _vssRvm_0_io_read_data_bits;
	wire _vssRvm_0_io_write_address_ready;
	wire _vssRvm_0_io_write_data_ready;
	wire _vssRvm_0_axi_ar_valid;
	wire [63:0] _vssRvm_0_axi_ar_bits_addr;
	wire [7:0] _vssRvm_0_axi_ar_bits_len;
	wire _vssRvm_0_axi_r_ready;
	wire _vssRvm_0_axi_aw_valid;
	wire [63:0] _vssRvm_0_axi_aw_bits_addr;
	wire [7:0] _vssRvm_0_axi_aw_bits_len;
	wire _vssRvm_0_axi_w_valid;
	wire [127:0] _vssRvm_0_axi_w_bits_data;
	wire _vssRvm_0_axi_w_bits_last;
	wire _virtualStealServers_1_io_connNetwork_ctrl_serveStealReq_valid;
	wire _virtualStealServers_1_io_connNetwork_data_availableTask_ready;
	wire _virtualStealServers_1_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _virtualStealServers_1_io_connNetwork_data_qOutTask_bits;
	wire _virtualStealServers_1_io_read_address_valid;
	wire [63:0] _virtualStealServers_1_io_read_address_bits;
	wire _virtualStealServers_1_io_read_data_ready;
	wire [3:0] _virtualStealServers_1_io_read_burst_len;
	wire _virtualStealServers_1_io_write_address_valid;
	wire [63:0] _virtualStealServers_1_io_write_address_bits;
	wire _virtualStealServers_1_io_write_data_valid;
	wire [127:0] _virtualStealServers_1_io_write_data_bits;
	wire [3:0] _virtualStealServers_1_io_write_burst_len;
	wire _virtualStealServers_1_io_write_last;
	wire _virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _virtualStealServers_0_io_connNetwork_data_availableTask_ready;
	wire _virtualStealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _virtualStealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _virtualStealServers_0_io_read_address_valid;
	wire [63:0] _virtualStealServers_0_io_read_address_bits;
	wire _virtualStealServers_0_io_read_data_ready;
	wire [3:0] _virtualStealServers_0_io_read_burst_len;
	wire _virtualStealServers_0_io_write_address_valid;
	wire [63:0] _virtualStealServers_0_io_write_address_bits;
	wire _virtualStealServers_0_io_write_data_valid;
	wire [127:0] _virtualStealServers_0_io_write_data_bits;
	wire [3:0] _virtualStealServers_0_io_write_burst_len;
	wire _virtualStealServers_0_io_write_last;
	wire _stealNW_TQ_io_connPE_0_push_ready;
	wire _stealNW_TQ_io_connPE_0_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_0_pop_bits;
	wire _stealNW_TQ_io_connPE_1_push_ready;
	wire _stealNW_TQ_io_connPE_1_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_1_pop_bits;
	wire _stealNW_TQ_io_connPE_2_push_ready;
	wire _stealNW_TQ_io_connPE_2_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_2_pop_bits;
	wire _stealNW_TQ_io_connPE_3_push_ready;
	wire _stealNW_TQ_io_connPE_3_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_3_pop_bits;
	wire _stealNW_TQ_io_connPE_4_push_ready;
	wire _stealNW_TQ_io_connPE_4_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_4_pop_bits;
	wire _stealNW_TQ_io_connPE_5_push_ready;
	wire _stealNW_TQ_io_connPE_5_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_5_pop_bits;
	wire _stealNW_TQ_io_connPE_6_push_ready;
	wire _stealNW_TQ_io_connPE_6_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_6_pop_bits;
	wire _stealNW_TQ_io_connPE_7_push_ready;
	wire _stealNW_TQ_io_connPE_7_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_7_pop_bits;
	wire _stealNW_TQ_io_connPE_8_push_ready;
	wire _stealNW_TQ_io_connPE_8_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_8_pop_bits;
	wire _stealNW_TQ_io_connPE_9_push_ready;
	wire _stealNW_TQ_io_connPE_9_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_9_pop_bits;
	wire _stealNW_TQ_io_connPE_10_push_ready;
	wire _stealNW_TQ_io_connPE_10_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_10_pop_bits;
	wire _stealNW_TQ_io_connPE_11_push_ready;
	wire _stealNW_TQ_io_connPE_11_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_11_pop_bits;
	wire _stealNW_TQ_io_connPE_12_push_ready;
	wire _stealNW_TQ_io_connPE_12_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_12_pop_bits;
	wire _stealNW_TQ_io_connPE_13_push_ready;
	wire _stealNW_TQ_io_connPE_13_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_13_pop_bits;
	wire _stealNW_TQ_io_connPE_14_push_ready;
	wire _stealNW_TQ_io_connPE_14_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_14_pop_bits;
	wire _stealNW_TQ_io_connPE_15_push_ready;
	wire _stealNW_TQ_io_connPE_15_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_15_pop_bits;
	wire _stealNW_TQ_io_connPE_16_push_ready;
	wire _stealNW_TQ_io_connPE_16_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_16_pop_bits;
	wire _stealNW_TQ_io_connPE_17_push_ready;
	wire _stealNW_TQ_io_connPE_17_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_17_pop_bits;
	wire _stealNW_TQ_io_connPE_18_push_ready;
	wire _stealNW_TQ_io_connPE_18_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_18_pop_bits;
	wire _stealNW_TQ_io_connPE_19_push_ready;
	wire _stealNW_TQ_io_connPE_19_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_19_pop_bits;
	wire _stealNW_TQ_io_connPE_20_push_ready;
	wire _stealNW_TQ_io_connPE_20_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_20_pop_bits;
	wire _stealNW_TQ_io_connPE_21_push_ready;
	wire _stealNW_TQ_io_connPE_21_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_21_pop_bits;
	wire _stealNW_TQ_io_connPE_22_push_ready;
	wire _stealNW_TQ_io_connPE_22_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_22_pop_bits;
	wire _stealNW_TQ_io_connPE_23_push_ready;
	wire _stealNW_TQ_io_connPE_23_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_23_pop_bits;
	wire _stealNW_TQ_io_connPE_24_push_ready;
	wire _stealNW_TQ_io_connPE_24_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_24_pop_bits;
	wire _stealNW_TQ_io_connPE_25_push_ready;
	wire _stealNW_TQ_io_connPE_25_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_25_pop_bits;
	wire _stealNW_TQ_io_connPE_26_push_ready;
	wire _stealNW_TQ_io_connPE_26_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_26_pop_bits;
	wire _stealNW_TQ_io_connPE_27_push_ready;
	wire _stealNW_TQ_io_connPE_27_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_27_pop_bits;
	wire _stealNW_TQ_io_connPE_28_push_ready;
	wire _stealNW_TQ_io_connPE_28_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_28_pop_bits;
	wire _stealNW_TQ_io_connPE_29_push_ready;
	wire _stealNW_TQ_io_connPE_29_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_29_pop_bits;
	wire _stealNW_TQ_io_connPE_30_push_ready;
	wire _stealNW_TQ_io_connPE_30_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_30_pop_bits;
	wire _stealNW_TQ_io_connPE_31_push_ready;
	wire _stealNW_TQ_io_connPE_31_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_31_pop_bits;
	wire _stealNW_TQ_io_connPE_32_push_ready;
	wire _stealNW_TQ_io_connPE_32_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_32_pop_bits;
	wire _stealNW_TQ_io_connPE_33_push_ready;
	wire _stealNW_TQ_io_connPE_33_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_33_pop_bits;
	wire _stealNW_TQ_io_connPE_34_push_ready;
	wire _stealNW_TQ_io_connPE_34_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_34_pop_bits;
	wire _stealNW_TQ_io_connPE_35_push_ready;
	wire _stealNW_TQ_io_connPE_35_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_35_pop_bits;
	wire _stealNW_TQ_io_connPE_36_push_ready;
	wire _stealNW_TQ_io_connPE_36_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_36_pop_bits;
	wire _stealNW_TQ_io_connPE_37_push_ready;
	wire _stealNW_TQ_io_connPE_37_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_37_pop_bits;
	wire _stealNW_TQ_io_connPE_38_push_ready;
	wire _stealNW_TQ_io_connPE_38_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_38_pop_bits;
	wire _stealNW_TQ_io_connPE_39_push_ready;
	wire _stealNW_TQ_io_connPE_39_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_39_pop_bits;
	wire _stealNW_TQ_io_connPE_40_push_ready;
	wire _stealNW_TQ_io_connPE_40_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_40_pop_bits;
	wire _stealNW_TQ_io_connPE_41_push_ready;
	wire _stealNW_TQ_io_connPE_41_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_41_pop_bits;
	wire _stealNW_TQ_io_connPE_42_push_ready;
	wire _stealNW_TQ_io_connPE_42_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_42_pop_bits;
	wire _stealNW_TQ_io_connPE_43_push_ready;
	wire _stealNW_TQ_io_connPE_43_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_43_pop_bits;
	wire _stealNW_TQ_io_connPE_44_push_ready;
	wire _stealNW_TQ_io_connPE_44_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_44_pop_bits;
	wire _stealNW_TQ_io_connPE_45_push_ready;
	wire _stealNW_TQ_io_connPE_45_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_45_pop_bits;
	wire _stealNW_TQ_io_connPE_46_push_ready;
	wire _stealNW_TQ_io_connPE_46_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_46_pop_bits;
	wire _stealNW_TQ_io_connPE_47_push_ready;
	wire _stealNW_TQ_io_connPE_47_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_47_pop_bits;
	wire _stealNW_TQ_io_connPE_48_push_ready;
	wire _stealNW_TQ_io_connPE_48_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_48_pop_bits;
	wire _stealNW_TQ_io_connPE_49_push_ready;
	wire _stealNW_TQ_io_connPE_49_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_49_pop_bits;
	wire _stealNW_TQ_io_connPE_50_push_ready;
	wire _stealNW_TQ_io_connPE_50_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_50_pop_bits;
	wire _stealNW_TQ_io_connPE_51_push_ready;
	wire _stealNW_TQ_io_connPE_51_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_51_pop_bits;
	wire _stealNW_TQ_io_connPE_52_push_ready;
	wire _stealNW_TQ_io_connPE_52_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_52_pop_bits;
	wire _stealNW_TQ_io_connPE_53_push_ready;
	wire _stealNW_TQ_io_connPE_53_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_53_pop_bits;
	wire _stealNW_TQ_io_connPE_54_push_ready;
	wire _stealNW_TQ_io_connPE_54_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_54_pop_bits;
	wire _stealNW_TQ_io_connPE_55_push_ready;
	wire _stealNW_TQ_io_connPE_55_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_55_pop_bits;
	wire _stealNW_TQ_io_connPE_56_push_ready;
	wire _stealNW_TQ_io_connPE_56_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_56_pop_bits;
	wire _stealNW_TQ_io_connPE_57_push_ready;
	wire _stealNW_TQ_io_connPE_57_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_57_pop_bits;
	wire _stealNW_TQ_io_connPE_58_push_ready;
	wire _stealNW_TQ_io_connPE_58_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_58_pop_bits;
	wire _stealNW_TQ_io_connPE_59_push_ready;
	wire _stealNW_TQ_io_connPE_59_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_59_pop_bits;
	wire _stealNW_TQ_io_connPE_60_push_ready;
	wire _stealNW_TQ_io_connPE_60_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_60_pop_bits;
	wire _stealNW_TQ_io_connPE_61_push_ready;
	wire _stealNW_TQ_io_connPE_61_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_61_pop_bits;
	wire _stealNW_TQ_io_connPE_62_push_ready;
	wire _stealNW_TQ_io_connPE_62_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_62_pop_bits;
	wire _stealNW_TQ_io_connPE_63_push_ready;
	wire _stealNW_TQ_io_connPE_63_pop_valid;
	wire [127:0] _stealNW_TQ_io_connPE_63_pop_bits;
	wire _stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready;
	wire _stealNW_TQ_io_connVSS_0_data_availableTask_valid;
	wire [127:0] _stealNW_TQ_io_connVSS_0_data_availableTask_bits;
	wire _stealNW_TQ_io_connVSS_0_data_qOutTask_ready;
	wire _stealNW_TQ_io_connVSS_1_ctrl_serveStealReq_ready;
	wire _stealNW_TQ_io_connVSS_1_data_availableTask_valid;
	wire [127:0] _stealNW_TQ_io_connVSS_1_data_availableTask_bits;
	wire _stealNW_TQ_io_connVSS_1_data_qOutTask_ready;
	wire _stealNW_TQ_io_ntwDataUnitOccupancyVSS_0;
	wire _stealNW_TQ_io_ntwDataUnitOccupancyVSS_1;
	SchedulerLocalNetwork stealNW_TQ(
		.clock(clock),
		.reset(reset),
		.io_connPE_0_push_ready(_stealNW_TQ_io_connPE_0_push_ready),
		.io_connPE_0_push_valid(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_connPE_0_push_bits(_axis_stream_converters_in_0_io_dataOut_TDATA),
		.io_connPE_0_pop_ready(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_connPE_0_pop_valid(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_connPE_0_pop_bits(_stealNW_TQ_io_connPE_0_pop_bits),
		.io_connPE_1_push_ready(_stealNW_TQ_io_connPE_1_push_ready),
		.io_connPE_1_push_valid(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_connPE_1_push_bits(_axis_stream_converters_in_1_io_dataOut_TDATA),
		.io_connPE_1_pop_ready(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_connPE_1_pop_valid(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_connPE_1_pop_bits(_stealNW_TQ_io_connPE_1_pop_bits),
		.io_connPE_2_push_ready(_stealNW_TQ_io_connPE_2_push_ready),
		.io_connPE_2_push_valid(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_connPE_2_push_bits(_axis_stream_converters_in_2_io_dataOut_TDATA),
		.io_connPE_2_pop_ready(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_connPE_2_pop_valid(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_connPE_2_pop_bits(_stealNW_TQ_io_connPE_2_pop_bits),
		.io_connPE_3_push_ready(_stealNW_TQ_io_connPE_3_push_ready),
		.io_connPE_3_push_valid(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_connPE_3_push_bits(_axis_stream_converters_in_3_io_dataOut_TDATA),
		.io_connPE_3_pop_ready(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_connPE_3_pop_valid(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_connPE_3_pop_bits(_stealNW_TQ_io_connPE_3_pop_bits),
		.io_connPE_4_push_ready(_stealNW_TQ_io_connPE_4_push_ready),
		.io_connPE_4_push_valid(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_connPE_4_push_bits(_axis_stream_converters_in_4_io_dataOut_TDATA),
		.io_connPE_4_pop_ready(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_connPE_4_pop_valid(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_connPE_4_pop_bits(_stealNW_TQ_io_connPE_4_pop_bits),
		.io_connPE_5_push_ready(_stealNW_TQ_io_connPE_5_push_ready),
		.io_connPE_5_push_valid(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_connPE_5_push_bits(_axis_stream_converters_in_5_io_dataOut_TDATA),
		.io_connPE_5_pop_ready(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_connPE_5_pop_valid(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_connPE_5_pop_bits(_stealNW_TQ_io_connPE_5_pop_bits),
		.io_connPE_6_push_ready(_stealNW_TQ_io_connPE_6_push_ready),
		.io_connPE_6_push_valid(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_connPE_6_push_bits(_axis_stream_converters_in_6_io_dataOut_TDATA),
		.io_connPE_6_pop_ready(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_connPE_6_pop_valid(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_connPE_6_pop_bits(_stealNW_TQ_io_connPE_6_pop_bits),
		.io_connPE_7_push_ready(_stealNW_TQ_io_connPE_7_push_ready),
		.io_connPE_7_push_valid(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_connPE_7_push_bits(_axis_stream_converters_in_7_io_dataOut_TDATA),
		.io_connPE_7_pop_ready(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_connPE_7_pop_valid(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_connPE_7_pop_bits(_stealNW_TQ_io_connPE_7_pop_bits),
		.io_connPE_8_push_ready(_stealNW_TQ_io_connPE_8_push_ready),
		.io_connPE_8_push_valid(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_connPE_8_push_bits(_axis_stream_converters_in_8_io_dataOut_TDATA),
		.io_connPE_8_pop_ready(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_connPE_8_pop_valid(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_connPE_8_pop_bits(_stealNW_TQ_io_connPE_8_pop_bits),
		.io_connPE_9_push_ready(_stealNW_TQ_io_connPE_9_push_ready),
		.io_connPE_9_push_valid(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_connPE_9_push_bits(_axis_stream_converters_in_9_io_dataOut_TDATA),
		.io_connPE_9_pop_ready(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_connPE_9_pop_valid(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_connPE_9_pop_bits(_stealNW_TQ_io_connPE_9_pop_bits),
		.io_connPE_10_push_ready(_stealNW_TQ_io_connPE_10_push_ready),
		.io_connPE_10_push_valid(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_connPE_10_push_bits(_axis_stream_converters_in_10_io_dataOut_TDATA),
		.io_connPE_10_pop_ready(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_connPE_10_pop_valid(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_connPE_10_pop_bits(_stealNW_TQ_io_connPE_10_pop_bits),
		.io_connPE_11_push_ready(_stealNW_TQ_io_connPE_11_push_ready),
		.io_connPE_11_push_valid(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_connPE_11_push_bits(_axis_stream_converters_in_11_io_dataOut_TDATA),
		.io_connPE_11_pop_ready(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_connPE_11_pop_valid(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_connPE_11_pop_bits(_stealNW_TQ_io_connPE_11_pop_bits),
		.io_connPE_12_push_ready(_stealNW_TQ_io_connPE_12_push_ready),
		.io_connPE_12_push_valid(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_connPE_12_push_bits(_axis_stream_converters_in_12_io_dataOut_TDATA),
		.io_connPE_12_pop_ready(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_connPE_12_pop_valid(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_connPE_12_pop_bits(_stealNW_TQ_io_connPE_12_pop_bits),
		.io_connPE_13_push_ready(_stealNW_TQ_io_connPE_13_push_ready),
		.io_connPE_13_push_valid(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_connPE_13_push_bits(_axis_stream_converters_in_13_io_dataOut_TDATA),
		.io_connPE_13_pop_ready(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_connPE_13_pop_valid(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_connPE_13_pop_bits(_stealNW_TQ_io_connPE_13_pop_bits),
		.io_connPE_14_push_ready(_stealNW_TQ_io_connPE_14_push_ready),
		.io_connPE_14_push_valid(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_connPE_14_push_bits(_axis_stream_converters_in_14_io_dataOut_TDATA),
		.io_connPE_14_pop_ready(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_connPE_14_pop_valid(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_connPE_14_pop_bits(_stealNW_TQ_io_connPE_14_pop_bits),
		.io_connPE_15_push_ready(_stealNW_TQ_io_connPE_15_push_ready),
		.io_connPE_15_push_valid(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_connPE_15_push_bits(_axis_stream_converters_in_15_io_dataOut_TDATA),
		.io_connPE_15_pop_ready(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_connPE_15_pop_valid(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_connPE_15_pop_bits(_stealNW_TQ_io_connPE_15_pop_bits),
		.io_connPE_16_push_ready(_stealNW_TQ_io_connPE_16_push_ready),
		.io_connPE_16_push_valid(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_connPE_16_push_bits(_axis_stream_converters_in_16_io_dataOut_TDATA),
		.io_connPE_16_pop_ready(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_connPE_16_pop_valid(_stealNW_TQ_io_connPE_16_pop_valid),
		.io_connPE_16_pop_bits(_stealNW_TQ_io_connPE_16_pop_bits),
		.io_connPE_17_push_ready(_stealNW_TQ_io_connPE_17_push_ready),
		.io_connPE_17_push_valid(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_connPE_17_push_bits(_axis_stream_converters_in_17_io_dataOut_TDATA),
		.io_connPE_17_pop_ready(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_connPE_17_pop_valid(_stealNW_TQ_io_connPE_17_pop_valid),
		.io_connPE_17_pop_bits(_stealNW_TQ_io_connPE_17_pop_bits),
		.io_connPE_18_push_ready(_stealNW_TQ_io_connPE_18_push_ready),
		.io_connPE_18_push_valid(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_connPE_18_push_bits(_axis_stream_converters_in_18_io_dataOut_TDATA),
		.io_connPE_18_pop_ready(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_connPE_18_pop_valid(_stealNW_TQ_io_connPE_18_pop_valid),
		.io_connPE_18_pop_bits(_stealNW_TQ_io_connPE_18_pop_bits),
		.io_connPE_19_push_ready(_stealNW_TQ_io_connPE_19_push_ready),
		.io_connPE_19_push_valid(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_connPE_19_push_bits(_axis_stream_converters_in_19_io_dataOut_TDATA),
		.io_connPE_19_pop_ready(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_connPE_19_pop_valid(_stealNW_TQ_io_connPE_19_pop_valid),
		.io_connPE_19_pop_bits(_stealNW_TQ_io_connPE_19_pop_bits),
		.io_connPE_20_push_ready(_stealNW_TQ_io_connPE_20_push_ready),
		.io_connPE_20_push_valid(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_connPE_20_push_bits(_axis_stream_converters_in_20_io_dataOut_TDATA),
		.io_connPE_20_pop_ready(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_connPE_20_pop_valid(_stealNW_TQ_io_connPE_20_pop_valid),
		.io_connPE_20_pop_bits(_stealNW_TQ_io_connPE_20_pop_bits),
		.io_connPE_21_push_ready(_stealNW_TQ_io_connPE_21_push_ready),
		.io_connPE_21_push_valid(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_connPE_21_push_bits(_axis_stream_converters_in_21_io_dataOut_TDATA),
		.io_connPE_21_pop_ready(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_connPE_21_pop_valid(_stealNW_TQ_io_connPE_21_pop_valid),
		.io_connPE_21_pop_bits(_stealNW_TQ_io_connPE_21_pop_bits),
		.io_connPE_22_push_ready(_stealNW_TQ_io_connPE_22_push_ready),
		.io_connPE_22_push_valid(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_connPE_22_push_bits(_axis_stream_converters_in_22_io_dataOut_TDATA),
		.io_connPE_22_pop_ready(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_connPE_22_pop_valid(_stealNW_TQ_io_connPE_22_pop_valid),
		.io_connPE_22_pop_bits(_stealNW_TQ_io_connPE_22_pop_bits),
		.io_connPE_23_push_ready(_stealNW_TQ_io_connPE_23_push_ready),
		.io_connPE_23_push_valid(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_connPE_23_push_bits(_axis_stream_converters_in_23_io_dataOut_TDATA),
		.io_connPE_23_pop_ready(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_connPE_23_pop_valid(_stealNW_TQ_io_connPE_23_pop_valid),
		.io_connPE_23_pop_bits(_stealNW_TQ_io_connPE_23_pop_bits),
		.io_connPE_24_push_ready(_stealNW_TQ_io_connPE_24_push_ready),
		.io_connPE_24_push_valid(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_connPE_24_push_bits(_axis_stream_converters_in_24_io_dataOut_TDATA),
		.io_connPE_24_pop_ready(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_connPE_24_pop_valid(_stealNW_TQ_io_connPE_24_pop_valid),
		.io_connPE_24_pop_bits(_stealNW_TQ_io_connPE_24_pop_bits),
		.io_connPE_25_push_ready(_stealNW_TQ_io_connPE_25_push_ready),
		.io_connPE_25_push_valid(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_connPE_25_push_bits(_axis_stream_converters_in_25_io_dataOut_TDATA),
		.io_connPE_25_pop_ready(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_connPE_25_pop_valid(_stealNW_TQ_io_connPE_25_pop_valid),
		.io_connPE_25_pop_bits(_stealNW_TQ_io_connPE_25_pop_bits),
		.io_connPE_26_push_ready(_stealNW_TQ_io_connPE_26_push_ready),
		.io_connPE_26_push_valid(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_connPE_26_push_bits(_axis_stream_converters_in_26_io_dataOut_TDATA),
		.io_connPE_26_pop_ready(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_connPE_26_pop_valid(_stealNW_TQ_io_connPE_26_pop_valid),
		.io_connPE_26_pop_bits(_stealNW_TQ_io_connPE_26_pop_bits),
		.io_connPE_27_push_ready(_stealNW_TQ_io_connPE_27_push_ready),
		.io_connPE_27_push_valid(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_connPE_27_push_bits(_axis_stream_converters_in_27_io_dataOut_TDATA),
		.io_connPE_27_pop_ready(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_connPE_27_pop_valid(_stealNW_TQ_io_connPE_27_pop_valid),
		.io_connPE_27_pop_bits(_stealNW_TQ_io_connPE_27_pop_bits),
		.io_connPE_28_push_ready(_stealNW_TQ_io_connPE_28_push_ready),
		.io_connPE_28_push_valid(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_connPE_28_push_bits(_axis_stream_converters_in_28_io_dataOut_TDATA),
		.io_connPE_28_pop_ready(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_connPE_28_pop_valid(_stealNW_TQ_io_connPE_28_pop_valid),
		.io_connPE_28_pop_bits(_stealNW_TQ_io_connPE_28_pop_bits),
		.io_connPE_29_push_ready(_stealNW_TQ_io_connPE_29_push_ready),
		.io_connPE_29_push_valid(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_connPE_29_push_bits(_axis_stream_converters_in_29_io_dataOut_TDATA),
		.io_connPE_29_pop_ready(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_connPE_29_pop_valid(_stealNW_TQ_io_connPE_29_pop_valid),
		.io_connPE_29_pop_bits(_stealNW_TQ_io_connPE_29_pop_bits),
		.io_connPE_30_push_ready(_stealNW_TQ_io_connPE_30_push_ready),
		.io_connPE_30_push_valid(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_connPE_30_push_bits(_axis_stream_converters_in_30_io_dataOut_TDATA),
		.io_connPE_30_pop_ready(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_connPE_30_pop_valid(_stealNW_TQ_io_connPE_30_pop_valid),
		.io_connPE_30_pop_bits(_stealNW_TQ_io_connPE_30_pop_bits),
		.io_connPE_31_push_ready(_stealNW_TQ_io_connPE_31_push_ready),
		.io_connPE_31_push_valid(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_connPE_31_push_bits(_axis_stream_converters_in_31_io_dataOut_TDATA),
		.io_connPE_31_pop_ready(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_connPE_31_pop_valid(_stealNW_TQ_io_connPE_31_pop_valid),
		.io_connPE_31_pop_bits(_stealNW_TQ_io_connPE_31_pop_bits),
		.io_connPE_32_push_ready(_stealNW_TQ_io_connPE_32_push_ready),
		.io_connPE_32_push_valid(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_connPE_32_push_bits(_axis_stream_converters_in_32_io_dataOut_TDATA),
		.io_connPE_32_pop_ready(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_connPE_32_pop_valid(_stealNW_TQ_io_connPE_32_pop_valid),
		.io_connPE_32_pop_bits(_stealNW_TQ_io_connPE_32_pop_bits),
		.io_connPE_33_push_ready(_stealNW_TQ_io_connPE_33_push_ready),
		.io_connPE_33_push_valid(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_connPE_33_push_bits(_axis_stream_converters_in_33_io_dataOut_TDATA),
		.io_connPE_33_pop_ready(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_connPE_33_pop_valid(_stealNW_TQ_io_connPE_33_pop_valid),
		.io_connPE_33_pop_bits(_stealNW_TQ_io_connPE_33_pop_bits),
		.io_connPE_34_push_ready(_stealNW_TQ_io_connPE_34_push_ready),
		.io_connPE_34_push_valid(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_connPE_34_push_bits(_axis_stream_converters_in_34_io_dataOut_TDATA),
		.io_connPE_34_pop_ready(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_connPE_34_pop_valid(_stealNW_TQ_io_connPE_34_pop_valid),
		.io_connPE_34_pop_bits(_stealNW_TQ_io_connPE_34_pop_bits),
		.io_connPE_35_push_ready(_stealNW_TQ_io_connPE_35_push_ready),
		.io_connPE_35_push_valid(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_connPE_35_push_bits(_axis_stream_converters_in_35_io_dataOut_TDATA),
		.io_connPE_35_pop_ready(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_connPE_35_pop_valid(_stealNW_TQ_io_connPE_35_pop_valid),
		.io_connPE_35_pop_bits(_stealNW_TQ_io_connPE_35_pop_bits),
		.io_connPE_36_push_ready(_stealNW_TQ_io_connPE_36_push_ready),
		.io_connPE_36_push_valid(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_connPE_36_push_bits(_axis_stream_converters_in_36_io_dataOut_TDATA),
		.io_connPE_36_pop_ready(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_connPE_36_pop_valid(_stealNW_TQ_io_connPE_36_pop_valid),
		.io_connPE_36_pop_bits(_stealNW_TQ_io_connPE_36_pop_bits),
		.io_connPE_37_push_ready(_stealNW_TQ_io_connPE_37_push_ready),
		.io_connPE_37_push_valid(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_connPE_37_push_bits(_axis_stream_converters_in_37_io_dataOut_TDATA),
		.io_connPE_37_pop_ready(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_connPE_37_pop_valid(_stealNW_TQ_io_connPE_37_pop_valid),
		.io_connPE_37_pop_bits(_stealNW_TQ_io_connPE_37_pop_bits),
		.io_connPE_38_push_ready(_stealNW_TQ_io_connPE_38_push_ready),
		.io_connPE_38_push_valid(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_connPE_38_push_bits(_axis_stream_converters_in_38_io_dataOut_TDATA),
		.io_connPE_38_pop_ready(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_connPE_38_pop_valid(_stealNW_TQ_io_connPE_38_pop_valid),
		.io_connPE_38_pop_bits(_stealNW_TQ_io_connPE_38_pop_bits),
		.io_connPE_39_push_ready(_stealNW_TQ_io_connPE_39_push_ready),
		.io_connPE_39_push_valid(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_connPE_39_push_bits(_axis_stream_converters_in_39_io_dataOut_TDATA),
		.io_connPE_39_pop_ready(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_connPE_39_pop_valid(_stealNW_TQ_io_connPE_39_pop_valid),
		.io_connPE_39_pop_bits(_stealNW_TQ_io_connPE_39_pop_bits),
		.io_connPE_40_push_ready(_stealNW_TQ_io_connPE_40_push_ready),
		.io_connPE_40_push_valid(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_connPE_40_push_bits(_axis_stream_converters_in_40_io_dataOut_TDATA),
		.io_connPE_40_pop_ready(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_connPE_40_pop_valid(_stealNW_TQ_io_connPE_40_pop_valid),
		.io_connPE_40_pop_bits(_stealNW_TQ_io_connPE_40_pop_bits),
		.io_connPE_41_push_ready(_stealNW_TQ_io_connPE_41_push_ready),
		.io_connPE_41_push_valid(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_connPE_41_push_bits(_axis_stream_converters_in_41_io_dataOut_TDATA),
		.io_connPE_41_pop_ready(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_connPE_41_pop_valid(_stealNW_TQ_io_connPE_41_pop_valid),
		.io_connPE_41_pop_bits(_stealNW_TQ_io_connPE_41_pop_bits),
		.io_connPE_42_push_ready(_stealNW_TQ_io_connPE_42_push_ready),
		.io_connPE_42_push_valid(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_connPE_42_push_bits(_axis_stream_converters_in_42_io_dataOut_TDATA),
		.io_connPE_42_pop_ready(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_connPE_42_pop_valid(_stealNW_TQ_io_connPE_42_pop_valid),
		.io_connPE_42_pop_bits(_stealNW_TQ_io_connPE_42_pop_bits),
		.io_connPE_43_push_ready(_stealNW_TQ_io_connPE_43_push_ready),
		.io_connPE_43_push_valid(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_connPE_43_push_bits(_axis_stream_converters_in_43_io_dataOut_TDATA),
		.io_connPE_43_pop_ready(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_connPE_43_pop_valid(_stealNW_TQ_io_connPE_43_pop_valid),
		.io_connPE_43_pop_bits(_stealNW_TQ_io_connPE_43_pop_bits),
		.io_connPE_44_push_ready(_stealNW_TQ_io_connPE_44_push_ready),
		.io_connPE_44_push_valid(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_connPE_44_push_bits(_axis_stream_converters_in_44_io_dataOut_TDATA),
		.io_connPE_44_pop_ready(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_connPE_44_pop_valid(_stealNW_TQ_io_connPE_44_pop_valid),
		.io_connPE_44_pop_bits(_stealNW_TQ_io_connPE_44_pop_bits),
		.io_connPE_45_push_ready(_stealNW_TQ_io_connPE_45_push_ready),
		.io_connPE_45_push_valid(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_connPE_45_push_bits(_axis_stream_converters_in_45_io_dataOut_TDATA),
		.io_connPE_45_pop_ready(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_connPE_45_pop_valid(_stealNW_TQ_io_connPE_45_pop_valid),
		.io_connPE_45_pop_bits(_stealNW_TQ_io_connPE_45_pop_bits),
		.io_connPE_46_push_ready(_stealNW_TQ_io_connPE_46_push_ready),
		.io_connPE_46_push_valid(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_connPE_46_push_bits(_axis_stream_converters_in_46_io_dataOut_TDATA),
		.io_connPE_46_pop_ready(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_connPE_46_pop_valid(_stealNW_TQ_io_connPE_46_pop_valid),
		.io_connPE_46_pop_bits(_stealNW_TQ_io_connPE_46_pop_bits),
		.io_connPE_47_push_ready(_stealNW_TQ_io_connPE_47_push_ready),
		.io_connPE_47_push_valid(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_connPE_47_push_bits(_axis_stream_converters_in_47_io_dataOut_TDATA),
		.io_connPE_47_pop_ready(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_connPE_47_pop_valid(_stealNW_TQ_io_connPE_47_pop_valid),
		.io_connPE_47_pop_bits(_stealNW_TQ_io_connPE_47_pop_bits),
		.io_connPE_48_push_ready(_stealNW_TQ_io_connPE_48_push_ready),
		.io_connPE_48_push_valid(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_connPE_48_push_bits(_axis_stream_converters_in_48_io_dataOut_TDATA),
		.io_connPE_48_pop_ready(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_connPE_48_pop_valid(_stealNW_TQ_io_connPE_48_pop_valid),
		.io_connPE_48_pop_bits(_stealNW_TQ_io_connPE_48_pop_bits),
		.io_connPE_49_push_ready(_stealNW_TQ_io_connPE_49_push_ready),
		.io_connPE_49_push_valid(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_connPE_49_push_bits(_axis_stream_converters_in_49_io_dataOut_TDATA),
		.io_connPE_49_pop_ready(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_connPE_49_pop_valid(_stealNW_TQ_io_connPE_49_pop_valid),
		.io_connPE_49_pop_bits(_stealNW_TQ_io_connPE_49_pop_bits),
		.io_connPE_50_push_ready(_stealNW_TQ_io_connPE_50_push_ready),
		.io_connPE_50_push_valid(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_connPE_50_push_bits(_axis_stream_converters_in_50_io_dataOut_TDATA),
		.io_connPE_50_pop_ready(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_connPE_50_pop_valid(_stealNW_TQ_io_connPE_50_pop_valid),
		.io_connPE_50_pop_bits(_stealNW_TQ_io_connPE_50_pop_bits),
		.io_connPE_51_push_ready(_stealNW_TQ_io_connPE_51_push_ready),
		.io_connPE_51_push_valid(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_connPE_51_push_bits(_axis_stream_converters_in_51_io_dataOut_TDATA),
		.io_connPE_51_pop_ready(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_connPE_51_pop_valid(_stealNW_TQ_io_connPE_51_pop_valid),
		.io_connPE_51_pop_bits(_stealNW_TQ_io_connPE_51_pop_bits),
		.io_connPE_52_push_ready(_stealNW_TQ_io_connPE_52_push_ready),
		.io_connPE_52_push_valid(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_connPE_52_push_bits(_axis_stream_converters_in_52_io_dataOut_TDATA),
		.io_connPE_52_pop_ready(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_connPE_52_pop_valid(_stealNW_TQ_io_connPE_52_pop_valid),
		.io_connPE_52_pop_bits(_stealNW_TQ_io_connPE_52_pop_bits),
		.io_connPE_53_push_ready(_stealNW_TQ_io_connPE_53_push_ready),
		.io_connPE_53_push_valid(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_connPE_53_push_bits(_axis_stream_converters_in_53_io_dataOut_TDATA),
		.io_connPE_53_pop_ready(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_connPE_53_pop_valid(_stealNW_TQ_io_connPE_53_pop_valid),
		.io_connPE_53_pop_bits(_stealNW_TQ_io_connPE_53_pop_bits),
		.io_connPE_54_push_ready(_stealNW_TQ_io_connPE_54_push_ready),
		.io_connPE_54_push_valid(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_connPE_54_push_bits(_axis_stream_converters_in_54_io_dataOut_TDATA),
		.io_connPE_54_pop_ready(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_connPE_54_pop_valid(_stealNW_TQ_io_connPE_54_pop_valid),
		.io_connPE_54_pop_bits(_stealNW_TQ_io_connPE_54_pop_bits),
		.io_connPE_55_push_ready(_stealNW_TQ_io_connPE_55_push_ready),
		.io_connPE_55_push_valid(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_connPE_55_push_bits(_axis_stream_converters_in_55_io_dataOut_TDATA),
		.io_connPE_55_pop_ready(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_connPE_55_pop_valid(_stealNW_TQ_io_connPE_55_pop_valid),
		.io_connPE_55_pop_bits(_stealNW_TQ_io_connPE_55_pop_bits),
		.io_connPE_56_push_ready(_stealNW_TQ_io_connPE_56_push_ready),
		.io_connPE_56_push_valid(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_connPE_56_push_bits(_axis_stream_converters_in_56_io_dataOut_TDATA),
		.io_connPE_56_pop_ready(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_connPE_56_pop_valid(_stealNW_TQ_io_connPE_56_pop_valid),
		.io_connPE_56_pop_bits(_stealNW_TQ_io_connPE_56_pop_bits),
		.io_connPE_57_push_ready(_stealNW_TQ_io_connPE_57_push_ready),
		.io_connPE_57_push_valid(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_connPE_57_push_bits(_axis_stream_converters_in_57_io_dataOut_TDATA),
		.io_connPE_57_pop_ready(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_connPE_57_pop_valid(_stealNW_TQ_io_connPE_57_pop_valid),
		.io_connPE_57_pop_bits(_stealNW_TQ_io_connPE_57_pop_bits),
		.io_connPE_58_push_ready(_stealNW_TQ_io_connPE_58_push_ready),
		.io_connPE_58_push_valid(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_connPE_58_push_bits(_axis_stream_converters_in_58_io_dataOut_TDATA),
		.io_connPE_58_pop_ready(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_connPE_58_pop_valid(_stealNW_TQ_io_connPE_58_pop_valid),
		.io_connPE_58_pop_bits(_stealNW_TQ_io_connPE_58_pop_bits),
		.io_connPE_59_push_ready(_stealNW_TQ_io_connPE_59_push_ready),
		.io_connPE_59_push_valid(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_connPE_59_push_bits(_axis_stream_converters_in_59_io_dataOut_TDATA),
		.io_connPE_59_pop_ready(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_connPE_59_pop_valid(_stealNW_TQ_io_connPE_59_pop_valid),
		.io_connPE_59_pop_bits(_stealNW_TQ_io_connPE_59_pop_bits),
		.io_connPE_60_push_ready(_stealNW_TQ_io_connPE_60_push_ready),
		.io_connPE_60_push_valid(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_connPE_60_push_bits(_axis_stream_converters_in_60_io_dataOut_TDATA),
		.io_connPE_60_pop_ready(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_connPE_60_pop_valid(_stealNW_TQ_io_connPE_60_pop_valid),
		.io_connPE_60_pop_bits(_stealNW_TQ_io_connPE_60_pop_bits),
		.io_connPE_61_push_ready(_stealNW_TQ_io_connPE_61_push_ready),
		.io_connPE_61_push_valid(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_connPE_61_push_bits(_axis_stream_converters_in_61_io_dataOut_TDATA),
		.io_connPE_61_pop_ready(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_connPE_61_pop_valid(_stealNW_TQ_io_connPE_61_pop_valid),
		.io_connPE_61_pop_bits(_stealNW_TQ_io_connPE_61_pop_bits),
		.io_connPE_62_push_ready(_stealNW_TQ_io_connPE_62_push_ready),
		.io_connPE_62_push_valid(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_connPE_62_push_bits(_axis_stream_converters_in_62_io_dataOut_TDATA),
		.io_connPE_62_pop_ready(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_connPE_62_pop_valid(_stealNW_TQ_io_connPE_62_pop_valid),
		.io_connPE_62_pop_bits(_stealNW_TQ_io_connPE_62_pop_bits),
		.io_connPE_63_push_ready(_stealNW_TQ_io_connPE_63_push_ready),
		.io_connPE_63_push_valid(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_connPE_63_push_bits(_axis_stream_converters_in_63_io_dataOut_TDATA),
		.io_connPE_63_pop_ready(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_connPE_63_pop_valid(_stealNW_TQ_io_connPE_63_pop_valid),
		.io_connPE_63_pop_bits(_stealNW_TQ_io_connPE_63_pop_bits),
		.io_connVSS_0_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connVSS_0_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connVSS_0_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connVSS_0_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connVSS_0_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connVSS_0_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connVSS_0_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connVSS_0_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connVSS_1_ctrl_serveStealReq_valid(_virtualStealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connVSS_1_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_1_ctrl_serveStealReq_ready),
		.io_connVSS_1_data_availableTask_ready(_virtualStealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connVSS_1_data_availableTask_valid(_stealNW_TQ_io_connVSS_1_data_availableTask_valid),
		.io_connVSS_1_data_availableTask_bits(_stealNW_TQ_io_connVSS_1_data_availableTask_bits),
		.io_connVSS_1_data_qOutTask_ready(_stealNW_TQ_io_connVSS_1_data_qOutTask_ready),
		.io_connVSS_1_data_qOutTask_valid(_virtualStealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connVSS_1_data_qOutTask_bits(_virtualStealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0),
		.io_ntwDataUnitOccupancyVSS_1(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_1)
	);
	SchedulerServer virtualStealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connNetwork_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vss_0_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vss_0_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vss_0_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vss_0_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vss_0_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vss_0_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vss_0_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vss_0_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vss_0_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vss_0_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vss_0_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vss_0_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vss_0_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vss_0_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vss_0_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vss_0_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vss_0_b_bits_resp),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_read_burst_len(_virtualStealServers_0_io_read_burst_len),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_write_burst_len(_virtualStealServers_0_io_write_burst_len),
		.io_write_last(_virtualStealServers_0_io_write_last),
		.io_ntwDataUnitOccupancy(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerServer virtualStealServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_virtualStealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_1_ctrl_serveStealReq_ready),
		.io_connNetwork_data_availableTask_ready(_virtualStealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNW_TQ_io_connVSS_1_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNW_TQ_io_connVSS_1_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNW_TQ_io_connVSS_1_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_virtualStealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_virtualStealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vss_1_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vss_1_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vss_1_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vss_1_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vss_1_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vss_1_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vss_1_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vss_1_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vss_1_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vss_1_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vss_1_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vss_1_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vss_1_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vss_1_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vss_1_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vss_1_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vss_1_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vss_1_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vss_1_b_bits_resp),
		.io_read_address_ready(_vssRvm_1_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_1_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_1_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_1_io_read_data_ready),
		.io_read_data_valid(_vssRvm_1_io_read_data_valid),
		.io_read_data_bits(_vssRvm_1_io_read_data_bits),
		.io_read_burst_len(_virtualStealServers_1_io_read_burst_len),
		.io_write_address_ready(_vssRvm_1_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_1_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_1_io_write_address_bits),
		.io_write_data_ready(_vssRvm_1_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_1_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_1_io_write_data_bits),
		.io_write_burst_len(_virtualStealServers_1_io_write_burst_len),
		.io_write_last(_virtualStealServers_1_io_write_last),
		.io_ntwDataUnitOccupancy(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_1)
	);
	RVtoAXIBridge vssRvm_0(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_writeBurst_len(_virtualStealServers_0_io_write_burst_len),
		.io_writeBurst_last(_virtualStealServers_0_io_write_last),
		.io_readBurst_len(_virtualStealServers_0_io_read_burst_len),
		.axi_ar_ready(_module_s_axi_ar_ready),
		.axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.axi_r_ready(_vssRvm_0_axi_r_ready),
		.axi_r_valid(_module_s_axi_r_valid),
		.axi_r_bits_data(_module_s_axi_r_bits_data),
		.axi_aw_ready(_module_s_axi_aw_ready),
		.axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.axi_aw_bits_len(_vssRvm_0_axi_aw_bits_len),
		.axi_w_ready(_module_s_axi_w_ready),
		.axi_w_valid(_vssRvm_0_axi_w_valid),
		.axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.axi_b_valid(_module_s_axi_b_valid)
	);
	RVtoAXIBridge vssRvm_1(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_vssRvm_1_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_1_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_1_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_1_io_read_data_ready),
		.io_read_data_valid(_vssRvm_1_io_read_data_valid),
		.io_read_data_bits(_vssRvm_1_io_read_data_bits),
		.io_write_address_ready(_vssRvm_1_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_1_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_1_io_write_address_bits),
		.io_write_data_ready(_vssRvm_1_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_1_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_1_io_write_data_bits),
		.io_writeBurst_len(_virtualStealServers_1_io_write_burst_len),
		.io_writeBurst_last(_virtualStealServers_1_io_write_last),
		.io_readBurst_len(_virtualStealServers_1_io_read_burst_len),
		.axi_ar_ready(_module_1_s_axi_ar_ready),
		.axi_ar_valid(_vssRvm_1_axi_ar_valid),
		.axi_ar_bits_addr(_vssRvm_1_axi_ar_bits_addr),
		.axi_ar_bits_len(_vssRvm_1_axi_ar_bits_len),
		.axi_r_ready(_vssRvm_1_axi_r_ready),
		.axi_r_valid(_module_1_s_axi_r_valid),
		.axi_r_bits_data(_module_1_s_axi_r_bits_data),
		.axi_aw_ready(_module_1_s_axi_aw_ready),
		.axi_aw_valid(_vssRvm_1_axi_aw_valid),
		.axi_aw_bits_addr(_vssRvm_1_axi_aw_bits_addr),
		.axi_aw_bits_len(_vssRvm_1_axi_aw_bits_len),
		.axi_w_ready(_module_1_s_axi_w_ready),
		.axi_w_valid(_vssRvm_1_axi_w_valid),
		.axi_w_bits_data(_vssRvm_1_axi_w_bits_data),
		.axi_w_bits_last(_vssRvm_1_axi_w_bits_last),
		.axi_b_valid(_module_1_s_axi_b_valid)
	);
	axi4FullMux mux(
		.clock(clock),
		.reset(reset),
		.s_axi_0_ar_ready(_mux_s_axi_0_ar_ready),
		.s_axi_0_ar_valid(_module_m_axi_ar_valid),
		.s_axi_0_ar_bits_addr(_module_m_axi_ar_bits_addr),
		.s_axi_0_ar_bits_len(_module_m_axi_ar_bits_len),
		.s_axi_0_ar_bits_size(_module_m_axi_ar_bits_size),
		.s_axi_0_ar_bits_burst(_module_m_axi_ar_bits_burst),
		.s_axi_0_ar_bits_lock(_module_m_axi_ar_bits_lock),
		.s_axi_0_ar_bits_cache(_module_m_axi_ar_bits_cache),
		.s_axi_0_ar_bits_prot(_module_m_axi_ar_bits_prot),
		.s_axi_0_ar_bits_qos(_module_m_axi_ar_bits_qos),
		.s_axi_0_ar_bits_region(_module_m_axi_ar_bits_region),
		.s_axi_0_r_ready(_module_m_axi_r_ready),
		.s_axi_0_r_valid(_mux_s_axi_0_r_valid),
		.s_axi_0_r_bits_data(_mux_s_axi_0_r_bits_data),
		.s_axi_0_aw_ready(_mux_s_axi_0_aw_ready),
		.s_axi_0_aw_valid(_module_m_axi_aw_valid),
		.s_axi_0_aw_bits_addr(_module_m_axi_aw_bits_addr),
		.s_axi_0_aw_bits_len(_module_m_axi_aw_bits_len),
		.s_axi_0_aw_bits_size(_module_m_axi_aw_bits_size),
		.s_axi_0_aw_bits_burst(_module_m_axi_aw_bits_burst),
		.s_axi_0_aw_bits_lock(_module_m_axi_aw_bits_lock),
		.s_axi_0_aw_bits_cache(_module_m_axi_aw_bits_cache),
		.s_axi_0_aw_bits_prot(_module_m_axi_aw_bits_prot),
		.s_axi_0_aw_bits_qos(_module_m_axi_aw_bits_qos),
		.s_axi_0_aw_bits_region(_module_m_axi_aw_bits_region),
		.s_axi_0_w_ready(_mux_s_axi_0_w_ready),
		.s_axi_0_w_valid(_module_m_axi_w_valid),
		.s_axi_0_w_bits_data(_module_m_axi_w_bits_data),
		.s_axi_0_w_bits_last(_module_m_axi_w_bits_last),
		.s_axi_0_b_valid(_mux_s_axi_0_b_valid),
		.s_axi_1_ar_ready(_mux_s_axi_1_ar_ready),
		.s_axi_1_ar_valid(_module_1_m_axi_ar_valid),
		.s_axi_1_ar_bits_addr(_module_1_m_axi_ar_bits_addr),
		.s_axi_1_ar_bits_len(_module_1_m_axi_ar_bits_len),
		.s_axi_1_ar_bits_size(_module_1_m_axi_ar_bits_size),
		.s_axi_1_ar_bits_burst(_module_1_m_axi_ar_bits_burst),
		.s_axi_1_ar_bits_lock(_module_1_m_axi_ar_bits_lock),
		.s_axi_1_ar_bits_cache(_module_1_m_axi_ar_bits_cache),
		.s_axi_1_ar_bits_prot(_module_1_m_axi_ar_bits_prot),
		.s_axi_1_ar_bits_qos(_module_1_m_axi_ar_bits_qos),
		.s_axi_1_ar_bits_region(_module_1_m_axi_ar_bits_region),
		.s_axi_1_r_ready(_module_1_m_axi_r_ready),
		.s_axi_1_r_valid(_mux_s_axi_1_r_valid),
		.s_axi_1_r_bits_data(_mux_s_axi_1_r_bits_data),
		.s_axi_1_aw_ready(_mux_s_axi_1_aw_ready),
		.s_axi_1_aw_valid(_module_1_m_axi_aw_valid),
		.s_axi_1_aw_bits_addr(_module_1_m_axi_aw_bits_addr),
		.s_axi_1_aw_bits_len(_module_1_m_axi_aw_bits_len),
		.s_axi_1_aw_bits_size(_module_1_m_axi_aw_bits_size),
		.s_axi_1_aw_bits_burst(_module_1_m_axi_aw_bits_burst),
		.s_axi_1_aw_bits_lock(_module_1_m_axi_aw_bits_lock),
		.s_axi_1_aw_bits_cache(_module_1_m_axi_aw_bits_cache),
		.s_axi_1_aw_bits_prot(_module_1_m_axi_aw_bits_prot),
		.s_axi_1_aw_bits_qos(_module_1_m_axi_aw_bits_qos),
		.s_axi_1_aw_bits_region(_module_1_m_axi_aw_bits_region),
		.s_axi_1_w_ready(_mux_s_axi_1_w_ready),
		.s_axi_1_w_valid(_module_1_m_axi_w_valid),
		.s_axi_1_w_bits_data(_module_1_m_axi_w_bits_data),
		.s_axi_1_w_bits_last(_module_1_m_axi_w_bits_last),
		.s_axi_1_b_valid(_mux_s_axi_1_b_valid),
		.m_axi_ar_ready(io_internal_vss_axi_full_0_ar_ready),
		.m_axi_ar_valid(io_internal_vss_axi_full_0_ar_valid),
		.m_axi_ar_bits_id(io_internal_vss_axi_full_0_ar_bits_id),
		.m_axi_ar_bits_addr(io_internal_vss_axi_full_0_ar_bits_addr),
		.m_axi_ar_bits_len(io_internal_vss_axi_full_0_ar_bits_len),
		.m_axi_ar_bits_size(io_internal_vss_axi_full_0_ar_bits_size),
		.m_axi_ar_bits_burst(io_internal_vss_axi_full_0_ar_bits_burst),
		.m_axi_ar_bits_lock(io_internal_vss_axi_full_0_ar_bits_lock),
		.m_axi_ar_bits_cache(io_internal_vss_axi_full_0_ar_bits_cache),
		.m_axi_ar_bits_prot(io_internal_vss_axi_full_0_ar_bits_prot),
		.m_axi_ar_bits_qos(io_internal_vss_axi_full_0_ar_bits_qos),
		.m_axi_ar_bits_region(io_internal_vss_axi_full_0_ar_bits_region),
		.m_axi_r_ready(io_internal_vss_axi_full_0_r_ready),
		.m_axi_r_valid(io_internal_vss_axi_full_0_r_valid),
		.m_axi_r_bits_id(io_internal_vss_axi_full_0_r_bits_id),
		.m_axi_r_bits_data(io_internal_vss_axi_full_0_r_bits_data),
		.m_axi_r_bits_resp(io_internal_vss_axi_full_0_r_bits_resp),
		.m_axi_r_bits_last(io_internal_vss_axi_full_0_r_bits_last),
		.m_axi_aw_ready(io_internal_vss_axi_full_0_aw_ready),
		.m_axi_aw_valid(io_internal_vss_axi_full_0_aw_valid),
		.m_axi_aw_bits_id(io_internal_vss_axi_full_0_aw_bits_id),
		.m_axi_aw_bits_addr(io_internal_vss_axi_full_0_aw_bits_addr),
		.m_axi_aw_bits_len(io_internal_vss_axi_full_0_aw_bits_len),
		.m_axi_aw_bits_size(io_internal_vss_axi_full_0_aw_bits_size),
		.m_axi_aw_bits_burst(io_internal_vss_axi_full_0_aw_bits_burst),
		.m_axi_aw_bits_lock(io_internal_vss_axi_full_0_aw_bits_lock),
		.m_axi_aw_bits_cache(io_internal_vss_axi_full_0_aw_bits_cache),
		.m_axi_aw_bits_prot(io_internal_vss_axi_full_0_aw_bits_prot),
		.m_axi_aw_bits_qos(io_internal_vss_axi_full_0_aw_bits_qos),
		.m_axi_aw_bits_region(io_internal_vss_axi_full_0_aw_bits_region),
		.m_axi_w_ready(io_internal_vss_axi_full_0_w_ready),
		.m_axi_w_valid(io_internal_vss_axi_full_0_w_valid),
		.m_axi_w_bits_data(io_internal_vss_axi_full_0_w_bits_data),
		.m_axi_w_bits_strb(io_internal_vss_axi_full_0_w_bits_strb),
		.m_axi_w_bits_last(io_internal_vss_axi_full_0_w_bits_last),
		.m_axi_b_ready(io_internal_vss_axi_full_0_b_ready),
		.m_axi_b_valid(io_internal_vss_axi_full_0_b_valid),
		.m_axi_b_bits_id(io_internal_vss_axi_full_0_b_bits_id),
		.m_axi_b_bits_resp(io_internal_vss_axi_full_0_b_bits_resp)
	);
	AxiWriteBuffer module_0(
		.clock(clock),
		.reset(reset),
		.s_axi_ar_ready(_module_s_axi_ar_ready),
		.s_axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.s_axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.s_axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.s_axi_r_ready(_vssRvm_0_axi_r_ready),
		.s_axi_r_valid(_module_s_axi_r_valid),
		.s_axi_r_bits_data(_module_s_axi_r_bits_data),
		.s_axi_aw_ready(_module_s_axi_aw_ready),
		.s_axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.s_axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.s_axi_aw_bits_len(_vssRvm_0_axi_aw_bits_len),
		.s_axi_w_ready(_module_s_axi_w_ready),
		.s_axi_w_valid(_vssRvm_0_axi_w_valid),
		.s_axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.s_axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.s_axi_b_valid(_module_s_axi_b_valid),
		.m_axi_ar_ready(_mux_s_axi_0_ar_ready),
		.m_axi_ar_valid(_module_m_axi_ar_valid),
		.m_axi_ar_bits_addr(_module_m_axi_ar_bits_addr),
		.m_axi_ar_bits_len(_module_m_axi_ar_bits_len),
		.m_axi_ar_bits_size(_module_m_axi_ar_bits_size),
		.m_axi_ar_bits_burst(_module_m_axi_ar_bits_burst),
		.m_axi_ar_bits_lock(_module_m_axi_ar_bits_lock),
		.m_axi_ar_bits_cache(_module_m_axi_ar_bits_cache),
		.m_axi_ar_bits_prot(_module_m_axi_ar_bits_prot),
		.m_axi_ar_bits_qos(_module_m_axi_ar_bits_qos),
		.m_axi_ar_bits_region(_module_m_axi_ar_bits_region),
		.m_axi_r_ready(_module_m_axi_r_ready),
		.m_axi_r_valid(_mux_s_axi_0_r_valid),
		.m_axi_r_bits_data(_mux_s_axi_0_r_bits_data),
		.m_axi_aw_ready(_mux_s_axi_0_aw_ready),
		.m_axi_aw_valid(_module_m_axi_aw_valid),
		.m_axi_aw_bits_addr(_module_m_axi_aw_bits_addr),
		.m_axi_aw_bits_len(_module_m_axi_aw_bits_len),
		.m_axi_aw_bits_size(_module_m_axi_aw_bits_size),
		.m_axi_aw_bits_burst(_module_m_axi_aw_bits_burst),
		.m_axi_aw_bits_lock(_module_m_axi_aw_bits_lock),
		.m_axi_aw_bits_cache(_module_m_axi_aw_bits_cache),
		.m_axi_aw_bits_prot(_module_m_axi_aw_bits_prot),
		.m_axi_aw_bits_qos(_module_m_axi_aw_bits_qos),
		.m_axi_aw_bits_region(_module_m_axi_aw_bits_region),
		.m_axi_w_ready(_mux_s_axi_0_w_ready),
		.m_axi_w_valid(_module_m_axi_w_valid),
		.m_axi_w_bits_data(_module_m_axi_w_bits_data),
		.m_axi_w_bits_last(_module_m_axi_w_bits_last),
		.m_axi_b_valid(_mux_s_axi_0_b_valid)
	);
	AxiWriteBuffer module_1(
		.clock(clock),
		.reset(reset),
		.s_axi_ar_ready(_module_1_s_axi_ar_ready),
		.s_axi_ar_valid(_vssRvm_1_axi_ar_valid),
		.s_axi_ar_bits_addr(_vssRvm_1_axi_ar_bits_addr),
		.s_axi_ar_bits_len(_vssRvm_1_axi_ar_bits_len),
		.s_axi_r_ready(_vssRvm_1_axi_r_ready),
		.s_axi_r_valid(_module_1_s_axi_r_valid),
		.s_axi_r_bits_data(_module_1_s_axi_r_bits_data),
		.s_axi_aw_ready(_module_1_s_axi_aw_ready),
		.s_axi_aw_valid(_vssRvm_1_axi_aw_valid),
		.s_axi_aw_bits_addr(_vssRvm_1_axi_aw_bits_addr),
		.s_axi_aw_bits_len(_vssRvm_1_axi_aw_bits_len),
		.s_axi_w_ready(_module_1_s_axi_w_ready),
		.s_axi_w_valid(_vssRvm_1_axi_w_valid),
		.s_axi_w_bits_data(_vssRvm_1_axi_w_bits_data),
		.s_axi_w_bits_last(_vssRvm_1_axi_w_bits_last),
		.s_axi_b_valid(_module_1_s_axi_b_valid),
		.m_axi_ar_ready(_mux_s_axi_1_ar_ready),
		.m_axi_ar_valid(_module_1_m_axi_ar_valid),
		.m_axi_ar_bits_addr(_module_1_m_axi_ar_bits_addr),
		.m_axi_ar_bits_len(_module_1_m_axi_ar_bits_len),
		.m_axi_ar_bits_size(_module_1_m_axi_ar_bits_size),
		.m_axi_ar_bits_burst(_module_1_m_axi_ar_bits_burst),
		.m_axi_ar_bits_lock(_module_1_m_axi_ar_bits_lock),
		.m_axi_ar_bits_cache(_module_1_m_axi_ar_bits_cache),
		.m_axi_ar_bits_prot(_module_1_m_axi_ar_bits_prot),
		.m_axi_ar_bits_qos(_module_1_m_axi_ar_bits_qos),
		.m_axi_ar_bits_region(_module_1_m_axi_ar_bits_region),
		.m_axi_r_ready(_module_1_m_axi_r_ready),
		.m_axi_r_valid(_mux_s_axi_1_r_valid),
		.m_axi_r_bits_data(_mux_s_axi_1_r_bits_data),
		.m_axi_aw_ready(_mux_s_axi_1_aw_ready),
		.m_axi_aw_valid(_module_1_m_axi_aw_valid),
		.m_axi_aw_bits_addr(_module_1_m_axi_aw_bits_addr),
		.m_axi_aw_bits_len(_module_1_m_axi_aw_bits_len),
		.m_axi_aw_bits_size(_module_1_m_axi_aw_bits_size),
		.m_axi_aw_bits_burst(_module_1_m_axi_aw_bits_burst),
		.m_axi_aw_bits_lock(_module_1_m_axi_aw_bits_lock),
		.m_axi_aw_bits_cache(_module_1_m_axi_aw_bits_cache),
		.m_axi_aw_bits_prot(_module_1_m_axi_aw_bits_prot),
		.m_axi_aw_bits_qos(_module_1_m_axi_aw_bits_qos),
		.m_axi_aw_bits_region(_module_1_m_axi_aw_bits_region),
		.m_axi_w_ready(_mux_s_axi_1_w_ready),
		.m_axi_w_valid(_module_1_m_axi_w_valid),
		.m_axi_w_bits_data(_module_1_m_axi_w_bits_data),
		.m_axi_w_bits_last(_module_1_m_axi_w_bits_last),
		.m_axi_b_valid(_mux_s_axi_1_b_valid)
	);
	AxisDataWidthConverter axis_stream_converters_out_0(
		.io_dataIn_TREADY(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_0_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_0_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_0_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_0_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_1(
		.io_dataIn_TREADY(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_1_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_1_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_1_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_1_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_2(
		.io_dataIn_TREADY(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_2_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_2_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_2_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_2_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_3(
		.io_dataIn_TREADY(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_3_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_3_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_3_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_3_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_4(
		.io_dataIn_TREADY(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_4_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_4_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_4_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_4_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_5(
		.io_dataIn_TREADY(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_5_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_5_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_5_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_5_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_6(
		.io_dataIn_TREADY(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_6_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_6_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_6_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_6_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_7(
		.io_dataIn_TREADY(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_7_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_7_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_7_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_7_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_8(
		.io_dataIn_TREADY(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_8_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_8_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_8_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_8_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_9(
		.io_dataIn_TREADY(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_9_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_9_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_9_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_9_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_10(
		.io_dataIn_TREADY(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_10_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_10_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_10_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_10_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_11(
		.io_dataIn_TREADY(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_11_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_11_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_11_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_11_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_12(
		.io_dataIn_TREADY(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_12_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_12_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_12_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_12_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_13(
		.io_dataIn_TREADY(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_13_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_13_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_13_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_13_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_14(
		.io_dataIn_TREADY(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_14_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_14_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_14_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_14_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_15(
		.io_dataIn_TREADY(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_15_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_15_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_15_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_15_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_16(
		.io_dataIn_TREADY(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_16_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_16_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_16_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_16_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_16_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_17(
		.io_dataIn_TREADY(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_17_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_17_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_17_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_17_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_17_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_18(
		.io_dataIn_TREADY(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_18_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_18_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_18_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_18_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_18_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_19(
		.io_dataIn_TREADY(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_19_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_19_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_19_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_19_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_19_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_20(
		.io_dataIn_TREADY(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_20_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_20_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_20_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_20_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_20_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_21(
		.io_dataIn_TREADY(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_21_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_21_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_21_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_21_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_21_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_22(
		.io_dataIn_TREADY(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_22_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_22_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_22_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_22_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_22_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_23(
		.io_dataIn_TREADY(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_23_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_23_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_23_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_23_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_23_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_24(
		.io_dataIn_TREADY(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_24_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_24_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_24_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_24_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_24_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_25(
		.io_dataIn_TREADY(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_25_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_25_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_25_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_25_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_25_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_26(
		.io_dataIn_TREADY(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_26_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_26_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_26_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_26_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_26_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_27(
		.io_dataIn_TREADY(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_27_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_27_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_27_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_27_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_27_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_28(
		.io_dataIn_TREADY(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_28_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_28_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_28_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_28_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_28_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_29(
		.io_dataIn_TREADY(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_29_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_29_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_29_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_29_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_29_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_30(
		.io_dataIn_TREADY(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_30_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_30_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_30_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_30_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_30_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_31(
		.io_dataIn_TREADY(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_31_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_31_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_31_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_31_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_31_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_32(
		.io_dataIn_TREADY(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_32_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_32_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_32_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_32_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_32_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_33(
		.io_dataIn_TREADY(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_33_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_33_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_33_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_33_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_33_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_34(
		.io_dataIn_TREADY(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_34_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_34_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_34_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_34_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_34_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_35(
		.io_dataIn_TREADY(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_35_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_35_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_35_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_35_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_35_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_36(
		.io_dataIn_TREADY(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_36_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_36_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_36_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_36_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_36_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_37(
		.io_dataIn_TREADY(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_37_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_37_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_37_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_37_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_37_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_38(
		.io_dataIn_TREADY(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_38_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_38_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_38_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_38_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_38_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_39(
		.io_dataIn_TREADY(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_39_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_39_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_39_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_39_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_39_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_40(
		.io_dataIn_TREADY(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_40_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_40_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_40_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_40_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_40_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_41(
		.io_dataIn_TREADY(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_41_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_41_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_41_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_41_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_41_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_42(
		.io_dataIn_TREADY(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_42_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_42_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_42_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_42_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_42_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_43(
		.io_dataIn_TREADY(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_43_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_43_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_43_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_43_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_43_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_44(
		.io_dataIn_TREADY(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_44_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_44_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_44_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_44_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_44_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_45(
		.io_dataIn_TREADY(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_45_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_45_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_45_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_45_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_45_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_46(
		.io_dataIn_TREADY(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_46_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_46_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_46_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_46_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_46_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_47(
		.io_dataIn_TREADY(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_47_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_47_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_47_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_47_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_47_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_48(
		.io_dataIn_TREADY(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_48_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_48_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_48_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_48_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_48_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_49(
		.io_dataIn_TREADY(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_49_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_49_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_49_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_49_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_49_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_50(
		.io_dataIn_TREADY(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_50_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_50_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_50_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_50_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_50_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_51(
		.io_dataIn_TREADY(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_51_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_51_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_51_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_51_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_51_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_52(
		.io_dataIn_TREADY(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_52_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_52_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_52_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_52_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_52_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_53(
		.io_dataIn_TREADY(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_53_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_53_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_53_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_53_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_53_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_54(
		.io_dataIn_TREADY(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_54_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_54_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_54_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_54_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_54_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_55(
		.io_dataIn_TREADY(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_55_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_55_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_55_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_55_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_55_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_56(
		.io_dataIn_TREADY(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_56_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_56_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_56_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_56_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_56_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_57(
		.io_dataIn_TREADY(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_57_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_57_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_57_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_57_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_57_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_58(
		.io_dataIn_TREADY(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_58_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_58_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_58_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_58_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_58_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_59(
		.io_dataIn_TREADY(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_59_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_59_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_59_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_59_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_59_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_60(
		.io_dataIn_TREADY(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_60_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_60_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_60_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_60_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_60_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_61(
		.io_dataIn_TREADY(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_61_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_61_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_61_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_61_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_61_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_62(
		.io_dataIn_TREADY(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_62_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_62_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_62_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_62_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_62_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_out_63(
		.io_dataIn_TREADY(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_63_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_63_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_63_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_63_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_63_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_0(
		.io_dataIn_TREADY(io_export_taskIn_0_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_0_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_0_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_0_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_0_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_1(
		.io_dataIn_TREADY(io_export_taskIn_1_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_1_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_1_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_1_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_1_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_2(
		.io_dataIn_TREADY(io_export_taskIn_2_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_2_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_2_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_2_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_2_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_3(
		.io_dataIn_TREADY(io_export_taskIn_3_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_3_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_3_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_3_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_3_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_4(
		.io_dataIn_TREADY(io_export_taskIn_4_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_4_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_4_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_4_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_4_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_5(
		.io_dataIn_TREADY(io_export_taskIn_5_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_5_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_5_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_5_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_5_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_6(
		.io_dataIn_TREADY(io_export_taskIn_6_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_6_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_6_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_6_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_6_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_7(
		.io_dataIn_TREADY(io_export_taskIn_7_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_7_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_7_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_7_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_7_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_8(
		.io_dataIn_TREADY(io_export_taskIn_8_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_8_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_8_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_8_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_8_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_9(
		.io_dataIn_TREADY(io_export_taskIn_9_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_9_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_9_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_9_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_9_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_10(
		.io_dataIn_TREADY(io_export_taskIn_10_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_10_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_10_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_10_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_10_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_11(
		.io_dataIn_TREADY(io_export_taskIn_11_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_11_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_11_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_11_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_11_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_12(
		.io_dataIn_TREADY(io_export_taskIn_12_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_12_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_12_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_12_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_12_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_13(
		.io_dataIn_TREADY(io_export_taskIn_13_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_13_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_13_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_13_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_13_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_14(
		.io_dataIn_TREADY(io_export_taskIn_14_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_14_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_14_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_14_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_14_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_15(
		.io_dataIn_TREADY(io_export_taskIn_15_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_15_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_15_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_15_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_15_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_16(
		.io_dataIn_TREADY(io_export_taskIn_16_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_16_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_16_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_16_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_16_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_17(
		.io_dataIn_TREADY(io_export_taskIn_17_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_17_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_17_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_17_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_17_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_18(
		.io_dataIn_TREADY(io_export_taskIn_18_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_18_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_18_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_18_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_18_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_19(
		.io_dataIn_TREADY(io_export_taskIn_19_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_19_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_19_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_19_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_19_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_20(
		.io_dataIn_TREADY(io_export_taskIn_20_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_20_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_20_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_20_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_20_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_21(
		.io_dataIn_TREADY(io_export_taskIn_21_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_21_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_21_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_21_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_21_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_22(
		.io_dataIn_TREADY(io_export_taskIn_22_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_22_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_22_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_22_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_22_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_23(
		.io_dataIn_TREADY(io_export_taskIn_23_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_23_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_23_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_23_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_23_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_24(
		.io_dataIn_TREADY(io_export_taskIn_24_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_24_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_24_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_24_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_24_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_25(
		.io_dataIn_TREADY(io_export_taskIn_25_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_25_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_25_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_25_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_25_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_26(
		.io_dataIn_TREADY(io_export_taskIn_26_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_26_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_26_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_26_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_26_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_27(
		.io_dataIn_TREADY(io_export_taskIn_27_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_27_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_27_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_27_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_27_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_28(
		.io_dataIn_TREADY(io_export_taskIn_28_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_28_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_28_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_28_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_28_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_29(
		.io_dataIn_TREADY(io_export_taskIn_29_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_29_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_29_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_29_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_29_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_30(
		.io_dataIn_TREADY(io_export_taskIn_30_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_30_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_30_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_30_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_30_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_31(
		.io_dataIn_TREADY(io_export_taskIn_31_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_31_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_31_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_31_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_31_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_32(
		.io_dataIn_TREADY(io_export_taskIn_32_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_32_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_32_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_32_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_32_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_33(
		.io_dataIn_TREADY(io_export_taskIn_33_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_33_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_33_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_33_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_33_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_34(
		.io_dataIn_TREADY(io_export_taskIn_34_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_34_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_34_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_34_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_34_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_35(
		.io_dataIn_TREADY(io_export_taskIn_35_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_35_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_35_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_35_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_35_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_36(
		.io_dataIn_TREADY(io_export_taskIn_36_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_36_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_36_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_36_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_36_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_37(
		.io_dataIn_TREADY(io_export_taskIn_37_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_37_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_37_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_37_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_37_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_38(
		.io_dataIn_TREADY(io_export_taskIn_38_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_38_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_38_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_38_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_38_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_39(
		.io_dataIn_TREADY(io_export_taskIn_39_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_39_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_39_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_39_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_39_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_40(
		.io_dataIn_TREADY(io_export_taskIn_40_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_40_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_40_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_40_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_40_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_41(
		.io_dataIn_TREADY(io_export_taskIn_41_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_41_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_41_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_41_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_41_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_42(
		.io_dataIn_TREADY(io_export_taskIn_42_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_42_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_42_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_42_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_42_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_43(
		.io_dataIn_TREADY(io_export_taskIn_43_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_43_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_43_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_43_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_43_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_44(
		.io_dataIn_TREADY(io_export_taskIn_44_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_44_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_44_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_44_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_44_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_45(
		.io_dataIn_TREADY(io_export_taskIn_45_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_45_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_45_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_45_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_45_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_46(
		.io_dataIn_TREADY(io_export_taskIn_46_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_46_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_46_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_46_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_46_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_47(
		.io_dataIn_TREADY(io_export_taskIn_47_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_47_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_47_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_47_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_47_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_48(
		.io_dataIn_TREADY(io_export_taskIn_48_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_48_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_48_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_48_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_48_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_49(
		.io_dataIn_TREADY(io_export_taskIn_49_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_49_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_49_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_49_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_49_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_50(
		.io_dataIn_TREADY(io_export_taskIn_50_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_50_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_50_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_50_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_50_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_51(
		.io_dataIn_TREADY(io_export_taskIn_51_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_51_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_51_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_51_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_51_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_52(
		.io_dataIn_TREADY(io_export_taskIn_52_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_52_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_52_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_52_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_52_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_53(
		.io_dataIn_TREADY(io_export_taskIn_53_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_53_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_53_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_53_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_53_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_54(
		.io_dataIn_TREADY(io_export_taskIn_54_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_54_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_54_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_54_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_54_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_55(
		.io_dataIn_TREADY(io_export_taskIn_55_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_55_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_55_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_55_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_55_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_56(
		.io_dataIn_TREADY(io_export_taskIn_56_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_56_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_56_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_56_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_56_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_57(
		.io_dataIn_TREADY(io_export_taskIn_57_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_57_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_57_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_57_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_57_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_58(
		.io_dataIn_TREADY(io_export_taskIn_58_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_58_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_58_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_58_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_58_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_59(
		.io_dataIn_TREADY(io_export_taskIn_59_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_59_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_59_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_59_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_59_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_60(
		.io_dataIn_TREADY(io_export_taskIn_60_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_60_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_60_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_60_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_60_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_61(
		.io_dataIn_TREADY(io_export_taskIn_61_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_61_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_61_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_61_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_61_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_62(
		.io_dataIn_TREADY(io_export_taskIn_62_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_62_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_62_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_62_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_62_io_dataOut_TDATA)
	);
	AxisDataWidthConverter axis_stream_converters_in_63(
		.io_dataIn_TREADY(io_export_taskIn_63_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_63_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_63_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_63_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_63_io_dataOut_TDATA)
	);
endmodule
module SchedulerNetworkDataUnit_66 (
	clock,
	reset,
	io_taskIn,
	io_taskOut,
	io_validIn,
	io_validOut,
	io_connSS_availableTask_ready,
	io_connSS_availableTask_valid,
	io_connSS_availableTask_bits,
	io_connSS_qOutTask_ready,
	io_connSS_qOutTask_valid,
	io_connSS_qOutTask_bits,
	io_occupied
);
	input clock;
	input reset;
	input [255:0] io_taskIn;
	output wire [255:0] io_taskOut;
	input io_validIn;
	output wire io_validOut;
	input io_connSS_availableTask_ready;
	output wire io_connSS_availableTask_valid;
	output wire [255:0] io_connSS_availableTask_bits;
	output wire io_connSS_qOutTask_ready;
	input io_connSS_qOutTask_valid;
	input [255:0] io_connSS_qOutTask_bits;
	output wire io_occupied;
	reg [255:0] taskReg;
	reg validReg;
	wire io_connSS_availableTask_valid_0 = io_connSS_availableTask_ready & io_validIn;
	wire _GEN = io_connSS_qOutTask_valid & ~io_validIn;
	always @(posedge clock)
		if (reset) begin
			taskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			validReg <= 1'h0;
		end
		else begin
			taskReg <= (io_connSS_availableTask_valid_0 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : (_GEN ? io_connSS_qOutTask_bits : (io_validIn ? io_taskIn : 256'h0000000000000000000000000000000000000000000000000000000000000000)));
			validReg <= ~io_connSS_availableTask_valid_0 & (_GEN | io_validIn);
		end
	assign io_taskOut = taskReg;
	assign io_validOut = validReg;
	assign io_connSS_availableTask_valid = io_connSS_availableTask_valid_0;
	assign io_connSS_availableTask_bits = (io_connSS_availableTask_valid_0 ? io_taskIn : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	assign io_connSS_qOutTask_ready = ~io_connSS_availableTask_valid_0 & _GEN;
	assign io_occupied = validReg;
endmodule
module SchedulerNetwork_1 (
	clock,
	reset,
	io_connSS_0_ctrl_serveStealReq_valid,
	io_connSS_0_ctrl_serveStealReq_ready,
	io_connSS_0_data_availableTask_ready,
	io_connSS_0_data_availableTask_valid,
	io_connSS_0_data_availableTask_bits,
	io_connSS_0_data_qOutTask_ready,
	io_connSS_0_data_qOutTask_valid,
	io_connSS_0_data_qOutTask_bits,
	io_connSS_1_ctrl_serveStealReq_valid,
	io_connSS_1_ctrl_serveStealReq_ready,
	io_connSS_1_data_availableTask_ready,
	io_connSS_1_data_availableTask_valid,
	io_connSS_1_data_availableTask_bits,
	io_connSS_1_data_qOutTask_ready,
	io_connSS_1_data_qOutTask_valid,
	io_connSS_1_data_qOutTask_bits,
	io_connSS_2_ctrl_serveStealReq_valid,
	io_connSS_2_ctrl_serveStealReq_ready,
	io_connSS_2_data_qOutTask_ready,
	io_connSS_2_data_qOutTask_valid,
	io_connSS_2_data_qOutTask_bits,
	io_connSS_3_ctrl_serveStealReq_valid,
	io_connSS_3_ctrl_serveStealReq_ready,
	io_connSS_3_data_qOutTask_ready,
	io_connSS_3_data_qOutTask_valid,
	io_connSS_3_data_qOutTask_bits,
	io_connSS_4_ctrl_serveStealReq_valid,
	io_connSS_4_ctrl_serveStealReq_ready,
	io_connSS_4_data_qOutTask_ready,
	io_connSS_4_data_qOutTask_valid,
	io_connSS_4_data_qOutTask_bits,
	io_connSS_5_ctrl_serveStealReq_valid,
	io_connSS_5_ctrl_serveStealReq_ready,
	io_connSS_5_data_qOutTask_ready,
	io_connSS_5_data_qOutTask_valid,
	io_connSS_5_data_qOutTask_bits,
	io_connSS_6_ctrl_serveStealReq_valid,
	io_connSS_6_ctrl_serveStealReq_ready,
	io_connSS_6_data_qOutTask_ready,
	io_connSS_6_data_qOutTask_valid,
	io_connSS_6_data_qOutTask_bits,
	io_connSS_7_ctrl_serveStealReq_valid,
	io_connSS_7_ctrl_serveStealReq_ready,
	io_connSS_7_data_qOutTask_ready,
	io_connSS_7_data_qOutTask_valid,
	io_connSS_7_data_qOutTask_bits,
	io_connSS_8_ctrl_serveStealReq_valid,
	io_connSS_8_ctrl_serveStealReq_ready,
	io_connSS_8_data_qOutTask_ready,
	io_connSS_8_data_qOutTask_valid,
	io_connSS_8_data_qOutTask_bits,
	io_connSS_9_ctrl_serveStealReq_valid,
	io_connSS_9_ctrl_serveStealReq_ready,
	io_connSS_9_data_qOutTask_ready,
	io_connSS_9_data_qOutTask_valid,
	io_connSS_9_data_qOutTask_bits,
	io_connSS_10_ctrl_serveStealReq_valid,
	io_connSS_10_ctrl_serveStealReq_ready,
	io_connSS_10_data_qOutTask_ready,
	io_connSS_10_data_qOutTask_valid,
	io_connSS_10_data_qOutTask_bits,
	io_connSS_11_ctrl_serveStealReq_valid,
	io_connSS_11_ctrl_serveStealReq_ready,
	io_connSS_11_data_qOutTask_ready,
	io_connSS_11_data_qOutTask_valid,
	io_connSS_11_data_qOutTask_bits,
	io_connSS_12_ctrl_serveStealReq_valid,
	io_connSS_12_ctrl_serveStealReq_ready,
	io_connSS_12_data_qOutTask_ready,
	io_connSS_12_data_qOutTask_valid,
	io_connSS_12_data_qOutTask_bits,
	io_connSS_13_ctrl_serveStealReq_valid,
	io_connSS_13_ctrl_serveStealReq_ready,
	io_connSS_13_data_qOutTask_ready,
	io_connSS_13_data_qOutTask_valid,
	io_connSS_13_data_qOutTask_bits,
	io_connSS_14_ctrl_serveStealReq_valid,
	io_connSS_14_ctrl_serveStealReq_ready,
	io_connSS_14_data_qOutTask_ready,
	io_connSS_14_data_qOutTask_valid,
	io_connSS_14_data_qOutTask_bits,
	io_connSS_15_ctrl_serveStealReq_valid,
	io_connSS_15_ctrl_serveStealReq_ready,
	io_connSS_15_data_qOutTask_ready,
	io_connSS_15_data_qOutTask_valid,
	io_connSS_15_data_qOutTask_bits,
	io_connSS_16_ctrl_serveStealReq_valid,
	io_connSS_16_ctrl_serveStealReq_ready,
	io_connSS_16_data_qOutTask_ready,
	io_connSS_16_data_qOutTask_valid,
	io_connSS_16_data_qOutTask_bits,
	io_connSS_17_ctrl_serveStealReq_valid,
	io_connSS_17_ctrl_serveStealReq_ready,
	io_connSS_17_data_qOutTask_ready,
	io_connSS_17_data_qOutTask_valid,
	io_connSS_17_data_qOutTask_bits,
	io_connSS_18_ctrl_serveStealReq_valid,
	io_connSS_18_ctrl_serveStealReq_ready,
	io_connSS_18_ctrl_stealReq_valid,
	io_connSS_18_ctrl_stealReq_ready,
	io_connSS_18_data_availableTask_ready,
	io_connSS_18_data_availableTask_valid,
	io_connSS_18_data_availableTask_bits,
	io_connSS_18_data_qOutTask_ready,
	io_connSS_18_data_qOutTask_valid,
	io_connSS_18_data_qOutTask_bits,
	io_connSS_19_ctrl_serveStealReq_valid,
	io_connSS_19_ctrl_serveStealReq_ready,
	io_connSS_19_ctrl_stealReq_valid,
	io_connSS_19_ctrl_stealReq_ready,
	io_connSS_19_data_availableTask_ready,
	io_connSS_19_data_availableTask_valid,
	io_connSS_19_data_availableTask_bits,
	io_connSS_19_data_qOutTask_ready,
	io_connSS_19_data_qOutTask_valid,
	io_connSS_19_data_qOutTask_bits,
	io_connSS_20_ctrl_serveStealReq_valid,
	io_connSS_20_ctrl_serveStealReq_ready,
	io_connSS_20_ctrl_stealReq_valid,
	io_connSS_20_ctrl_stealReq_ready,
	io_connSS_20_data_availableTask_ready,
	io_connSS_20_data_availableTask_valid,
	io_connSS_20_data_availableTask_bits,
	io_connSS_20_data_qOutTask_ready,
	io_connSS_20_data_qOutTask_valid,
	io_connSS_20_data_qOutTask_bits,
	io_connSS_21_ctrl_serveStealReq_valid,
	io_connSS_21_ctrl_serveStealReq_ready,
	io_connSS_21_ctrl_stealReq_valid,
	io_connSS_21_ctrl_stealReq_ready,
	io_connSS_21_data_availableTask_ready,
	io_connSS_21_data_availableTask_valid,
	io_connSS_21_data_availableTask_bits,
	io_connSS_21_data_qOutTask_ready,
	io_connSS_21_data_qOutTask_valid,
	io_connSS_21_data_qOutTask_bits,
	io_connSS_22_ctrl_serveStealReq_valid,
	io_connSS_22_ctrl_serveStealReq_ready,
	io_connSS_22_ctrl_stealReq_valid,
	io_connSS_22_ctrl_stealReq_ready,
	io_connSS_22_data_availableTask_ready,
	io_connSS_22_data_availableTask_valid,
	io_connSS_22_data_availableTask_bits,
	io_connSS_22_data_qOutTask_ready,
	io_connSS_22_data_qOutTask_valid,
	io_connSS_22_data_qOutTask_bits,
	io_connSS_23_ctrl_serveStealReq_valid,
	io_connSS_23_ctrl_serveStealReq_ready,
	io_connSS_23_ctrl_stealReq_valid,
	io_connSS_23_ctrl_stealReq_ready,
	io_connSS_23_data_availableTask_ready,
	io_connSS_23_data_availableTask_valid,
	io_connSS_23_data_availableTask_bits,
	io_connSS_23_data_qOutTask_ready,
	io_connSS_23_data_qOutTask_valid,
	io_connSS_23_data_qOutTask_bits,
	io_connSS_24_ctrl_serveStealReq_valid,
	io_connSS_24_ctrl_serveStealReq_ready,
	io_connSS_24_ctrl_stealReq_valid,
	io_connSS_24_ctrl_stealReq_ready,
	io_connSS_24_data_availableTask_ready,
	io_connSS_24_data_availableTask_valid,
	io_connSS_24_data_availableTask_bits,
	io_connSS_24_data_qOutTask_ready,
	io_connSS_24_data_qOutTask_valid,
	io_connSS_24_data_qOutTask_bits,
	io_connSS_25_ctrl_serveStealReq_valid,
	io_connSS_25_ctrl_serveStealReq_ready,
	io_connSS_25_ctrl_stealReq_valid,
	io_connSS_25_ctrl_stealReq_ready,
	io_connSS_25_data_availableTask_ready,
	io_connSS_25_data_availableTask_valid,
	io_connSS_25_data_availableTask_bits,
	io_connSS_25_data_qOutTask_ready,
	io_connSS_25_data_qOutTask_valid,
	io_connSS_25_data_qOutTask_bits,
	io_connSS_26_ctrl_serveStealReq_valid,
	io_connSS_26_ctrl_serveStealReq_ready,
	io_connSS_26_ctrl_stealReq_valid,
	io_connSS_26_ctrl_stealReq_ready,
	io_connSS_26_data_availableTask_ready,
	io_connSS_26_data_availableTask_valid,
	io_connSS_26_data_availableTask_bits,
	io_connSS_26_data_qOutTask_ready,
	io_connSS_26_data_qOutTask_valid,
	io_connSS_26_data_qOutTask_bits,
	io_connSS_27_ctrl_serveStealReq_valid,
	io_connSS_27_ctrl_serveStealReq_ready,
	io_connSS_27_ctrl_stealReq_valid,
	io_connSS_27_ctrl_stealReq_ready,
	io_connSS_27_data_availableTask_ready,
	io_connSS_27_data_availableTask_valid,
	io_connSS_27_data_availableTask_bits,
	io_connSS_27_data_qOutTask_ready,
	io_connSS_27_data_qOutTask_valid,
	io_connSS_27_data_qOutTask_bits,
	io_connSS_28_ctrl_serveStealReq_valid,
	io_connSS_28_ctrl_serveStealReq_ready,
	io_connSS_28_ctrl_stealReq_valid,
	io_connSS_28_ctrl_stealReq_ready,
	io_connSS_28_data_availableTask_ready,
	io_connSS_28_data_availableTask_valid,
	io_connSS_28_data_availableTask_bits,
	io_connSS_28_data_qOutTask_ready,
	io_connSS_28_data_qOutTask_valid,
	io_connSS_28_data_qOutTask_bits,
	io_connSS_29_ctrl_serveStealReq_valid,
	io_connSS_29_ctrl_serveStealReq_ready,
	io_connSS_29_ctrl_stealReq_valid,
	io_connSS_29_ctrl_stealReq_ready,
	io_connSS_29_data_availableTask_ready,
	io_connSS_29_data_availableTask_valid,
	io_connSS_29_data_availableTask_bits,
	io_connSS_29_data_qOutTask_ready,
	io_connSS_29_data_qOutTask_valid,
	io_connSS_29_data_qOutTask_bits,
	io_connSS_30_ctrl_serveStealReq_valid,
	io_connSS_30_ctrl_serveStealReq_ready,
	io_connSS_30_ctrl_stealReq_valid,
	io_connSS_30_ctrl_stealReq_ready,
	io_connSS_30_data_availableTask_ready,
	io_connSS_30_data_availableTask_valid,
	io_connSS_30_data_availableTask_bits,
	io_connSS_30_data_qOutTask_ready,
	io_connSS_30_data_qOutTask_valid,
	io_connSS_30_data_qOutTask_bits,
	io_connSS_31_ctrl_serveStealReq_valid,
	io_connSS_31_ctrl_serveStealReq_ready,
	io_connSS_31_ctrl_stealReq_valid,
	io_connSS_31_ctrl_stealReq_ready,
	io_connSS_31_data_availableTask_ready,
	io_connSS_31_data_availableTask_valid,
	io_connSS_31_data_availableTask_bits,
	io_connSS_31_data_qOutTask_ready,
	io_connSS_31_data_qOutTask_valid,
	io_connSS_31_data_qOutTask_bits,
	io_connSS_32_ctrl_serveStealReq_valid,
	io_connSS_32_ctrl_serveStealReq_ready,
	io_connSS_32_ctrl_stealReq_valid,
	io_connSS_32_ctrl_stealReq_ready,
	io_connSS_32_data_availableTask_ready,
	io_connSS_32_data_availableTask_valid,
	io_connSS_32_data_availableTask_bits,
	io_connSS_32_data_qOutTask_ready,
	io_connSS_32_data_qOutTask_valid,
	io_connSS_32_data_qOutTask_bits,
	io_connSS_33_ctrl_serveStealReq_valid,
	io_connSS_33_ctrl_serveStealReq_ready,
	io_connSS_33_ctrl_stealReq_valid,
	io_connSS_33_ctrl_stealReq_ready,
	io_connSS_33_data_availableTask_ready,
	io_connSS_33_data_availableTask_valid,
	io_connSS_33_data_availableTask_bits,
	io_connSS_33_data_qOutTask_ready,
	io_connSS_33_data_qOutTask_valid,
	io_connSS_33_data_qOutTask_bits,
	io_connSS_34_ctrl_serveStealReq_valid,
	io_connSS_34_ctrl_serveStealReq_ready,
	io_connSS_34_ctrl_stealReq_valid,
	io_connSS_34_ctrl_stealReq_ready,
	io_connSS_34_data_availableTask_ready,
	io_connSS_34_data_availableTask_valid,
	io_connSS_34_data_availableTask_bits,
	io_connSS_34_data_qOutTask_ready,
	io_connSS_34_data_qOutTask_valid,
	io_connSS_34_data_qOutTask_bits,
	io_connSS_35_ctrl_serveStealReq_valid,
	io_connSS_35_ctrl_serveStealReq_ready,
	io_connSS_35_ctrl_stealReq_valid,
	io_connSS_35_ctrl_stealReq_ready,
	io_connSS_35_data_availableTask_ready,
	io_connSS_35_data_availableTask_valid,
	io_connSS_35_data_availableTask_bits,
	io_connSS_35_data_qOutTask_ready,
	io_connSS_35_data_qOutTask_valid,
	io_connSS_35_data_qOutTask_bits,
	io_connSS_36_ctrl_serveStealReq_valid,
	io_connSS_36_ctrl_serveStealReq_ready,
	io_connSS_36_ctrl_stealReq_valid,
	io_connSS_36_ctrl_stealReq_ready,
	io_connSS_36_data_availableTask_ready,
	io_connSS_36_data_availableTask_valid,
	io_connSS_36_data_availableTask_bits,
	io_connSS_36_data_qOutTask_ready,
	io_connSS_36_data_qOutTask_valid,
	io_connSS_36_data_qOutTask_bits,
	io_connSS_37_ctrl_serveStealReq_valid,
	io_connSS_37_ctrl_serveStealReq_ready,
	io_connSS_37_ctrl_stealReq_valid,
	io_connSS_37_ctrl_stealReq_ready,
	io_connSS_37_data_availableTask_ready,
	io_connSS_37_data_availableTask_valid,
	io_connSS_37_data_availableTask_bits,
	io_connSS_37_data_qOutTask_ready,
	io_connSS_37_data_qOutTask_valid,
	io_connSS_37_data_qOutTask_bits,
	io_connSS_38_ctrl_serveStealReq_valid,
	io_connSS_38_ctrl_serveStealReq_ready,
	io_connSS_38_ctrl_stealReq_valid,
	io_connSS_38_ctrl_stealReq_ready,
	io_connSS_38_data_availableTask_ready,
	io_connSS_38_data_availableTask_valid,
	io_connSS_38_data_availableTask_bits,
	io_connSS_38_data_qOutTask_ready,
	io_connSS_38_data_qOutTask_valid,
	io_connSS_38_data_qOutTask_bits,
	io_connSS_39_ctrl_serveStealReq_valid,
	io_connSS_39_ctrl_serveStealReq_ready,
	io_connSS_39_ctrl_stealReq_valid,
	io_connSS_39_ctrl_stealReq_ready,
	io_connSS_39_data_availableTask_ready,
	io_connSS_39_data_availableTask_valid,
	io_connSS_39_data_availableTask_bits,
	io_connSS_39_data_qOutTask_ready,
	io_connSS_39_data_qOutTask_valid,
	io_connSS_39_data_qOutTask_bits,
	io_connSS_40_ctrl_serveStealReq_valid,
	io_connSS_40_ctrl_serveStealReq_ready,
	io_connSS_40_ctrl_stealReq_valid,
	io_connSS_40_ctrl_stealReq_ready,
	io_connSS_40_data_availableTask_ready,
	io_connSS_40_data_availableTask_valid,
	io_connSS_40_data_availableTask_bits,
	io_connSS_40_data_qOutTask_ready,
	io_connSS_40_data_qOutTask_valid,
	io_connSS_40_data_qOutTask_bits,
	io_connSS_41_ctrl_serveStealReq_valid,
	io_connSS_41_ctrl_serveStealReq_ready,
	io_connSS_41_ctrl_stealReq_valid,
	io_connSS_41_ctrl_stealReq_ready,
	io_connSS_41_data_availableTask_ready,
	io_connSS_41_data_availableTask_valid,
	io_connSS_41_data_availableTask_bits,
	io_connSS_41_data_qOutTask_ready,
	io_connSS_41_data_qOutTask_valid,
	io_connSS_41_data_qOutTask_bits,
	io_connSS_42_ctrl_serveStealReq_valid,
	io_connSS_42_ctrl_serveStealReq_ready,
	io_connSS_42_ctrl_stealReq_valid,
	io_connSS_42_ctrl_stealReq_ready,
	io_connSS_42_data_availableTask_ready,
	io_connSS_42_data_availableTask_valid,
	io_connSS_42_data_availableTask_bits,
	io_connSS_42_data_qOutTask_ready,
	io_connSS_42_data_qOutTask_valid,
	io_connSS_42_data_qOutTask_bits,
	io_connSS_43_ctrl_serveStealReq_valid,
	io_connSS_43_ctrl_serveStealReq_ready,
	io_connSS_43_ctrl_stealReq_valid,
	io_connSS_43_ctrl_stealReq_ready,
	io_connSS_43_data_availableTask_ready,
	io_connSS_43_data_availableTask_valid,
	io_connSS_43_data_availableTask_bits,
	io_connSS_43_data_qOutTask_ready,
	io_connSS_43_data_qOutTask_valid,
	io_connSS_43_data_qOutTask_bits,
	io_connSS_44_ctrl_serveStealReq_valid,
	io_connSS_44_ctrl_serveStealReq_ready,
	io_connSS_44_ctrl_stealReq_valid,
	io_connSS_44_ctrl_stealReq_ready,
	io_connSS_44_data_availableTask_ready,
	io_connSS_44_data_availableTask_valid,
	io_connSS_44_data_availableTask_bits,
	io_connSS_44_data_qOutTask_ready,
	io_connSS_44_data_qOutTask_valid,
	io_connSS_44_data_qOutTask_bits,
	io_connSS_45_ctrl_serveStealReq_valid,
	io_connSS_45_ctrl_serveStealReq_ready,
	io_connSS_45_ctrl_stealReq_valid,
	io_connSS_45_ctrl_stealReq_ready,
	io_connSS_45_data_availableTask_ready,
	io_connSS_45_data_availableTask_valid,
	io_connSS_45_data_availableTask_bits,
	io_connSS_45_data_qOutTask_ready,
	io_connSS_45_data_qOutTask_valid,
	io_connSS_45_data_qOutTask_bits,
	io_connSS_46_ctrl_serveStealReq_valid,
	io_connSS_46_ctrl_serveStealReq_ready,
	io_connSS_46_ctrl_stealReq_valid,
	io_connSS_46_ctrl_stealReq_ready,
	io_connSS_46_data_availableTask_ready,
	io_connSS_46_data_availableTask_valid,
	io_connSS_46_data_availableTask_bits,
	io_connSS_46_data_qOutTask_ready,
	io_connSS_46_data_qOutTask_valid,
	io_connSS_46_data_qOutTask_bits,
	io_connSS_47_ctrl_serveStealReq_valid,
	io_connSS_47_ctrl_serveStealReq_ready,
	io_connSS_47_ctrl_stealReq_valid,
	io_connSS_47_ctrl_stealReq_ready,
	io_connSS_47_data_availableTask_ready,
	io_connSS_47_data_availableTask_valid,
	io_connSS_47_data_availableTask_bits,
	io_connSS_47_data_qOutTask_ready,
	io_connSS_47_data_qOutTask_valid,
	io_connSS_47_data_qOutTask_bits,
	io_connSS_48_ctrl_serveStealReq_valid,
	io_connSS_48_ctrl_serveStealReq_ready,
	io_connSS_48_ctrl_stealReq_valid,
	io_connSS_48_ctrl_stealReq_ready,
	io_connSS_48_data_availableTask_ready,
	io_connSS_48_data_availableTask_valid,
	io_connSS_48_data_availableTask_bits,
	io_connSS_48_data_qOutTask_ready,
	io_connSS_48_data_qOutTask_valid,
	io_connSS_48_data_qOutTask_bits,
	io_connSS_49_ctrl_serveStealReq_valid,
	io_connSS_49_ctrl_serveStealReq_ready,
	io_connSS_49_ctrl_stealReq_valid,
	io_connSS_49_ctrl_stealReq_ready,
	io_connSS_49_data_availableTask_ready,
	io_connSS_49_data_availableTask_valid,
	io_connSS_49_data_availableTask_bits,
	io_connSS_49_data_qOutTask_ready,
	io_connSS_49_data_qOutTask_valid,
	io_connSS_49_data_qOutTask_bits,
	io_connSS_50_ctrl_serveStealReq_valid,
	io_connSS_50_ctrl_serveStealReq_ready,
	io_connSS_50_ctrl_stealReq_valid,
	io_connSS_50_ctrl_stealReq_ready,
	io_connSS_50_data_availableTask_ready,
	io_connSS_50_data_availableTask_valid,
	io_connSS_50_data_availableTask_bits,
	io_connSS_50_data_qOutTask_ready,
	io_connSS_50_data_qOutTask_valid,
	io_connSS_50_data_qOutTask_bits,
	io_connSS_51_ctrl_serveStealReq_valid,
	io_connSS_51_ctrl_serveStealReq_ready,
	io_connSS_51_ctrl_stealReq_valid,
	io_connSS_51_ctrl_stealReq_ready,
	io_connSS_51_data_availableTask_ready,
	io_connSS_51_data_availableTask_valid,
	io_connSS_51_data_availableTask_bits,
	io_connSS_51_data_qOutTask_ready,
	io_connSS_51_data_qOutTask_valid,
	io_connSS_51_data_qOutTask_bits,
	io_connSS_52_ctrl_serveStealReq_valid,
	io_connSS_52_ctrl_serveStealReq_ready,
	io_connSS_52_ctrl_stealReq_valid,
	io_connSS_52_ctrl_stealReq_ready,
	io_connSS_52_data_availableTask_ready,
	io_connSS_52_data_availableTask_valid,
	io_connSS_52_data_availableTask_bits,
	io_connSS_52_data_qOutTask_ready,
	io_connSS_52_data_qOutTask_valid,
	io_connSS_52_data_qOutTask_bits,
	io_connSS_53_ctrl_serveStealReq_valid,
	io_connSS_53_ctrl_serveStealReq_ready,
	io_connSS_53_ctrl_stealReq_valid,
	io_connSS_53_ctrl_stealReq_ready,
	io_connSS_53_data_availableTask_ready,
	io_connSS_53_data_availableTask_valid,
	io_connSS_53_data_availableTask_bits,
	io_connSS_53_data_qOutTask_ready,
	io_connSS_53_data_qOutTask_valid,
	io_connSS_53_data_qOutTask_bits,
	io_connSS_54_ctrl_serveStealReq_valid,
	io_connSS_54_ctrl_serveStealReq_ready,
	io_connSS_54_ctrl_stealReq_valid,
	io_connSS_54_ctrl_stealReq_ready,
	io_connSS_54_data_availableTask_ready,
	io_connSS_54_data_availableTask_valid,
	io_connSS_54_data_availableTask_bits,
	io_connSS_54_data_qOutTask_ready,
	io_connSS_54_data_qOutTask_valid,
	io_connSS_54_data_qOutTask_bits,
	io_connSS_55_ctrl_serveStealReq_valid,
	io_connSS_55_ctrl_serveStealReq_ready,
	io_connSS_55_ctrl_stealReq_valid,
	io_connSS_55_ctrl_stealReq_ready,
	io_connSS_55_data_availableTask_ready,
	io_connSS_55_data_availableTask_valid,
	io_connSS_55_data_availableTask_bits,
	io_connSS_55_data_qOutTask_ready,
	io_connSS_55_data_qOutTask_valid,
	io_connSS_55_data_qOutTask_bits,
	io_connSS_56_ctrl_serveStealReq_valid,
	io_connSS_56_ctrl_serveStealReq_ready,
	io_connSS_56_ctrl_stealReq_valid,
	io_connSS_56_ctrl_stealReq_ready,
	io_connSS_56_data_availableTask_ready,
	io_connSS_56_data_availableTask_valid,
	io_connSS_56_data_availableTask_bits,
	io_connSS_56_data_qOutTask_ready,
	io_connSS_56_data_qOutTask_valid,
	io_connSS_56_data_qOutTask_bits,
	io_connSS_57_ctrl_serveStealReq_valid,
	io_connSS_57_ctrl_serveStealReq_ready,
	io_connSS_57_ctrl_stealReq_valid,
	io_connSS_57_ctrl_stealReq_ready,
	io_connSS_57_data_availableTask_ready,
	io_connSS_57_data_availableTask_valid,
	io_connSS_57_data_availableTask_bits,
	io_connSS_57_data_qOutTask_ready,
	io_connSS_57_data_qOutTask_valid,
	io_connSS_57_data_qOutTask_bits,
	io_connSS_58_ctrl_serveStealReq_valid,
	io_connSS_58_ctrl_serveStealReq_ready,
	io_connSS_58_ctrl_stealReq_valid,
	io_connSS_58_ctrl_stealReq_ready,
	io_connSS_58_data_availableTask_ready,
	io_connSS_58_data_availableTask_valid,
	io_connSS_58_data_availableTask_bits,
	io_connSS_58_data_qOutTask_ready,
	io_connSS_58_data_qOutTask_valid,
	io_connSS_58_data_qOutTask_bits,
	io_connSS_59_ctrl_serveStealReq_valid,
	io_connSS_59_ctrl_serveStealReq_ready,
	io_connSS_59_ctrl_stealReq_valid,
	io_connSS_59_ctrl_stealReq_ready,
	io_connSS_59_data_availableTask_ready,
	io_connSS_59_data_availableTask_valid,
	io_connSS_59_data_availableTask_bits,
	io_connSS_59_data_qOutTask_ready,
	io_connSS_59_data_qOutTask_valid,
	io_connSS_59_data_qOutTask_bits,
	io_connSS_60_ctrl_serveStealReq_valid,
	io_connSS_60_ctrl_serveStealReq_ready,
	io_connSS_60_ctrl_stealReq_valid,
	io_connSS_60_ctrl_stealReq_ready,
	io_connSS_60_data_availableTask_ready,
	io_connSS_60_data_availableTask_valid,
	io_connSS_60_data_availableTask_bits,
	io_connSS_60_data_qOutTask_ready,
	io_connSS_60_data_qOutTask_valid,
	io_connSS_60_data_qOutTask_bits,
	io_connSS_61_ctrl_serveStealReq_valid,
	io_connSS_61_ctrl_serveStealReq_ready,
	io_connSS_61_ctrl_stealReq_valid,
	io_connSS_61_ctrl_stealReq_ready,
	io_connSS_61_data_availableTask_ready,
	io_connSS_61_data_availableTask_valid,
	io_connSS_61_data_availableTask_bits,
	io_connSS_61_data_qOutTask_ready,
	io_connSS_61_data_qOutTask_valid,
	io_connSS_61_data_qOutTask_bits,
	io_connSS_62_ctrl_serveStealReq_valid,
	io_connSS_62_ctrl_serveStealReq_ready,
	io_connSS_62_ctrl_stealReq_valid,
	io_connSS_62_ctrl_stealReq_ready,
	io_connSS_62_data_availableTask_ready,
	io_connSS_62_data_availableTask_valid,
	io_connSS_62_data_availableTask_bits,
	io_connSS_62_data_qOutTask_ready,
	io_connSS_62_data_qOutTask_valid,
	io_connSS_62_data_qOutTask_bits,
	io_connSS_63_ctrl_serveStealReq_valid,
	io_connSS_63_ctrl_serveStealReq_ready,
	io_connSS_63_ctrl_stealReq_valid,
	io_connSS_63_ctrl_stealReq_ready,
	io_connSS_63_data_availableTask_ready,
	io_connSS_63_data_availableTask_valid,
	io_connSS_63_data_availableTask_bits,
	io_connSS_63_data_qOutTask_ready,
	io_connSS_63_data_qOutTask_valid,
	io_connSS_63_data_qOutTask_bits,
	io_connSS_64_ctrl_serveStealReq_valid,
	io_connSS_64_ctrl_serveStealReq_ready,
	io_connSS_64_ctrl_stealReq_valid,
	io_connSS_64_ctrl_stealReq_ready,
	io_connSS_64_data_availableTask_ready,
	io_connSS_64_data_availableTask_valid,
	io_connSS_64_data_availableTask_bits,
	io_connSS_64_data_qOutTask_ready,
	io_connSS_64_data_qOutTask_valid,
	io_connSS_64_data_qOutTask_bits,
	io_connSS_65_ctrl_serveStealReq_valid,
	io_connSS_65_ctrl_serveStealReq_ready,
	io_connSS_65_ctrl_stealReq_valid,
	io_connSS_65_ctrl_stealReq_ready,
	io_connSS_65_data_availableTask_ready,
	io_connSS_65_data_availableTask_valid,
	io_connSS_65_data_availableTask_bits,
	io_connSS_65_data_qOutTask_ready,
	io_connSS_65_data_qOutTask_valid,
	io_connSS_65_data_qOutTask_bits,
	io_connSS_66_ctrl_serveStealReq_valid,
	io_connSS_66_ctrl_serveStealReq_ready,
	io_connSS_66_ctrl_stealReq_valid,
	io_connSS_66_ctrl_stealReq_ready,
	io_connSS_66_data_availableTask_ready,
	io_connSS_66_data_availableTask_valid,
	io_connSS_66_data_availableTask_bits,
	io_connSS_66_data_qOutTask_ready,
	io_connSS_66_data_qOutTask_valid,
	io_connSS_66_data_qOutTask_bits,
	io_connSS_67_ctrl_serveStealReq_valid,
	io_connSS_67_ctrl_serveStealReq_ready,
	io_connSS_67_ctrl_stealReq_valid,
	io_connSS_67_ctrl_stealReq_ready,
	io_connSS_67_data_availableTask_ready,
	io_connSS_67_data_availableTask_valid,
	io_connSS_67_data_availableTask_bits,
	io_connSS_67_data_qOutTask_ready,
	io_connSS_67_data_qOutTask_valid,
	io_connSS_67_data_qOutTask_bits,
	io_connSS_68_ctrl_serveStealReq_valid,
	io_connSS_68_ctrl_serveStealReq_ready,
	io_connSS_68_ctrl_stealReq_valid,
	io_connSS_68_ctrl_stealReq_ready,
	io_connSS_68_data_availableTask_ready,
	io_connSS_68_data_availableTask_valid,
	io_connSS_68_data_availableTask_bits,
	io_connSS_68_data_qOutTask_ready,
	io_connSS_68_data_qOutTask_valid,
	io_connSS_68_data_qOutTask_bits,
	io_connSS_69_ctrl_serveStealReq_valid,
	io_connSS_69_ctrl_serveStealReq_ready,
	io_connSS_69_ctrl_stealReq_valid,
	io_connSS_69_ctrl_stealReq_ready,
	io_connSS_69_data_availableTask_ready,
	io_connSS_69_data_availableTask_valid,
	io_connSS_69_data_availableTask_bits,
	io_connSS_69_data_qOutTask_ready,
	io_connSS_69_data_qOutTask_valid,
	io_connSS_69_data_qOutTask_bits,
	io_connSS_70_ctrl_serveStealReq_valid,
	io_connSS_70_ctrl_serveStealReq_ready,
	io_connSS_70_ctrl_stealReq_valid,
	io_connSS_70_ctrl_stealReq_ready,
	io_connSS_70_data_availableTask_ready,
	io_connSS_70_data_availableTask_valid,
	io_connSS_70_data_availableTask_bits,
	io_connSS_70_data_qOutTask_ready,
	io_connSS_70_data_qOutTask_valid,
	io_connSS_70_data_qOutTask_bits,
	io_connSS_71_ctrl_serveStealReq_valid,
	io_connSS_71_ctrl_serveStealReq_ready,
	io_connSS_71_ctrl_stealReq_valid,
	io_connSS_71_ctrl_stealReq_ready,
	io_connSS_71_data_availableTask_ready,
	io_connSS_71_data_availableTask_valid,
	io_connSS_71_data_availableTask_bits,
	io_connSS_71_data_qOutTask_ready,
	io_connSS_71_data_qOutTask_valid,
	io_connSS_71_data_qOutTask_bits,
	io_connSS_72_ctrl_serveStealReq_valid,
	io_connSS_72_ctrl_serveStealReq_ready,
	io_connSS_72_ctrl_stealReq_valid,
	io_connSS_72_ctrl_stealReq_ready,
	io_connSS_72_data_availableTask_ready,
	io_connSS_72_data_availableTask_valid,
	io_connSS_72_data_availableTask_bits,
	io_connSS_72_data_qOutTask_ready,
	io_connSS_72_data_qOutTask_valid,
	io_connSS_72_data_qOutTask_bits,
	io_connSS_73_ctrl_serveStealReq_valid,
	io_connSS_73_ctrl_serveStealReq_ready,
	io_connSS_73_ctrl_stealReq_valid,
	io_connSS_73_ctrl_stealReq_ready,
	io_connSS_73_data_availableTask_ready,
	io_connSS_73_data_availableTask_valid,
	io_connSS_73_data_availableTask_bits,
	io_connSS_73_data_qOutTask_ready,
	io_connSS_73_data_qOutTask_valid,
	io_connSS_73_data_qOutTask_bits,
	io_connSS_74_ctrl_serveStealReq_valid,
	io_connSS_74_ctrl_serveStealReq_ready,
	io_connSS_74_ctrl_stealReq_valid,
	io_connSS_74_ctrl_stealReq_ready,
	io_connSS_74_data_availableTask_ready,
	io_connSS_74_data_availableTask_valid,
	io_connSS_74_data_availableTask_bits,
	io_connSS_74_data_qOutTask_ready,
	io_connSS_74_data_qOutTask_valid,
	io_connSS_74_data_qOutTask_bits,
	io_connSS_75_ctrl_serveStealReq_valid,
	io_connSS_75_ctrl_serveStealReq_ready,
	io_connSS_75_ctrl_stealReq_valid,
	io_connSS_75_ctrl_stealReq_ready,
	io_connSS_75_data_availableTask_ready,
	io_connSS_75_data_availableTask_valid,
	io_connSS_75_data_availableTask_bits,
	io_connSS_75_data_qOutTask_ready,
	io_connSS_75_data_qOutTask_valid,
	io_connSS_75_data_qOutTask_bits,
	io_connSS_76_ctrl_serveStealReq_valid,
	io_connSS_76_ctrl_serveStealReq_ready,
	io_connSS_76_ctrl_stealReq_valid,
	io_connSS_76_ctrl_stealReq_ready,
	io_connSS_76_data_availableTask_ready,
	io_connSS_76_data_availableTask_valid,
	io_connSS_76_data_availableTask_bits,
	io_connSS_76_data_qOutTask_ready,
	io_connSS_76_data_qOutTask_valid,
	io_connSS_76_data_qOutTask_bits,
	io_connSS_77_ctrl_serveStealReq_valid,
	io_connSS_77_ctrl_serveStealReq_ready,
	io_connSS_77_ctrl_stealReq_valid,
	io_connSS_77_ctrl_stealReq_ready,
	io_connSS_77_data_availableTask_ready,
	io_connSS_77_data_availableTask_valid,
	io_connSS_77_data_availableTask_bits,
	io_connSS_77_data_qOutTask_ready,
	io_connSS_77_data_qOutTask_valid,
	io_connSS_77_data_qOutTask_bits,
	io_connSS_78_ctrl_serveStealReq_valid,
	io_connSS_78_ctrl_serveStealReq_ready,
	io_connSS_78_ctrl_stealReq_valid,
	io_connSS_78_ctrl_stealReq_ready,
	io_connSS_78_data_availableTask_ready,
	io_connSS_78_data_availableTask_valid,
	io_connSS_78_data_availableTask_bits,
	io_connSS_78_data_qOutTask_ready,
	io_connSS_78_data_qOutTask_valid,
	io_connSS_78_data_qOutTask_bits,
	io_connSS_79_ctrl_serveStealReq_valid,
	io_connSS_79_ctrl_serveStealReq_ready,
	io_connSS_79_ctrl_stealReq_valid,
	io_connSS_79_ctrl_stealReq_ready,
	io_connSS_79_data_availableTask_ready,
	io_connSS_79_data_availableTask_valid,
	io_connSS_79_data_availableTask_bits,
	io_connSS_79_data_qOutTask_ready,
	io_connSS_79_data_qOutTask_valid,
	io_connSS_79_data_qOutTask_bits,
	io_connSS_80_ctrl_serveStealReq_valid,
	io_connSS_80_ctrl_serveStealReq_ready,
	io_connSS_80_ctrl_stealReq_valid,
	io_connSS_80_ctrl_stealReq_ready,
	io_connSS_80_data_availableTask_ready,
	io_connSS_80_data_availableTask_valid,
	io_connSS_80_data_availableTask_bits,
	io_connSS_80_data_qOutTask_ready,
	io_connSS_80_data_qOutTask_valid,
	io_connSS_80_data_qOutTask_bits,
	io_connSS_81_ctrl_serveStealReq_valid,
	io_connSS_81_ctrl_serveStealReq_ready,
	io_connSS_81_ctrl_stealReq_valid,
	io_connSS_81_ctrl_stealReq_ready,
	io_connSS_81_data_availableTask_ready,
	io_connSS_81_data_availableTask_valid,
	io_connSS_81_data_availableTask_bits,
	io_connSS_81_data_qOutTask_ready,
	io_connSS_81_data_qOutTask_valid,
	io_connSS_81_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0,
	io_ntwDataUnitOccupancyVSS_1
);
	input clock;
	input reset;
	input io_connSS_0_ctrl_serveStealReq_valid;
	output wire io_connSS_0_ctrl_serveStealReq_ready;
	input io_connSS_0_data_availableTask_ready;
	output wire io_connSS_0_data_availableTask_valid;
	output wire [255:0] io_connSS_0_data_availableTask_bits;
	output wire io_connSS_0_data_qOutTask_ready;
	input io_connSS_0_data_qOutTask_valid;
	input [255:0] io_connSS_0_data_qOutTask_bits;
	input io_connSS_1_ctrl_serveStealReq_valid;
	output wire io_connSS_1_ctrl_serveStealReq_ready;
	input io_connSS_1_data_availableTask_ready;
	output wire io_connSS_1_data_availableTask_valid;
	output wire [255:0] io_connSS_1_data_availableTask_bits;
	output wire io_connSS_1_data_qOutTask_ready;
	input io_connSS_1_data_qOutTask_valid;
	input [255:0] io_connSS_1_data_qOutTask_bits;
	input io_connSS_2_ctrl_serveStealReq_valid;
	output wire io_connSS_2_ctrl_serveStealReq_ready;
	output wire io_connSS_2_data_qOutTask_ready;
	input io_connSS_2_data_qOutTask_valid;
	input [255:0] io_connSS_2_data_qOutTask_bits;
	input io_connSS_3_ctrl_serveStealReq_valid;
	output wire io_connSS_3_ctrl_serveStealReq_ready;
	output wire io_connSS_3_data_qOutTask_ready;
	input io_connSS_3_data_qOutTask_valid;
	input [255:0] io_connSS_3_data_qOutTask_bits;
	input io_connSS_4_ctrl_serveStealReq_valid;
	output wire io_connSS_4_ctrl_serveStealReq_ready;
	output wire io_connSS_4_data_qOutTask_ready;
	input io_connSS_4_data_qOutTask_valid;
	input [255:0] io_connSS_4_data_qOutTask_bits;
	input io_connSS_5_ctrl_serveStealReq_valid;
	output wire io_connSS_5_ctrl_serveStealReq_ready;
	output wire io_connSS_5_data_qOutTask_ready;
	input io_connSS_5_data_qOutTask_valid;
	input [255:0] io_connSS_5_data_qOutTask_bits;
	input io_connSS_6_ctrl_serveStealReq_valid;
	output wire io_connSS_6_ctrl_serveStealReq_ready;
	output wire io_connSS_6_data_qOutTask_ready;
	input io_connSS_6_data_qOutTask_valid;
	input [255:0] io_connSS_6_data_qOutTask_bits;
	input io_connSS_7_ctrl_serveStealReq_valid;
	output wire io_connSS_7_ctrl_serveStealReq_ready;
	output wire io_connSS_7_data_qOutTask_ready;
	input io_connSS_7_data_qOutTask_valid;
	input [255:0] io_connSS_7_data_qOutTask_bits;
	input io_connSS_8_ctrl_serveStealReq_valid;
	output wire io_connSS_8_ctrl_serveStealReq_ready;
	output wire io_connSS_8_data_qOutTask_ready;
	input io_connSS_8_data_qOutTask_valid;
	input [255:0] io_connSS_8_data_qOutTask_bits;
	input io_connSS_9_ctrl_serveStealReq_valid;
	output wire io_connSS_9_ctrl_serveStealReq_ready;
	output wire io_connSS_9_data_qOutTask_ready;
	input io_connSS_9_data_qOutTask_valid;
	input [255:0] io_connSS_9_data_qOutTask_bits;
	input io_connSS_10_ctrl_serveStealReq_valid;
	output wire io_connSS_10_ctrl_serveStealReq_ready;
	output wire io_connSS_10_data_qOutTask_ready;
	input io_connSS_10_data_qOutTask_valid;
	input [255:0] io_connSS_10_data_qOutTask_bits;
	input io_connSS_11_ctrl_serveStealReq_valid;
	output wire io_connSS_11_ctrl_serveStealReq_ready;
	output wire io_connSS_11_data_qOutTask_ready;
	input io_connSS_11_data_qOutTask_valid;
	input [255:0] io_connSS_11_data_qOutTask_bits;
	input io_connSS_12_ctrl_serveStealReq_valid;
	output wire io_connSS_12_ctrl_serveStealReq_ready;
	output wire io_connSS_12_data_qOutTask_ready;
	input io_connSS_12_data_qOutTask_valid;
	input [255:0] io_connSS_12_data_qOutTask_bits;
	input io_connSS_13_ctrl_serveStealReq_valid;
	output wire io_connSS_13_ctrl_serveStealReq_ready;
	output wire io_connSS_13_data_qOutTask_ready;
	input io_connSS_13_data_qOutTask_valid;
	input [255:0] io_connSS_13_data_qOutTask_bits;
	input io_connSS_14_ctrl_serveStealReq_valid;
	output wire io_connSS_14_ctrl_serveStealReq_ready;
	output wire io_connSS_14_data_qOutTask_ready;
	input io_connSS_14_data_qOutTask_valid;
	input [255:0] io_connSS_14_data_qOutTask_bits;
	input io_connSS_15_ctrl_serveStealReq_valid;
	output wire io_connSS_15_ctrl_serveStealReq_ready;
	output wire io_connSS_15_data_qOutTask_ready;
	input io_connSS_15_data_qOutTask_valid;
	input [255:0] io_connSS_15_data_qOutTask_bits;
	input io_connSS_16_ctrl_serveStealReq_valid;
	output wire io_connSS_16_ctrl_serveStealReq_ready;
	output wire io_connSS_16_data_qOutTask_ready;
	input io_connSS_16_data_qOutTask_valid;
	input [255:0] io_connSS_16_data_qOutTask_bits;
	input io_connSS_17_ctrl_serveStealReq_valid;
	output wire io_connSS_17_ctrl_serveStealReq_ready;
	output wire io_connSS_17_data_qOutTask_ready;
	input io_connSS_17_data_qOutTask_valid;
	input [255:0] io_connSS_17_data_qOutTask_bits;
	input io_connSS_18_ctrl_serveStealReq_valid;
	output wire io_connSS_18_ctrl_serveStealReq_ready;
	input io_connSS_18_ctrl_stealReq_valid;
	output wire io_connSS_18_ctrl_stealReq_ready;
	input io_connSS_18_data_availableTask_ready;
	output wire io_connSS_18_data_availableTask_valid;
	output wire [255:0] io_connSS_18_data_availableTask_bits;
	output wire io_connSS_18_data_qOutTask_ready;
	input io_connSS_18_data_qOutTask_valid;
	input [255:0] io_connSS_18_data_qOutTask_bits;
	input io_connSS_19_ctrl_serveStealReq_valid;
	output wire io_connSS_19_ctrl_serveStealReq_ready;
	input io_connSS_19_ctrl_stealReq_valid;
	output wire io_connSS_19_ctrl_stealReq_ready;
	input io_connSS_19_data_availableTask_ready;
	output wire io_connSS_19_data_availableTask_valid;
	output wire [255:0] io_connSS_19_data_availableTask_bits;
	output wire io_connSS_19_data_qOutTask_ready;
	input io_connSS_19_data_qOutTask_valid;
	input [255:0] io_connSS_19_data_qOutTask_bits;
	input io_connSS_20_ctrl_serveStealReq_valid;
	output wire io_connSS_20_ctrl_serveStealReq_ready;
	input io_connSS_20_ctrl_stealReq_valid;
	output wire io_connSS_20_ctrl_stealReq_ready;
	input io_connSS_20_data_availableTask_ready;
	output wire io_connSS_20_data_availableTask_valid;
	output wire [255:0] io_connSS_20_data_availableTask_bits;
	output wire io_connSS_20_data_qOutTask_ready;
	input io_connSS_20_data_qOutTask_valid;
	input [255:0] io_connSS_20_data_qOutTask_bits;
	input io_connSS_21_ctrl_serveStealReq_valid;
	output wire io_connSS_21_ctrl_serveStealReq_ready;
	input io_connSS_21_ctrl_stealReq_valid;
	output wire io_connSS_21_ctrl_stealReq_ready;
	input io_connSS_21_data_availableTask_ready;
	output wire io_connSS_21_data_availableTask_valid;
	output wire [255:0] io_connSS_21_data_availableTask_bits;
	output wire io_connSS_21_data_qOutTask_ready;
	input io_connSS_21_data_qOutTask_valid;
	input [255:0] io_connSS_21_data_qOutTask_bits;
	input io_connSS_22_ctrl_serveStealReq_valid;
	output wire io_connSS_22_ctrl_serveStealReq_ready;
	input io_connSS_22_ctrl_stealReq_valid;
	output wire io_connSS_22_ctrl_stealReq_ready;
	input io_connSS_22_data_availableTask_ready;
	output wire io_connSS_22_data_availableTask_valid;
	output wire [255:0] io_connSS_22_data_availableTask_bits;
	output wire io_connSS_22_data_qOutTask_ready;
	input io_connSS_22_data_qOutTask_valid;
	input [255:0] io_connSS_22_data_qOutTask_bits;
	input io_connSS_23_ctrl_serveStealReq_valid;
	output wire io_connSS_23_ctrl_serveStealReq_ready;
	input io_connSS_23_ctrl_stealReq_valid;
	output wire io_connSS_23_ctrl_stealReq_ready;
	input io_connSS_23_data_availableTask_ready;
	output wire io_connSS_23_data_availableTask_valid;
	output wire [255:0] io_connSS_23_data_availableTask_bits;
	output wire io_connSS_23_data_qOutTask_ready;
	input io_connSS_23_data_qOutTask_valid;
	input [255:0] io_connSS_23_data_qOutTask_bits;
	input io_connSS_24_ctrl_serveStealReq_valid;
	output wire io_connSS_24_ctrl_serveStealReq_ready;
	input io_connSS_24_ctrl_stealReq_valid;
	output wire io_connSS_24_ctrl_stealReq_ready;
	input io_connSS_24_data_availableTask_ready;
	output wire io_connSS_24_data_availableTask_valid;
	output wire [255:0] io_connSS_24_data_availableTask_bits;
	output wire io_connSS_24_data_qOutTask_ready;
	input io_connSS_24_data_qOutTask_valid;
	input [255:0] io_connSS_24_data_qOutTask_bits;
	input io_connSS_25_ctrl_serveStealReq_valid;
	output wire io_connSS_25_ctrl_serveStealReq_ready;
	input io_connSS_25_ctrl_stealReq_valid;
	output wire io_connSS_25_ctrl_stealReq_ready;
	input io_connSS_25_data_availableTask_ready;
	output wire io_connSS_25_data_availableTask_valid;
	output wire [255:0] io_connSS_25_data_availableTask_bits;
	output wire io_connSS_25_data_qOutTask_ready;
	input io_connSS_25_data_qOutTask_valid;
	input [255:0] io_connSS_25_data_qOutTask_bits;
	input io_connSS_26_ctrl_serveStealReq_valid;
	output wire io_connSS_26_ctrl_serveStealReq_ready;
	input io_connSS_26_ctrl_stealReq_valid;
	output wire io_connSS_26_ctrl_stealReq_ready;
	input io_connSS_26_data_availableTask_ready;
	output wire io_connSS_26_data_availableTask_valid;
	output wire [255:0] io_connSS_26_data_availableTask_bits;
	output wire io_connSS_26_data_qOutTask_ready;
	input io_connSS_26_data_qOutTask_valid;
	input [255:0] io_connSS_26_data_qOutTask_bits;
	input io_connSS_27_ctrl_serveStealReq_valid;
	output wire io_connSS_27_ctrl_serveStealReq_ready;
	input io_connSS_27_ctrl_stealReq_valid;
	output wire io_connSS_27_ctrl_stealReq_ready;
	input io_connSS_27_data_availableTask_ready;
	output wire io_connSS_27_data_availableTask_valid;
	output wire [255:0] io_connSS_27_data_availableTask_bits;
	output wire io_connSS_27_data_qOutTask_ready;
	input io_connSS_27_data_qOutTask_valid;
	input [255:0] io_connSS_27_data_qOutTask_bits;
	input io_connSS_28_ctrl_serveStealReq_valid;
	output wire io_connSS_28_ctrl_serveStealReq_ready;
	input io_connSS_28_ctrl_stealReq_valid;
	output wire io_connSS_28_ctrl_stealReq_ready;
	input io_connSS_28_data_availableTask_ready;
	output wire io_connSS_28_data_availableTask_valid;
	output wire [255:0] io_connSS_28_data_availableTask_bits;
	output wire io_connSS_28_data_qOutTask_ready;
	input io_connSS_28_data_qOutTask_valid;
	input [255:0] io_connSS_28_data_qOutTask_bits;
	input io_connSS_29_ctrl_serveStealReq_valid;
	output wire io_connSS_29_ctrl_serveStealReq_ready;
	input io_connSS_29_ctrl_stealReq_valid;
	output wire io_connSS_29_ctrl_stealReq_ready;
	input io_connSS_29_data_availableTask_ready;
	output wire io_connSS_29_data_availableTask_valid;
	output wire [255:0] io_connSS_29_data_availableTask_bits;
	output wire io_connSS_29_data_qOutTask_ready;
	input io_connSS_29_data_qOutTask_valid;
	input [255:0] io_connSS_29_data_qOutTask_bits;
	input io_connSS_30_ctrl_serveStealReq_valid;
	output wire io_connSS_30_ctrl_serveStealReq_ready;
	input io_connSS_30_ctrl_stealReq_valid;
	output wire io_connSS_30_ctrl_stealReq_ready;
	input io_connSS_30_data_availableTask_ready;
	output wire io_connSS_30_data_availableTask_valid;
	output wire [255:0] io_connSS_30_data_availableTask_bits;
	output wire io_connSS_30_data_qOutTask_ready;
	input io_connSS_30_data_qOutTask_valid;
	input [255:0] io_connSS_30_data_qOutTask_bits;
	input io_connSS_31_ctrl_serveStealReq_valid;
	output wire io_connSS_31_ctrl_serveStealReq_ready;
	input io_connSS_31_ctrl_stealReq_valid;
	output wire io_connSS_31_ctrl_stealReq_ready;
	input io_connSS_31_data_availableTask_ready;
	output wire io_connSS_31_data_availableTask_valid;
	output wire [255:0] io_connSS_31_data_availableTask_bits;
	output wire io_connSS_31_data_qOutTask_ready;
	input io_connSS_31_data_qOutTask_valid;
	input [255:0] io_connSS_31_data_qOutTask_bits;
	input io_connSS_32_ctrl_serveStealReq_valid;
	output wire io_connSS_32_ctrl_serveStealReq_ready;
	input io_connSS_32_ctrl_stealReq_valid;
	output wire io_connSS_32_ctrl_stealReq_ready;
	input io_connSS_32_data_availableTask_ready;
	output wire io_connSS_32_data_availableTask_valid;
	output wire [255:0] io_connSS_32_data_availableTask_bits;
	output wire io_connSS_32_data_qOutTask_ready;
	input io_connSS_32_data_qOutTask_valid;
	input [255:0] io_connSS_32_data_qOutTask_bits;
	input io_connSS_33_ctrl_serveStealReq_valid;
	output wire io_connSS_33_ctrl_serveStealReq_ready;
	input io_connSS_33_ctrl_stealReq_valid;
	output wire io_connSS_33_ctrl_stealReq_ready;
	input io_connSS_33_data_availableTask_ready;
	output wire io_connSS_33_data_availableTask_valid;
	output wire [255:0] io_connSS_33_data_availableTask_bits;
	output wire io_connSS_33_data_qOutTask_ready;
	input io_connSS_33_data_qOutTask_valid;
	input [255:0] io_connSS_33_data_qOutTask_bits;
	input io_connSS_34_ctrl_serveStealReq_valid;
	output wire io_connSS_34_ctrl_serveStealReq_ready;
	input io_connSS_34_ctrl_stealReq_valid;
	output wire io_connSS_34_ctrl_stealReq_ready;
	input io_connSS_34_data_availableTask_ready;
	output wire io_connSS_34_data_availableTask_valid;
	output wire [255:0] io_connSS_34_data_availableTask_bits;
	output wire io_connSS_34_data_qOutTask_ready;
	input io_connSS_34_data_qOutTask_valid;
	input [255:0] io_connSS_34_data_qOutTask_bits;
	input io_connSS_35_ctrl_serveStealReq_valid;
	output wire io_connSS_35_ctrl_serveStealReq_ready;
	input io_connSS_35_ctrl_stealReq_valid;
	output wire io_connSS_35_ctrl_stealReq_ready;
	input io_connSS_35_data_availableTask_ready;
	output wire io_connSS_35_data_availableTask_valid;
	output wire [255:0] io_connSS_35_data_availableTask_bits;
	output wire io_connSS_35_data_qOutTask_ready;
	input io_connSS_35_data_qOutTask_valid;
	input [255:0] io_connSS_35_data_qOutTask_bits;
	input io_connSS_36_ctrl_serveStealReq_valid;
	output wire io_connSS_36_ctrl_serveStealReq_ready;
	input io_connSS_36_ctrl_stealReq_valid;
	output wire io_connSS_36_ctrl_stealReq_ready;
	input io_connSS_36_data_availableTask_ready;
	output wire io_connSS_36_data_availableTask_valid;
	output wire [255:0] io_connSS_36_data_availableTask_bits;
	output wire io_connSS_36_data_qOutTask_ready;
	input io_connSS_36_data_qOutTask_valid;
	input [255:0] io_connSS_36_data_qOutTask_bits;
	input io_connSS_37_ctrl_serveStealReq_valid;
	output wire io_connSS_37_ctrl_serveStealReq_ready;
	input io_connSS_37_ctrl_stealReq_valid;
	output wire io_connSS_37_ctrl_stealReq_ready;
	input io_connSS_37_data_availableTask_ready;
	output wire io_connSS_37_data_availableTask_valid;
	output wire [255:0] io_connSS_37_data_availableTask_bits;
	output wire io_connSS_37_data_qOutTask_ready;
	input io_connSS_37_data_qOutTask_valid;
	input [255:0] io_connSS_37_data_qOutTask_bits;
	input io_connSS_38_ctrl_serveStealReq_valid;
	output wire io_connSS_38_ctrl_serveStealReq_ready;
	input io_connSS_38_ctrl_stealReq_valid;
	output wire io_connSS_38_ctrl_stealReq_ready;
	input io_connSS_38_data_availableTask_ready;
	output wire io_connSS_38_data_availableTask_valid;
	output wire [255:0] io_connSS_38_data_availableTask_bits;
	output wire io_connSS_38_data_qOutTask_ready;
	input io_connSS_38_data_qOutTask_valid;
	input [255:0] io_connSS_38_data_qOutTask_bits;
	input io_connSS_39_ctrl_serveStealReq_valid;
	output wire io_connSS_39_ctrl_serveStealReq_ready;
	input io_connSS_39_ctrl_stealReq_valid;
	output wire io_connSS_39_ctrl_stealReq_ready;
	input io_connSS_39_data_availableTask_ready;
	output wire io_connSS_39_data_availableTask_valid;
	output wire [255:0] io_connSS_39_data_availableTask_bits;
	output wire io_connSS_39_data_qOutTask_ready;
	input io_connSS_39_data_qOutTask_valid;
	input [255:0] io_connSS_39_data_qOutTask_bits;
	input io_connSS_40_ctrl_serveStealReq_valid;
	output wire io_connSS_40_ctrl_serveStealReq_ready;
	input io_connSS_40_ctrl_stealReq_valid;
	output wire io_connSS_40_ctrl_stealReq_ready;
	input io_connSS_40_data_availableTask_ready;
	output wire io_connSS_40_data_availableTask_valid;
	output wire [255:0] io_connSS_40_data_availableTask_bits;
	output wire io_connSS_40_data_qOutTask_ready;
	input io_connSS_40_data_qOutTask_valid;
	input [255:0] io_connSS_40_data_qOutTask_bits;
	input io_connSS_41_ctrl_serveStealReq_valid;
	output wire io_connSS_41_ctrl_serveStealReq_ready;
	input io_connSS_41_ctrl_stealReq_valid;
	output wire io_connSS_41_ctrl_stealReq_ready;
	input io_connSS_41_data_availableTask_ready;
	output wire io_connSS_41_data_availableTask_valid;
	output wire [255:0] io_connSS_41_data_availableTask_bits;
	output wire io_connSS_41_data_qOutTask_ready;
	input io_connSS_41_data_qOutTask_valid;
	input [255:0] io_connSS_41_data_qOutTask_bits;
	input io_connSS_42_ctrl_serveStealReq_valid;
	output wire io_connSS_42_ctrl_serveStealReq_ready;
	input io_connSS_42_ctrl_stealReq_valid;
	output wire io_connSS_42_ctrl_stealReq_ready;
	input io_connSS_42_data_availableTask_ready;
	output wire io_connSS_42_data_availableTask_valid;
	output wire [255:0] io_connSS_42_data_availableTask_bits;
	output wire io_connSS_42_data_qOutTask_ready;
	input io_connSS_42_data_qOutTask_valid;
	input [255:0] io_connSS_42_data_qOutTask_bits;
	input io_connSS_43_ctrl_serveStealReq_valid;
	output wire io_connSS_43_ctrl_serveStealReq_ready;
	input io_connSS_43_ctrl_stealReq_valid;
	output wire io_connSS_43_ctrl_stealReq_ready;
	input io_connSS_43_data_availableTask_ready;
	output wire io_connSS_43_data_availableTask_valid;
	output wire [255:0] io_connSS_43_data_availableTask_bits;
	output wire io_connSS_43_data_qOutTask_ready;
	input io_connSS_43_data_qOutTask_valid;
	input [255:0] io_connSS_43_data_qOutTask_bits;
	input io_connSS_44_ctrl_serveStealReq_valid;
	output wire io_connSS_44_ctrl_serveStealReq_ready;
	input io_connSS_44_ctrl_stealReq_valid;
	output wire io_connSS_44_ctrl_stealReq_ready;
	input io_connSS_44_data_availableTask_ready;
	output wire io_connSS_44_data_availableTask_valid;
	output wire [255:0] io_connSS_44_data_availableTask_bits;
	output wire io_connSS_44_data_qOutTask_ready;
	input io_connSS_44_data_qOutTask_valid;
	input [255:0] io_connSS_44_data_qOutTask_bits;
	input io_connSS_45_ctrl_serveStealReq_valid;
	output wire io_connSS_45_ctrl_serveStealReq_ready;
	input io_connSS_45_ctrl_stealReq_valid;
	output wire io_connSS_45_ctrl_stealReq_ready;
	input io_connSS_45_data_availableTask_ready;
	output wire io_connSS_45_data_availableTask_valid;
	output wire [255:0] io_connSS_45_data_availableTask_bits;
	output wire io_connSS_45_data_qOutTask_ready;
	input io_connSS_45_data_qOutTask_valid;
	input [255:0] io_connSS_45_data_qOutTask_bits;
	input io_connSS_46_ctrl_serveStealReq_valid;
	output wire io_connSS_46_ctrl_serveStealReq_ready;
	input io_connSS_46_ctrl_stealReq_valid;
	output wire io_connSS_46_ctrl_stealReq_ready;
	input io_connSS_46_data_availableTask_ready;
	output wire io_connSS_46_data_availableTask_valid;
	output wire [255:0] io_connSS_46_data_availableTask_bits;
	output wire io_connSS_46_data_qOutTask_ready;
	input io_connSS_46_data_qOutTask_valid;
	input [255:0] io_connSS_46_data_qOutTask_bits;
	input io_connSS_47_ctrl_serveStealReq_valid;
	output wire io_connSS_47_ctrl_serveStealReq_ready;
	input io_connSS_47_ctrl_stealReq_valid;
	output wire io_connSS_47_ctrl_stealReq_ready;
	input io_connSS_47_data_availableTask_ready;
	output wire io_connSS_47_data_availableTask_valid;
	output wire [255:0] io_connSS_47_data_availableTask_bits;
	output wire io_connSS_47_data_qOutTask_ready;
	input io_connSS_47_data_qOutTask_valid;
	input [255:0] io_connSS_47_data_qOutTask_bits;
	input io_connSS_48_ctrl_serveStealReq_valid;
	output wire io_connSS_48_ctrl_serveStealReq_ready;
	input io_connSS_48_ctrl_stealReq_valid;
	output wire io_connSS_48_ctrl_stealReq_ready;
	input io_connSS_48_data_availableTask_ready;
	output wire io_connSS_48_data_availableTask_valid;
	output wire [255:0] io_connSS_48_data_availableTask_bits;
	output wire io_connSS_48_data_qOutTask_ready;
	input io_connSS_48_data_qOutTask_valid;
	input [255:0] io_connSS_48_data_qOutTask_bits;
	input io_connSS_49_ctrl_serveStealReq_valid;
	output wire io_connSS_49_ctrl_serveStealReq_ready;
	input io_connSS_49_ctrl_stealReq_valid;
	output wire io_connSS_49_ctrl_stealReq_ready;
	input io_connSS_49_data_availableTask_ready;
	output wire io_connSS_49_data_availableTask_valid;
	output wire [255:0] io_connSS_49_data_availableTask_bits;
	output wire io_connSS_49_data_qOutTask_ready;
	input io_connSS_49_data_qOutTask_valid;
	input [255:0] io_connSS_49_data_qOutTask_bits;
	input io_connSS_50_ctrl_serveStealReq_valid;
	output wire io_connSS_50_ctrl_serveStealReq_ready;
	input io_connSS_50_ctrl_stealReq_valid;
	output wire io_connSS_50_ctrl_stealReq_ready;
	input io_connSS_50_data_availableTask_ready;
	output wire io_connSS_50_data_availableTask_valid;
	output wire [255:0] io_connSS_50_data_availableTask_bits;
	output wire io_connSS_50_data_qOutTask_ready;
	input io_connSS_50_data_qOutTask_valid;
	input [255:0] io_connSS_50_data_qOutTask_bits;
	input io_connSS_51_ctrl_serveStealReq_valid;
	output wire io_connSS_51_ctrl_serveStealReq_ready;
	input io_connSS_51_ctrl_stealReq_valid;
	output wire io_connSS_51_ctrl_stealReq_ready;
	input io_connSS_51_data_availableTask_ready;
	output wire io_connSS_51_data_availableTask_valid;
	output wire [255:0] io_connSS_51_data_availableTask_bits;
	output wire io_connSS_51_data_qOutTask_ready;
	input io_connSS_51_data_qOutTask_valid;
	input [255:0] io_connSS_51_data_qOutTask_bits;
	input io_connSS_52_ctrl_serveStealReq_valid;
	output wire io_connSS_52_ctrl_serveStealReq_ready;
	input io_connSS_52_ctrl_stealReq_valid;
	output wire io_connSS_52_ctrl_stealReq_ready;
	input io_connSS_52_data_availableTask_ready;
	output wire io_connSS_52_data_availableTask_valid;
	output wire [255:0] io_connSS_52_data_availableTask_bits;
	output wire io_connSS_52_data_qOutTask_ready;
	input io_connSS_52_data_qOutTask_valid;
	input [255:0] io_connSS_52_data_qOutTask_bits;
	input io_connSS_53_ctrl_serveStealReq_valid;
	output wire io_connSS_53_ctrl_serveStealReq_ready;
	input io_connSS_53_ctrl_stealReq_valid;
	output wire io_connSS_53_ctrl_stealReq_ready;
	input io_connSS_53_data_availableTask_ready;
	output wire io_connSS_53_data_availableTask_valid;
	output wire [255:0] io_connSS_53_data_availableTask_bits;
	output wire io_connSS_53_data_qOutTask_ready;
	input io_connSS_53_data_qOutTask_valid;
	input [255:0] io_connSS_53_data_qOutTask_bits;
	input io_connSS_54_ctrl_serveStealReq_valid;
	output wire io_connSS_54_ctrl_serveStealReq_ready;
	input io_connSS_54_ctrl_stealReq_valid;
	output wire io_connSS_54_ctrl_stealReq_ready;
	input io_connSS_54_data_availableTask_ready;
	output wire io_connSS_54_data_availableTask_valid;
	output wire [255:0] io_connSS_54_data_availableTask_bits;
	output wire io_connSS_54_data_qOutTask_ready;
	input io_connSS_54_data_qOutTask_valid;
	input [255:0] io_connSS_54_data_qOutTask_bits;
	input io_connSS_55_ctrl_serveStealReq_valid;
	output wire io_connSS_55_ctrl_serveStealReq_ready;
	input io_connSS_55_ctrl_stealReq_valid;
	output wire io_connSS_55_ctrl_stealReq_ready;
	input io_connSS_55_data_availableTask_ready;
	output wire io_connSS_55_data_availableTask_valid;
	output wire [255:0] io_connSS_55_data_availableTask_bits;
	output wire io_connSS_55_data_qOutTask_ready;
	input io_connSS_55_data_qOutTask_valid;
	input [255:0] io_connSS_55_data_qOutTask_bits;
	input io_connSS_56_ctrl_serveStealReq_valid;
	output wire io_connSS_56_ctrl_serveStealReq_ready;
	input io_connSS_56_ctrl_stealReq_valid;
	output wire io_connSS_56_ctrl_stealReq_ready;
	input io_connSS_56_data_availableTask_ready;
	output wire io_connSS_56_data_availableTask_valid;
	output wire [255:0] io_connSS_56_data_availableTask_bits;
	output wire io_connSS_56_data_qOutTask_ready;
	input io_connSS_56_data_qOutTask_valid;
	input [255:0] io_connSS_56_data_qOutTask_bits;
	input io_connSS_57_ctrl_serveStealReq_valid;
	output wire io_connSS_57_ctrl_serveStealReq_ready;
	input io_connSS_57_ctrl_stealReq_valid;
	output wire io_connSS_57_ctrl_stealReq_ready;
	input io_connSS_57_data_availableTask_ready;
	output wire io_connSS_57_data_availableTask_valid;
	output wire [255:0] io_connSS_57_data_availableTask_bits;
	output wire io_connSS_57_data_qOutTask_ready;
	input io_connSS_57_data_qOutTask_valid;
	input [255:0] io_connSS_57_data_qOutTask_bits;
	input io_connSS_58_ctrl_serveStealReq_valid;
	output wire io_connSS_58_ctrl_serveStealReq_ready;
	input io_connSS_58_ctrl_stealReq_valid;
	output wire io_connSS_58_ctrl_stealReq_ready;
	input io_connSS_58_data_availableTask_ready;
	output wire io_connSS_58_data_availableTask_valid;
	output wire [255:0] io_connSS_58_data_availableTask_bits;
	output wire io_connSS_58_data_qOutTask_ready;
	input io_connSS_58_data_qOutTask_valid;
	input [255:0] io_connSS_58_data_qOutTask_bits;
	input io_connSS_59_ctrl_serveStealReq_valid;
	output wire io_connSS_59_ctrl_serveStealReq_ready;
	input io_connSS_59_ctrl_stealReq_valid;
	output wire io_connSS_59_ctrl_stealReq_ready;
	input io_connSS_59_data_availableTask_ready;
	output wire io_connSS_59_data_availableTask_valid;
	output wire [255:0] io_connSS_59_data_availableTask_bits;
	output wire io_connSS_59_data_qOutTask_ready;
	input io_connSS_59_data_qOutTask_valid;
	input [255:0] io_connSS_59_data_qOutTask_bits;
	input io_connSS_60_ctrl_serveStealReq_valid;
	output wire io_connSS_60_ctrl_serveStealReq_ready;
	input io_connSS_60_ctrl_stealReq_valid;
	output wire io_connSS_60_ctrl_stealReq_ready;
	input io_connSS_60_data_availableTask_ready;
	output wire io_connSS_60_data_availableTask_valid;
	output wire [255:0] io_connSS_60_data_availableTask_bits;
	output wire io_connSS_60_data_qOutTask_ready;
	input io_connSS_60_data_qOutTask_valid;
	input [255:0] io_connSS_60_data_qOutTask_bits;
	input io_connSS_61_ctrl_serveStealReq_valid;
	output wire io_connSS_61_ctrl_serveStealReq_ready;
	input io_connSS_61_ctrl_stealReq_valid;
	output wire io_connSS_61_ctrl_stealReq_ready;
	input io_connSS_61_data_availableTask_ready;
	output wire io_connSS_61_data_availableTask_valid;
	output wire [255:0] io_connSS_61_data_availableTask_bits;
	output wire io_connSS_61_data_qOutTask_ready;
	input io_connSS_61_data_qOutTask_valid;
	input [255:0] io_connSS_61_data_qOutTask_bits;
	input io_connSS_62_ctrl_serveStealReq_valid;
	output wire io_connSS_62_ctrl_serveStealReq_ready;
	input io_connSS_62_ctrl_stealReq_valid;
	output wire io_connSS_62_ctrl_stealReq_ready;
	input io_connSS_62_data_availableTask_ready;
	output wire io_connSS_62_data_availableTask_valid;
	output wire [255:0] io_connSS_62_data_availableTask_bits;
	output wire io_connSS_62_data_qOutTask_ready;
	input io_connSS_62_data_qOutTask_valid;
	input [255:0] io_connSS_62_data_qOutTask_bits;
	input io_connSS_63_ctrl_serveStealReq_valid;
	output wire io_connSS_63_ctrl_serveStealReq_ready;
	input io_connSS_63_ctrl_stealReq_valid;
	output wire io_connSS_63_ctrl_stealReq_ready;
	input io_connSS_63_data_availableTask_ready;
	output wire io_connSS_63_data_availableTask_valid;
	output wire [255:0] io_connSS_63_data_availableTask_bits;
	output wire io_connSS_63_data_qOutTask_ready;
	input io_connSS_63_data_qOutTask_valid;
	input [255:0] io_connSS_63_data_qOutTask_bits;
	input io_connSS_64_ctrl_serveStealReq_valid;
	output wire io_connSS_64_ctrl_serveStealReq_ready;
	input io_connSS_64_ctrl_stealReq_valid;
	output wire io_connSS_64_ctrl_stealReq_ready;
	input io_connSS_64_data_availableTask_ready;
	output wire io_connSS_64_data_availableTask_valid;
	output wire [255:0] io_connSS_64_data_availableTask_bits;
	output wire io_connSS_64_data_qOutTask_ready;
	input io_connSS_64_data_qOutTask_valid;
	input [255:0] io_connSS_64_data_qOutTask_bits;
	input io_connSS_65_ctrl_serveStealReq_valid;
	output wire io_connSS_65_ctrl_serveStealReq_ready;
	input io_connSS_65_ctrl_stealReq_valid;
	output wire io_connSS_65_ctrl_stealReq_ready;
	input io_connSS_65_data_availableTask_ready;
	output wire io_connSS_65_data_availableTask_valid;
	output wire [255:0] io_connSS_65_data_availableTask_bits;
	output wire io_connSS_65_data_qOutTask_ready;
	input io_connSS_65_data_qOutTask_valid;
	input [255:0] io_connSS_65_data_qOutTask_bits;
	input io_connSS_66_ctrl_serveStealReq_valid;
	output wire io_connSS_66_ctrl_serveStealReq_ready;
	input io_connSS_66_ctrl_stealReq_valid;
	output wire io_connSS_66_ctrl_stealReq_ready;
	input io_connSS_66_data_availableTask_ready;
	output wire io_connSS_66_data_availableTask_valid;
	output wire [255:0] io_connSS_66_data_availableTask_bits;
	output wire io_connSS_66_data_qOutTask_ready;
	input io_connSS_66_data_qOutTask_valid;
	input [255:0] io_connSS_66_data_qOutTask_bits;
	input io_connSS_67_ctrl_serveStealReq_valid;
	output wire io_connSS_67_ctrl_serveStealReq_ready;
	input io_connSS_67_ctrl_stealReq_valid;
	output wire io_connSS_67_ctrl_stealReq_ready;
	input io_connSS_67_data_availableTask_ready;
	output wire io_connSS_67_data_availableTask_valid;
	output wire [255:0] io_connSS_67_data_availableTask_bits;
	output wire io_connSS_67_data_qOutTask_ready;
	input io_connSS_67_data_qOutTask_valid;
	input [255:0] io_connSS_67_data_qOutTask_bits;
	input io_connSS_68_ctrl_serveStealReq_valid;
	output wire io_connSS_68_ctrl_serveStealReq_ready;
	input io_connSS_68_ctrl_stealReq_valid;
	output wire io_connSS_68_ctrl_stealReq_ready;
	input io_connSS_68_data_availableTask_ready;
	output wire io_connSS_68_data_availableTask_valid;
	output wire [255:0] io_connSS_68_data_availableTask_bits;
	output wire io_connSS_68_data_qOutTask_ready;
	input io_connSS_68_data_qOutTask_valid;
	input [255:0] io_connSS_68_data_qOutTask_bits;
	input io_connSS_69_ctrl_serveStealReq_valid;
	output wire io_connSS_69_ctrl_serveStealReq_ready;
	input io_connSS_69_ctrl_stealReq_valid;
	output wire io_connSS_69_ctrl_stealReq_ready;
	input io_connSS_69_data_availableTask_ready;
	output wire io_connSS_69_data_availableTask_valid;
	output wire [255:0] io_connSS_69_data_availableTask_bits;
	output wire io_connSS_69_data_qOutTask_ready;
	input io_connSS_69_data_qOutTask_valid;
	input [255:0] io_connSS_69_data_qOutTask_bits;
	input io_connSS_70_ctrl_serveStealReq_valid;
	output wire io_connSS_70_ctrl_serveStealReq_ready;
	input io_connSS_70_ctrl_stealReq_valid;
	output wire io_connSS_70_ctrl_stealReq_ready;
	input io_connSS_70_data_availableTask_ready;
	output wire io_connSS_70_data_availableTask_valid;
	output wire [255:0] io_connSS_70_data_availableTask_bits;
	output wire io_connSS_70_data_qOutTask_ready;
	input io_connSS_70_data_qOutTask_valid;
	input [255:0] io_connSS_70_data_qOutTask_bits;
	input io_connSS_71_ctrl_serveStealReq_valid;
	output wire io_connSS_71_ctrl_serveStealReq_ready;
	input io_connSS_71_ctrl_stealReq_valid;
	output wire io_connSS_71_ctrl_stealReq_ready;
	input io_connSS_71_data_availableTask_ready;
	output wire io_connSS_71_data_availableTask_valid;
	output wire [255:0] io_connSS_71_data_availableTask_bits;
	output wire io_connSS_71_data_qOutTask_ready;
	input io_connSS_71_data_qOutTask_valid;
	input [255:0] io_connSS_71_data_qOutTask_bits;
	input io_connSS_72_ctrl_serveStealReq_valid;
	output wire io_connSS_72_ctrl_serveStealReq_ready;
	input io_connSS_72_ctrl_stealReq_valid;
	output wire io_connSS_72_ctrl_stealReq_ready;
	input io_connSS_72_data_availableTask_ready;
	output wire io_connSS_72_data_availableTask_valid;
	output wire [255:0] io_connSS_72_data_availableTask_bits;
	output wire io_connSS_72_data_qOutTask_ready;
	input io_connSS_72_data_qOutTask_valid;
	input [255:0] io_connSS_72_data_qOutTask_bits;
	input io_connSS_73_ctrl_serveStealReq_valid;
	output wire io_connSS_73_ctrl_serveStealReq_ready;
	input io_connSS_73_ctrl_stealReq_valid;
	output wire io_connSS_73_ctrl_stealReq_ready;
	input io_connSS_73_data_availableTask_ready;
	output wire io_connSS_73_data_availableTask_valid;
	output wire [255:0] io_connSS_73_data_availableTask_bits;
	output wire io_connSS_73_data_qOutTask_ready;
	input io_connSS_73_data_qOutTask_valid;
	input [255:0] io_connSS_73_data_qOutTask_bits;
	input io_connSS_74_ctrl_serveStealReq_valid;
	output wire io_connSS_74_ctrl_serveStealReq_ready;
	input io_connSS_74_ctrl_stealReq_valid;
	output wire io_connSS_74_ctrl_stealReq_ready;
	input io_connSS_74_data_availableTask_ready;
	output wire io_connSS_74_data_availableTask_valid;
	output wire [255:0] io_connSS_74_data_availableTask_bits;
	output wire io_connSS_74_data_qOutTask_ready;
	input io_connSS_74_data_qOutTask_valid;
	input [255:0] io_connSS_74_data_qOutTask_bits;
	input io_connSS_75_ctrl_serveStealReq_valid;
	output wire io_connSS_75_ctrl_serveStealReq_ready;
	input io_connSS_75_ctrl_stealReq_valid;
	output wire io_connSS_75_ctrl_stealReq_ready;
	input io_connSS_75_data_availableTask_ready;
	output wire io_connSS_75_data_availableTask_valid;
	output wire [255:0] io_connSS_75_data_availableTask_bits;
	output wire io_connSS_75_data_qOutTask_ready;
	input io_connSS_75_data_qOutTask_valid;
	input [255:0] io_connSS_75_data_qOutTask_bits;
	input io_connSS_76_ctrl_serveStealReq_valid;
	output wire io_connSS_76_ctrl_serveStealReq_ready;
	input io_connSS_76_ctrl_stealReq_valid;
	output wire io_connSS_76_ctrl_stealReq_ready;
	input io_connSS_76_data_availableTask_ready;
	output wire io_connSS_76_data_availableTask_valid;
	output wire [255:0] io_connSS_76_data_availableTask_bits;
	output wire io_connSS_76_data_qOutTask_ready;
	input io_connSS_76_data_qOutTask_valid;
	input [255:0] io_connSS_76_data_qOutTask_bits;
	input io_connSS_77_ctrl_serveStealReq_valid;
	output wire io_connSS_77_ctrl_serveStealReq_ready;
	input io_connSS_77_ctrl_stealReq_valid;
	output wire io_connSS_77_ctrl_stealReq_ready;
	input io_connSS_77_data_availableTask_ready;
	output wire io_connSS_77_data_availableTask_valid;
	output wire [255:0] io_connSS_77_data_availableTask_bits;
	output wire io_connSS_77_data_qOutTask_ready;
	input io_connSS_77_data_qOutTask_valid;
	input [255:0] io_connSS_77_data_qOutTask_bits;
	input io_connSS_78_ctrl_serveStealReq_valid;
	output wire io_connSS_78_ctrl_serveStealReq_ready;
	input io_connSS_78_ctrl_stealReq_valid;
	output wire io_connSS_78_ctrl_stealReq_ready;
	input io_connSS_78_data_availableTask_ready;
	output wire io_connSS_78_data_availableTask_valid;
	output wire [255:0] io_connSS_78_data_availableTask_bits;
	output wire io_connSS_78_data_qOutTask_ready;
	input io_connSS_78_data_qOutTask_valid;
	input [255:0] io_connSS_78_data_qOutTask_bits;
	input io_connSS_79_ctrl_serveStealReq_valid;
	output wire io_connSS_79_ctrl_serveStealReq_ready;
	input io_connSS_79_ctrl_stealReq_valid;
	output wire io_connSS_79_ctrl_stealReq_ready;
	input io_connSS_79_data_availableTask_ready;
	output wire io_connSS_79_data_availableTask_valid;
	output wire [255:0] io_connSS_79_data_availableTask_bits;
	output wire io_connSS_79_data_qOutTask_ready;
	input io_connSS_79_data_qOutTask_valid;
	input [255:0] io_connSS_79_data_qOutTask_bits;
	input io_connSS_80_ctrl_serveStealReq_valid;
	output wire io_connSS_80_ctrl_serveStealReq_ready;
	input io_connSS_80_ctrl_stealReq_valid;
	output wire io_connSS_80_ctrl_stealReq_ready;
	input io_connSS_80_data_availableTask_ready;
	output wire io_connSS_80_data_availableTask_valid;
	output wire [255:0] io_connSS_80_data_availableTask_bits;
	output wire io_connSS_80_data_qOutTask_ready;
	input io_connSS_80_data_qOutTask_valid;
	input [255:0] io_connSS_80_data_qOutTask_bits;
	input io_connSS_81_ctrl_serveStealReq_valid;
	output wire io_connSS_81_ctrl_serveStealReq_ready;
	input io_connSS_81_ctrl_stealReq_valid;
	output wire io_connSS_81_ctrl_stealReq_ready;
	input io_connSS_81_data_availableTask_ready;
	output wire io_connSS_81_data_availableTask_valid;
	output wire [255:0] io_connSS_81_data_availableTask_bits;
	output wire io_connSS_81_data_qOutTask_ready;
	input io_connSS_81_data_qOutTask_valid;
	input [255:0] io_connSS_81_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	output wire io_ntwDataUnitOccupancyVSS_1;
	wire _ctrlunits_81_io_reqTaskOut;
	wire _ctrlunits_80_io_reqTaskOut;
	wire _ctrlunits_79_io_reqTaskOut;
	wire _ctrlunits_78_io_reqTaskOut;
	wire _ctrlunits_77_io_reqTaskOut;
	wire _ctrlunits_76_io_reqTaskOut;
	wire _ctrlunits_75_io_reqTaskOut;
	wire _ctrlunits_74_io_reqTaskOut;
	wire _ctrlunits_73_io_reqTaskOut;
	wire _ctrlunits_72_io_reqTaskOut;
	wire _ctrlunits_71_io_reqTaskOut;
	wire _ctrlunits_70_io_reqTaskOut;
	wire _ctrlunits_69_io_reqTaskOut;
	wire _ctrlunits_68_io_reqTaskOut;
	wire _ctrlunits_67_io_reqTaskOut;
	wire _ctrlunits_66_io_reqTaskOut;
	wire _ctrlunits_65_io_reqTaskOut;
	wire _ctrlunits_64_io_reqTaskOut;
	wire _ctrlunits_63_io_reqTaskOut;
	wire _ctrlunits_62_io_reqTaskOut;
	wire _ctrlunits_61_io_reqTaskOut;
	wire _ctrlunits_60_io_reqTaskOut;
	wire _ctrlunits_59_io_reqTaskOut;
	wire _ctrlunits_58_io_reqTaskOut;
	wire _ctrlunits_57_io_reqTaskOut;
	wire _ctrlunits_56_io_reqTaskOut;
	wire _ctrlunits_55_io_reqTaskOut;
	wire _ctrlunits_54_io_reqTaskOut;
	wire _ctrlunits_53_io_reqTaskOut;
	wire _ctrlunits_52_io_reqTaskOut;
	wire _ctrlunits_51_io_reqTaskOut;
	wire _ctrlunits_50_io_reqTaskOut;
	wire _ctrlunits_49_io_reqTaskOut;
	wire _ctrlunits_48_io_reqTaskOut;
	wire _ctrlunits_47_io_reqTaskOut;
	wire _ctrlunits_46_io_reqTaskOut;
	wire _ctrlunits_45_io_reqTaskOut;
	wire _ctrlunits_44_io_reqTaskOut;
	wire _ctrlunits_43_io_reqTaskOut;
	wire _ctrlunits_42_io_reqTaskOut;
	wire _ctrlunits_41_io_reqTaskOut;
	wire _ctrlunits_40_io_reqTaskOut;
	wire _ctrlunits_39_io_reqTaskOut;
	wire _ctrlunits_38_io_reqTaskOut;
	wire _ctrlunits_37_io_reqTaskOut;
	wire _ctrlunits_36_io_reqTaskOut;
	wire _ctrlunits_35_io_reqTaskOut;
	wire _ctrlunits_34_io_reqTaskOut;
	wire _ctrlunits_33_io_reqTaskOut;
	wire _ctrlunits_32_io_reqTaskOut;
	wire _ctrlunits_31_io_reqTaskOut;
	wire _ctrlunits_30_io_reqTaskOut;
	wire _ctrlunits_29_io_reqTaskOut;
	wire _ctrlunits_28_io_reqTaskOut;
	wire _ctrlunits_27_io_reqTaskOut;
	wire _ctrlunits_26_io_reqTaskOut;
	wire _ctrlunits_25_io_reqTaskOut;
	wire _ctrlunits_24_io_reqTaskOut;
	wire _ctrlunits_23_io_reqTaskOut;
	wire _ctrlunits_22_io_reqTaskOut;
	wire _ctrlunits_21_io_reqTaskOut;
	wire _ctrlunits_20_io_reqTaskOut;
	wire _ctrlunits_19_io_reqTaskOut;
	wire _ctrlunits_18_io_reqTaskOut;
	wire _ctrlunits_17_io_reqTaskOut;
	wire _ctrlunits_16_io_reqTaskOut;
	wire _ctrlunits_15_io_reqTaskOut;
	wire _ctrlunits_14_io_reqTaskOut;
	wire _ctrlunits_13_io_reqTaskOut;
	wire _ctrlunits_12_io_reqTaskOut;
	wire _ctrlunits_11_io_reqTaskOut;
	wire _ctrlunits_10_io_reqTaskOut;
	wire _ctrlunits_9_io_reqTaskOut;
	wire _ctrlunits_8_io_reqTaskOut;
	wire _ctrlunits_7_io_reqTaskOut;
	wire _ctrlunits_6_io_reqTaskOut;
	wire _ctrlunits_5_io_reqTaskOut;
	wire _ctrlunits_4_io_reqTaskOut;
	wire _ctrlunits_3_io_reqTaskOut;
	wire _ctrlunits_2_io_reqTaskOut;
	wire _ctrlunits_1_io_reqTaskOut;
	wire _ctrlunits_0_io_reqTaskOut;
	wire [255:0] _dataUnits_81_io_taskOut;
	wire _dataUnits_81_io_validOut;
	wire [255:0] _dataUnits_80_io_taskOut;
	wire _dataUnits_80_io_validOut;
	wire [255:0] _dataUnits_79_io_taskOut;
	wire _dataUnits_79_io_validOut;
	wire [255:0] _dataUnits_78_io_taskOut;
	wire _dataUnits_78_io_validOut;
	wire [255:0] _dataUnits_77_io_taskOut;
	wire _dataUnits_77_io_validOut;
	wire [255:0] _dataUnits_76_io_taskOut;
	wire _dataUnits_76_io_validOut;
	wire [255:0] _dataUnits_75_io_taskOut;
	wire _dataUnits_75_io_validOut;
	wire [255:0] _dataUnits_74_io_taskOut;
	wire _dataUnits_74_io_validOut;
	wire [255:0] _dataUnits_73_io_taskOut;
	wire _dataUnits_73_io_validOut;
	wire [255:0] _dataUnits_72_io_taskOut;
	wire _dataUnits_72_io_validOut;
	wire [255:0] _dataUnits_71_io_taskOut;
	wire _dataUnits_71_io_validOut;
	wire [255:0] _dataUnits_70_io_taskOut;
	wire _dataUnits_70_io_validOut;
	wire [255:0] _dataUnits_69_io_taskOut;
	wire _dataUnits_69_io_validOut;
	wire [255:0] _dataUnits_68_io_taskOut;
	wire _dataUnits_68_io_validOut;
	wire [255:0] _dataUnits_67_io_taskOut;
	wire _dataUnits_67_io_validOut;
	wire [255:0] _dataUnits_66_io_taskOut;
	wire _dataUnits_66_io_validOut;
	wire [255:0] _dataUnits_65_io_taskOut;
	wire _dataUnits_65_io_validOut;
	wire [255:0] _dataUnits_64_io_taskOut;
	wire _dataUnits_64_io_validOut;
	wire [255:0] _dataUnits_63_io_taskOut;
	wire _dataUnits_63_io_validOut;
	wire [255:0] _dataUnits_62_io_taskOut;
	wire _dataUnits_62_io_validOut;
	wire [255:0] _dataUnits_61_io_taskOut;
	wire _dataUnits_61_io_validOut;
	wire [255:0] _dataUnits_60_io_taskOut;
	wire _dataUnits_60_io_validOut;
	wire [255:0] _dataUnits_59_io_taskOut;
	wire _dataUnits_59_io_validOut;
	wire [255:0] _dataUnits_58_io_taskOut;
	wire _dataUnits_58_io_validOut;
	wire [255:0] _dataUnits_57_io_taskOut;
	wire _dataUnits_57_io_validOut;
	wire [255:0] _dataUnits_56_io_taskOut;
	wire _dataUnits_56_io_validOut;
	wire [255:0] _dataUnits_55_io_taskOut;
	wire _dataUnits_55_io_validOut;
	wire [255:0] _dataUnits_54_io_taskOut;
	wire _dataUnits_54_io_validOut;
	wire [255:0] _dataUnits_53_io_taskOut;
	wire _dataUnits_53_io_validOut;
	wire [255:0] _dataUnits_52_io_taskOut;
	wire _dataUnits_52_io_validOut;
	wire [255:0] _dataUnits_51_io_taskOut;
	wire _dataUnits_51_io_validOut;
	wire [255:0] _dataUnits_50_io_taskOut;
	wire _dataUnits_50_io_validOut;
	wire [255:0] _dataUnits_49_io_taskOut;
	wire _dataUnits_49_io_validOut;
	wire [255:0] _dataUnits_48_io_taskOut;
	wire _dataUnits_48_io_validOut;
	wire [255:0] _dataUnits_47_io_taskOut;
	wire _dataUnits_47_io_validOut;
	wire [255:0] _dataUnits_46_io_taskOut;
	wire _dataUnits_46_io_validOut;
	wire [255:0] _dataUnits_45_io_taskOut;
	wire _dataUnits_45_io_validOut;
	wire [255:0] _dataUnits_44_io_taskOut;
	wire _dataUnits_44_io_validOut;
	wire [255:0] _dataUnits_43_io_taskOut;
	wire _dataUnits_43_io_validOut;
	wire [255:0] _dataUnits_42_io_taskOut;
	wire _dataUnits_42_io_validOut;
	wire [255:0] _dataUnits_41_io_taskOut;
	wire _dataUnits_41_io_validOut;
	wire [255:0] _dataUnits_40_io_taskOut;
	wire _dataUnits_40_io_validOut;
	wire [255:0] _dataUnits_39_io_taskOut;
	wire _dataUnits_39_io_validOut;
	wire [255:0] _dataUnits_38_io_taskOut;
	wire _dataUnits_38_io_validOut;
	wire [255:0] _dataUnits_37_io_taskOut;
	wire _dataUnits_37_io_validOut;
	wire [255:0] _dataUnits_36_io_taskOut;
	wire _dataUnits_36_io_validOut;
	wire [255:0] _dataUnits_35_io_taskOut;
	wire _dataUnits_35_io_validOut;
	wire [255:0] _dataUnits_34_io_taskOut;
	wire _dataUnits_34_io_validOut;
	wire [255:0] _dataUnits_33_io_taskOut;
	wire _dataUnits_33_io_validOut;
	wire [255:0] _dataUnits_32_io_taskOut;
	wire _dataUnits_32_io_validOut;
	wire [255:0] _dataUnits_31_io_taskOut;
	wire _dataUnits_31_io_validOut;
	wire [255:0] _dataUnits_30_io_taskOut;
	wire _dataUnits_30_io_validOut;
	wire [255:0] _dataUnits_29_io_taskOut;
	wire _dataUnits_29_io_validOut;
	wire [255:0] _dataUnits_28_io_taskOut;
	wire _dataUnits_28_io_validOut;
	wire [255:0] _dataUnits_27_io_taskOut;
	wire _dataUnits_27_io_validOut;
	wire [255:0] _dataUnits_26_io_taskOut;
	wire _dataUnits_26_io_validOut;
	wire [255:0] _dataUnits_25_io_taskOut;
	wire _dataUnits_25_io_validOut;
	wire [255:0] _dataUnits_24_io_taskOut;
	wire _dataUnits_24_io_validOut;
	wire [255:0] _dataUnits_23_io_taskOut;
	wire _dataUnits_23_io_validOut;
	wire [255:0] _dataUnits_22_io_taskOut;
	wire _dataUnits_22_io_validOut;
	wire [255:0] _dataUnits_21_io_taskOut;
	wire _dataUnits_21_io_validOut;
	wire [255:0] _dataUnits_20_io_taskOut;
	wire _dataUnits_20_io_validOut;
	wire [255:0] _dataUnits_19_io_taskOut;
	wire _dataUnits_19_io_validOut;
	wire [255:0] _dataUnits_18_io_taskOut;
	wire _dataUnits_18_io_validOut;
	wire [255:0] _dataUnits_17_io_taskOut;
	wire _dataUnits_17_io_validOut;
	wire [255:0] _dataUnits_16_io_taskOut;
	wire _dataUnits_16_io_validOut;
	wire [255:0] _dataUnits_15_io_taskOut;
	wire _dataUnits_15_io_validOut;
	wire [255:0] _dataUnits_14_io_taskOut;
	wire _dataUnits_14_io_validOut;
	wire [255:0] _dataUnits_13_io_taskOut;
	wire _dataUnits_13_io_validOut;
	wire [255:0] _dataUnits_12_io_taskOut;
	wire _dataUnits_12_io_validOut;
	wire [255:0] _dataUnits_11_io_taskOut;
	wire _dataUnits_11_io_validOut;
	wire [255:0] _dataUnits_10_io_taskOut;
	wire _dataUnits_10_io_validOut;
	wire [255:0] _dataUnits_9_io_taskOut;
	wire _dataUnits_9_io_validOut;
	wire [255:0] _dataUnits_8_io_taskOut;
	wire _dataUnits_8_io_validOut;
	wire [255:0] _dataUnits_7_io_taskOut;
	wire _dataUnits_7_io_validOut;
	wire [255:0] _dataUnits_6_io_taskOut;
	wire _dataUnits_6_io_validOut;
	wire [255:0] _dataUnits_5_io_taskOut;
	wire _dataUnits_5_io_validOut;
	wire [255:0] _dataUnits_4_io_taskOut;
	wire _dataUnits_4_io_validOut;
	wire [255:0] _dataUnits_3_io_taskOut;
	wire _dataUnits_3_io_validOut;
	wire [255:0] _dataUnits_2_io_taskOut;
	wire _dataUnits_2_io_validOut;
	wire [255:0] _dataUnits_1_io_taskOut;
	wire _dataUnits_1_io_validOut;
	wire [255:0] _dataUnits_0_io_taskOut;
	wire _dataUnits_0_io_validOut;
	SchedulerNetworkDataUnit_66 dataUnits_0(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_81_io_taskOut),
		.io_taskOut(_dataUnits_0_io_taskOut),
		.io_validIn(_dataUnits_81_io_validOut),
		.io_validOut(_dataUnits_0_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_0_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_0_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_0_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_0_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_0_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_0_data_qOutTask_bits),
		.io_occupied(io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerNetworkDataUnit_66 dataUnits_1(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_0_io_taskOut),
		.io_taskOut(_dataUnits_1_io_taskOut),
		.io_validIn(_dataUnits_0_io_validOut),
		.io_validOut(_dataUnits_1_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_1_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_1_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_1_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_1_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_1_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_1_data_qOutTask_bits),
		.io_occupied(io_ntwDataUnitOccupancyVSS_1)
	);
	SchedulerNetworkDataUnit_66 dataUnits_2(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_1_io_taskOut),
		.io_taskOut(_dataUnits_2_io_taskOut),
		.io_validIn(_dataUnits_1_io_validOut),
		.io_validOut(_dataUnits_2_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_2_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_2_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_2_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_3(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_2_io_taskOut),
		.io_taskOut(_dataUnits_3_io_taskOut),
		.io_validIn(_dataUnits_2_io_validOut),
		.io_validOut(_dataUnits_3_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_3_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_3_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_3_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_4(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_3_io_taskOut),
		.io_taskOut(_dataUnits_4_io_taskOut),
		.io_validIn(_dataUnits_3_io_validOut),
		.io_validOut(_dataUnits_4_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_4_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_4_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_4_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_5(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_4_io_taskOut),
		.io_taskOut(_dataUnits_5_io_taskOut),
		.io_validIn(_dataUnits_4_io_validOut),
		.io_validOut(_dataUnits_5_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_5_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_5_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_5_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_6(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_5_io_taskOut),
		.io_taskOut(_dataUnits_6_io_taskOut),
		.io_validIn(_dataUnits_5_io_validOut),
		.io_validOut(_dataUnits_6_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_6_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_6_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_6_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_7(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_6_io_taskOut),
		.io_taskOut(_dataUnits_7_io_taskOut),
		.io_validIn(_dataUnits_6_io_validOut),
		.io_validOut(_dataUnits_7_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_7_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_7_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_7_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_8(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_7_io_taskOut),
		.io_taskOut(_dataUnits_8_io_taskOut),
		.io_validIn(_dataUnits_7_io_validOut),
		.io_validOut(_dataUnits_8_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_8_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_8_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_8_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_9(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_8_io_taskOut),
		.io_taskOut(_dataUnits_9_io_taskOut),
		.io_validIn(_dataUnits_8_io_validOut),
		.io_validOut(_dataUnits_9_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_9_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_9_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_9_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_10(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_9_io_taskOut),
		.io_taskOut(_dataUnits_10_io_taskOut),
		.io_validIn(_dataUnits_9_io_validOut),
		.io_validOut(_dataUnits_10_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_10_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_10_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_10_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_11(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_10_io_taskOut),
		.io_taskOut(_dataUnits_11_io_taskOut),
		.io_validIn(_dataUnits_10_io_validOut),
		.io_validOut(_dataUnits_11_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_11_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_11_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_11_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_12(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_11_io_taskOut),
		.io_taskOut(_dataUnits_12_io_taskOut),
		.io_validIn(_dataUnits_11_io_validOut),
		.io_validOut(_dataUnits_12_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_12_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_12_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_12_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_13(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_12_io_taskOut),
		.io_taskOut(_dataUnits_13_io_taskOut),
		.io_validIn(_dataUnits_12_io_validOut),
		.io_validOut(_dataUnits_13_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_13_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_13_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_13_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_14(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_13_io_taskOut),
		.io_taskOut(_dataUnits_14_io_taskOut),
		.io_validIn(_dataUnits_13_io_validOut),
		.io_validOut(_dataUnits_14_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_14_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_14_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_14_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_15(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_14_io_taskOut),
		.io_taskOut(_dataUnits_15_io_taskOut),
		.io_validIn(_dataUnits_14_io_validOut),
		.io_validOut(_dataUnits_15_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_15_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_15_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_15_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_16(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_15_io_taskOut),
		.io_taskOut(_dataUnits_16_io_taskOut),
		.io_validIn(_dataUnits_15_io_validOut),
		.io_validOut(_dataUnits_16_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_16_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_16_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_16_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_17(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_16_io_taskOut),
		.io_taskOut(_dataUnits_17_io_taskOut),
		.io_validIn(_dataUnits_16_io_validOut),
		.io_validOut(_dataUnits_17_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_17_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_17_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_17_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_18(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_17_io_taskOut),
		.io_taskOut(_dataUnits_18_io_taskOut),
		.io_validIn(_dataUnits_17_io_validOut),
		.io_validOut(_dataUnits_18_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_18_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_18_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_18_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_18_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_18_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_18_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_19(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_18_io_taskOut),
		.io_taskOut(_dataUnits_19_io_taskOut),
		.io_validIn(_dataUnits_18_io_validOut),
		.io_validOut(_dataUnits_19_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_19_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_19_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_19_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_19_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_19_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_19_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_20(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_19_io_taskOut),
		.io_taskOut(_dataUnits_20_io_taskOut),
		.io_validIn(_dataUnits_19_io_validOut),
		.io_validOut(_dataUnits_20_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_20_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_20_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_20_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_20_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_20_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_20_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_21(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_20_io_taskOut),
		.io_taskOut(_dataUnits_21_io_taskOut),
		.io_validIn(_dataUnits_20_io_validOut),
		.io_validOut(_dataUnits_21_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_21_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_21_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_21_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_21_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_21_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_21_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_22(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_21_io_taskOut),
		.io_taskOut(_dataUnits_22_io_taskOut),
		.io_validIn(_dataUnits_21_io_validOut),
		.io_validOut(_dataUnits_22_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_22_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_22_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_22_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_22_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_22_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_22_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_23(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_22_io_taskOut),
		.io_taskOut(_dataUnits_23_io_taskOut),
		.io_validIn(_dataUnits_22_io_validOut),
		.io_validOut(_dataUnits_23_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_23_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_23_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_23_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_23_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_23_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_23_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_24(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_23_io_taskOut),
		.io_taskOut(_dataUnits_24_io_taskOut),
		.io_validIn(_dataUnits_23_io_validOut),
		.io_validOut(_dataUnits_24_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_24_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_24_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_24_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_24_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_24_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_24_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_25(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_24_io_taskOut),
		.io_taskOut(_dataUnits_25_io_taskOut),
		.io_validIn(_dataUnits_24_io_validOut),
		.io_validOut(_dataUnits_25_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_25_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_25_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_25_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_25_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_25_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_25_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_26(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_25_io_taskOut),
		.io_taskOut(_dataUnits_26_io_taskOut),
		.io_validIn(_dataUnits_25_io_validOut),
		.io_validOut(_dataUnits_26_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_26_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_26_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_26_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_26_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_26_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_26_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_27(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_26_io_taskOut),
		.io_taskOut(_dataUnits_27_io_taskOut),
		.io_validIn(_dataUnits_26_io_validOut),
		.io_validOut(_dataUnits_27_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_27_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_27_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_27_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_27_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_27_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_27_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_28(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_27_io_taskOut),
		.io_taskOut(_dataUnits_28_io_taskOut),
		.io_validIn(_dataUnits_27_io_validOut),
		.io_validOut(_dataUnits_28_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_28_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_28_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_28_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_28_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_28_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_28_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_29(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_28_io_taskOut),
		.io_taskOut(_dataUnits_29_io_taskOut),
		.io_validIn(_dataUnits_28_io_validOut),
		.io_validOut(_dataUnits_29_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_29_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_29_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_29_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_29_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_29_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_29_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_30(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_29_io_taskOut),
		.io_taskOut(_dataUnits_30_io_taskOut),
		.io_validIn(_dataUnits_29_io_validOut),
		.io_validOut(_dataUnits_30_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_30_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_30_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_30_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_30_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_30_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_30_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_31(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_30_io_taskOut),
		.io_taskOut(_dataUnits_31_io_taskOut),
		.io_validIn(_dataUnits_30_io_validOut),
		.io_validOut(_dataUnits_31_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_31_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_31_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_31_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_31_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_31_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_31_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_32(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_31_io_taskOut),
		.io_taskOut(_dataUnits_32_io_taskOut),
		.io_validIn(_dataUnits_31_io_validOut),
		.io_validOut(_dataUnits_32_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_32_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_32_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_32_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_32_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_32_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_32_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_33(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_32_io_taskOut),
		.io_taskOut(_dataUnits_33_io_taskOut),
		.io_validIn(_dataUnits_32_io_validOut),
		.io_validOut(_dataUnits_33_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_33_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_33_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_33_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_33_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_33_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_33_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_34(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_33_io_taskOut),
		.io_taskOut(_dataUnits_34_io_taskOut),
		.io_validIn(_dataUnits_33_io_validOut),
		.io_validOut(_dataUnits_34_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_34_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_34_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_34_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_34_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_34_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_34_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_35(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_34_io_taskOut),
		.io_taskOut(_dataUnits_35_io_taskOut),
		.io_validIn(_dataUnits_34_io_validOut),
		.io_validOut(_dataUnits_35_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_35_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_35_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_35_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_35_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_35_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_35_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_36(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_35_io_taskOut),
		.io_taskOut(_dataUnits_36_io_taskOut),
		.io_validIn(_dataUnits_35_io_validOut),
		.io_validOut(_dataUnits_36_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_36_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_36_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_36_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_36_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_36_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_36_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_37(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_36_io_taskOut),
		.io_taskOut(_dataUnits_37_io_taskOut),
		.io_validIn(_dataUnits_36_io_validOut),
		.io_validOut(_dataUnits_37_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_37_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_37_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_37_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_37_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_37_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_37_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_38(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_37_io_taskOut),
		.io_taskOut(_dataUnits_38_io_taskOut),
		.io_validIn(_dataUnits_37_io_validOut),
		.io_validOut(_dataUnits_38_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_38_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_38_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_38_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_38_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_38_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_38_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_39(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_38_io_taskOut),
		.io_taskOut(_dataUnits_39_io_taskOut),
		.io_validIn(_dataUnits_38_io_validOut),
		.io_validOut(_dataUnits_39_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_39_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_39_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_39_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_39_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_39_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_39_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_40(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_39_io_taskOut),
		.io_taskOut(_dataUnits_40_io_taskOut),
		.io_validIn(_dataUnits_39_io_validOut),
		.io_validOut(_dataUnits_40_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_40_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_40_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_40_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_40_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_40_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_40_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_41(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_40_io_taskOut),
		.io_taskOut(_dataUnits_41_io_taskOut),
		.io_validIn(_dataUnits_40_io_validOut),
		.io_validOut(_dataUnits_41_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_41_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_41_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_41_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_41_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_41_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_41_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_42(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_41_io_taskOut),
		.io_taskOut(_dataUnits_42_io_taskOut),
		.io_validIn(_dataUnits_41_io_validOut),
		.io_validOut(_dataUnits_42_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_42_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_42_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_42_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_42_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_42_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_42_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_43(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_42_io_taskOut),
		.io_taskOut(_dataUnits_43_io_taskOut),
		.io_validIn(_dataUnits_42_io_validOut),
		.io_validOut(_dataUnits_43_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_43_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_43_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_43_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_43_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_43_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_43_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_44(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_43_io_taskOut),
		.io_taskOut(_dataUnits_44_io_taskOut),
		.io_validIn(_dataUnits_43_io_validOut),
		.io_validOut(_dataUnits_44_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_44_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_44_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_44_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_44_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_44_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_44_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_45(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_44_io_taskOut),
		.io_taskOut(_dataUnits_45_io_taskOut),
		.io_validIn(_dataUnits_44_io_validOut),
		.io_validOut(_dataUnits_45_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_45_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_45_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_45_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_45_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_45_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_45_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_46(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_45_io_taskOut),
		.io_taskOut(_dataUnits_46_io_taskOut),
		.io_validIn(_dataUnits_45_io_validOut),
		.io_validOut(_dataUnits_46_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_46_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_46_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_46_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_46_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_46_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_46_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_47(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_46_io_taskOut),
		.io_taskOut(_dataUnits_47_io_taskOut),
		.io_validIn(_dataUnits_46_io_validOut),
		.io_validOut(_dataUnits_47_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_47_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_47_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_47_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_47_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_47_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_47_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_48(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_47_io_taskOut),
		.io_taskOut(_dataUnits_48_io_taskOut),
		.io_validIn(_dataUnits_47_io_validOut),
		.io_validOut(_dataUnits_48_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_48_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_48_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_48_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_48_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_48_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_48_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_49(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_48_io_taskOut),
		.io_taskOut(_dataUnits_49_io_taskOut),
		.io_validIn(_dataUnits_48_io_validOut),
		.io_validOut(_dataUnits_49_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_49_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_49_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_49_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_49_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_49_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_49_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_50(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_49_io_taskOut),
		.io_taskOut(_dataUnits_50_io_taskOut),
		.io_validIn(_dataUnits_49_io_validOut),
		.io_validOut(_dataUnits_50_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_50_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_50_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_50_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_50_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_50_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_50_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_51(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_50_io_taskOut),
		.io_taskOut(_dataUnits_51_io_taskOut),
		.io_validIn(_dataUnits_50_io_validOut),
		.io_validOut(_dataUnits_51_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_51_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_51_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_51_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_51_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_51_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_51_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_52(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_51_io_taskOut),
		.io_taskOut(_dataUnits_52_io_taskOut),
		.io_validIn(_dataUnits_51_io_validOut),
		.io_validOut(_dataUnits_52_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_52_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_52_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_52_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_52_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_52_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_52_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_53(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_52_io_taskOut),
		.io_taskOut(_dataUnits_53_io_taskOut),
		.io_validIn(_dataUnits_52_io_validOut),
		.io_validOut(_dataUnits_53_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_53_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_53_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_53_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_53_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_53_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_53_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_54(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_53_io_taskOut),
		.io_taskOut(_dataUnits_54_io_taskOut),
		.io_validIn(_dataUnits_53_io_validOut),
		.io_validOut(_dataUnits_54_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_54_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_54_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_54_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_54_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_54_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_54_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_55(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_54_io_taskOut),
		.io_taskOut(_dataUnits_55_io_taskOut),
		.io_validIn(_dataUnits_54_io_validOut),
		.io_validOut(_dataUnits_55_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_55_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_55_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_55_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_55_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_55_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_55_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_56(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_55_io_taskOut),
		.io_taskOut(_dataUnits_56_io_taskOut),
		.io_validIn(_dataUnits_55_io_validOut),
		.io_validOut(_dataUnits_56_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_56_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_56_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_56_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_56_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_56_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_56_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_57(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_56_io_taskOut),
		.io_taskOut(_dataUnits_57_io_taskOut),
		.io_validIn(_dataUnits_56_io_validOut),
		.io_validOut(_dataUnits_57_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_57_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_57_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_57_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_57_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_57_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_57_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_58(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_57_io_taskOut),
		.io_taskOut(_dataUnits_58_io_taskOut),
		.io_validIn(_dataUnits_57_io_validOut),
		.io_validOut(_dataUnits_58_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_58_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_58_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_58_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_58_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_58_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_58_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_59(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_58_io_taskOut),
		.io_taskOut(_dataUnits_59_io_taskOut),
		.io_validIn(_dataUnits_58_io_validOut),
		.io_validOut(_dataUnits_59_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_59_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_59_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_59_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_59_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_59_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_59_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_60(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_59_io_taskOut),
		.io_taskOut(_dataUnits_60_io_taskOut),
		.io_validIn(_dataUnits_59_io_validOut),
		.io_validOut(_dataUnits_60_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_60_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_60_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_60_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_60_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_60_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_60_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_61(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_60_io_taskOut),
		.io_taskOut(_dataUnits_61_io_taskOut),
		.io_validIn(_dataUnits_60_io_validOut),
		.io_validOut(_dataUnits_61_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_61_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_61_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_61_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_61_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_61_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_61_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_62(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_61_io_taskOut),
		.io_taskOut(_dataUnits_62_io_taskOut),
		.io_validIn(_dataUnits_61_io_validOut),
		.io_validOut(_dataUnits_62_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_62_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_62_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_62_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_62_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_62_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_62_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_63(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_62_io_taskOut),
		.io_taskOut(_dataUnits_63_io_taskOut),
		.io_validIn(_dataUnits_62_io_validOut),
		.io_validOut(_dataUnits_63_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_63_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_63_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_63_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_63_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_63_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_63_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_64(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_63_io_taskOut),
		.io_taskOut(_dataUnits_64_io_taskOut),
		.io_validIn(_dataUnits_63_io_validOut),
		.io_validOut(_dataUnits_64_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_64_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_64_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_64_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_64_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_64_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_64_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_65(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_64_io_taskOut),
		.io_taskOut(_dataUnits_65_io_taskOut),
		.io_validIn(_dataUnits_64_io_validOut),
		.io_validOut(_dataUnits_65_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_65_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_65_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_65_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_65_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_65_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_65_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_66(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_65_io_taskOut),
		.io_taskOut(_dataUnits_66_io_taskOut),
		.io_validIn(_dataUnits_65_io_validOut),
		.io_validOut(_dataUnits_66_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_66_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_66_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_66_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_66_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_66_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_66_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_67(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_66_io_taskOut),
		.io_taskOut(_dataUnits_67_io_taskOut),
		.io_validIn(_dataUnits_66_io_validOut),
		.io_validOut(_dataUnits_67_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_67_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_67_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_67_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_67_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_67_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_67_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_68(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_67_io_taskOut),
		.io_taskOut(_dataUnits_68_io_taskOut),
		.io_validIn(_dataUnits_67_io_validOut),
		.io_validOut(_dataUnits_68_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_68_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_68_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_68_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_68_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_68_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_68_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_69(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_68_io_taskOut),
		.io_taskOut(_dataUnits_69_io_taskOut),
		.io_validIn(_dataUnits_68_io_validOut),
		.io_validOut(_dataUnits_69_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_69_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_69_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_69_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_69_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_69_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_69_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_70(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_69_io_taskOut),
		.io_taskOut(_dataUnits_70_io_taskOut),
		.io_validIn(_dataUnits_69_io_validOut),
		.io_validOut(_dataUnits_70_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_70_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_70_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_70_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_70_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_70_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_70_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_71(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_70_io_taskOut),
		.io_taskOut(_dataUnits_71_io_taskOut),
		.io_validIn(_dataUnits_70_io_validOut),
		.io_validOut(_dataUnits_71_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_71_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_71_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_71_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_71_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_71_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_71_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_72(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_71_io_taskOut),
		.io_taskOut(_dataUnits_72_io_taskOut),
		.io_validIn(_dataUnits_71_io_validOut),
		.io_validOut(_dataUnits_72_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_72_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_72_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_72_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_72_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_72_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_72_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_73(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_72_io_taskOut),
		.io_taskOut(_dataUnits_73_io_taskOut),
		.io_validIn(_dataUnits_72_io_validOut),
		.io_validOut(_dataUnits_73_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_73_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_73_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_73_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_73_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_73_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_73_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_74(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_73_io_taskOut),
		.io_taskOut(_dataUnits_74_io_taskOut),
		.io_validIn(_dataUnits_73_io_validOut),
		.io_validOut(_dataUnits_74_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_74_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_74_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_74_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_74_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_74_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_74_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_75(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_74_io_taskOut),
		.io_taskOut(_dataUnits_75_io_taskOut),
		.io_validIn(_dataUnits_74_io_validOut),
		.io_validOut(_dataUnits_75_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_75_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_75_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_75_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_75_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_75_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_75_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_76(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_75_io_taskOut),
		.io_taskOut(_dataUnits_76_io_taskOut),
		.io_validIn(_dataUnits_75_io_validOut),
		.io_validOut(_dataUnits_76_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_76_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_76_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_76_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_76_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_76_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_76_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_77(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_76_io_taskOut),
		.io_taskOut(_dataUnits_77_io_taskOut),
		.io_validIn(_dataUnits_76_io_validOut),
		.io_validOut(_dataUnits_77_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_77_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_77_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_77_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_77_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_77_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_77_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_78(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_77_io_taskOut),
		.io_taskOut(_dataUnits_78_io_taskOut),
		.io_validIn(_dataUnits_77_io_validOut),
		.io_validOut(_dataUnits_78_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_78_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_78_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_78_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_78_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_78_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_78_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_79(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_78_io_taskOut),
		.io_taskOut(_dataUnits_79_io_taskOut),
		.io_validIn(_dataUnits_78_io_validOut),
		.io_validOut(_dataUnits_79_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_79_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_79_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_79_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_79_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_79_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_79_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_80(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_79_io_taskOut),
		.io_taskOut(_dataUnits_80_io_taskOut),
		.io_validIn(_dataUnits_79_io_validOut),
		.io_validOut(_dataUnits_80_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_80_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_80_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_80_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_80_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_80_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_80_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_66 dataUnits_81(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_80_io_taskOut),
		.io_taskOut(_dataUnits_81_io_taskOut),
		.io_validIn(_dataUnits_80_io_validOut),
		.io_validOut(_dataUnits_81_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_81_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_81_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_81_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_81_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_81_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_81_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkControlUnit ctrlunits_0(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_1_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_0_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_0_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_0_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_1(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_2_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_1_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_1_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_1_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_2(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_3_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_2_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_2_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_2_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_3(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_4_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_3_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_3_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_3_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_4(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_5_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_4_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_4_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_4_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_5(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_6_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_5_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_5_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_5_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_6(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_7_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_6_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_6_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_6_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_7(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_8_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_7_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_7_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_7_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_8(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_9_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_8_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_8_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_8_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_9(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_10_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_9_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_9_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_9_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_10(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_11_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_10_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_10_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_10_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_11(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_12_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_11_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_11_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_11_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_12(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_13_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_12_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_12_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_12_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_13(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_14_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_13_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_13_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_13_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_14(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_15_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_14_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_14_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_14_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_15(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_16_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_15_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_15_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_15_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_16(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_17_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_16_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_16_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_16_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_17(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_18_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_17_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_17_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_18(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_19_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_18_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_18_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_18_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_18_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_19(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_20_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_19_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_19_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_19_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_19_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_20(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_21_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_20_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_20_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_20_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_20_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_21(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_22_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_21_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_21_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_21_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_21_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_22(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_23_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_22_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_22_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_22_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_22_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_23(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_24_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_23_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_23_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_23_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_23_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_24(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_25_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_24_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_24_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_24_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_24_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_25(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_26_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_25_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_25_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_25_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_25_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_26(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_27_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_26_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_26_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_26_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_26_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_27(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_28_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_27_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_27_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_27_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_27_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_28(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_29_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_28_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_28_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_28_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_28_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_29(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_30_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_29_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_29_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_29_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_29_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_30(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_31_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_30_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_30_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_30_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_30_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_31(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_32_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_31_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_31_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_31_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_31_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_32(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_33_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_32_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_32_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_32_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_32_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_33(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_34_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_33_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_33_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_33_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_33_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_33_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_34(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_35_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_34_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_34_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_34_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_34_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_34_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_35(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_36_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_35_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_35_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_35_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_35_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_35_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_36(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_37_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_36_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_36_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_36_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_36_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_36_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_37(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_38_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_37_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_37_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_37_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_37_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_37_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_38(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_39_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_38_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_38_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_38_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_38_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_38_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_39(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_40_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_39_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_39_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_39_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_39_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_39_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_40(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_41_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_40_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_40_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_40_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_40_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_40_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_41(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_42_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_41_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_41_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_41_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_41_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_41_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_42(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_43_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_42_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_42_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_42_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_42_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_42_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_43(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_44_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_43_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_43_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_43_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_43_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_43_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_44(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_45_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_44_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_44_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_44_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_44_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_44_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_45(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_46_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_45_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_45_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_45_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_45_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_45_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_46(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_47_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_46_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_46_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_46_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_46_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_46_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_47(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_48_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_47_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_47_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_47_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_47_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_47_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_48(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_49_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_48_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_48_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_48_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_48_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_48_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_49(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_50_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_49_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_49_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_49_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_49_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_49_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_50(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_51_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_50_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_50_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_50_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_50_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_50_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_51(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_52_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_51_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_51_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_51_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_51_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_51_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_52(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_53_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_52_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_52_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_52_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_52_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_52_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_53(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_54_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_53_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_53_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_53_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_53_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_53_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_54(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_55_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_54_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_54_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_54_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_54_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_54_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_55(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_56_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_55_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_55_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_55_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_55_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_55_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_56(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_57_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_56_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_56_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_56_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_56_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_56_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_57(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_58_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_57_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_57_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_57_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_57_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_57_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_58(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_59_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_58_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_58_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_58_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_58_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_58_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_59(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_60_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_59_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_59_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_59_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_59_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_59_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_60(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_61_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_60_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_60_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_60_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_60_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_60_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_61(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_62_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_61_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_61_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_61_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_61_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_61_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_62(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_63_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_62_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_62_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_62_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_62_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_62_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_63(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_64_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_63_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_63_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_63_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_63_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_63_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_64(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_65_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_64_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_64_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_64_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_64_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_64_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_65(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_66_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_65_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_65_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_65_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_65_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_65_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_66(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_67_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_66_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_66_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_66_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_66_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_66_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_67(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_68_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_67_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_67_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_67_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_67_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_67_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_68(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_69_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_68_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_68_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_68_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_68_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_68_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_69(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_70_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_69_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_69_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_69_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_69_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_69_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_70(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_71_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_70_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_70_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_70_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_70_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_70_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_71(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_72_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_71_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_71_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_71_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_71_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_71_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_72(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_73_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_72_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_72_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_72_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_72_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_72_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_73(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_74_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_73_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_73_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_73_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_73_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_73_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_74(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_75_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_74_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_74_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_74_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_74_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_74_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_75(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_76_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_75_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_75_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_75_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_75_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_75_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_76(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_77_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_76_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_76_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_76_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_76_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_76_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_77(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_78_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_77_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_77_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_77_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_77_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_77_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_78(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_79_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_78_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_78_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_78_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_78_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_78_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_79(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_80_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_79_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_79_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_79_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_79_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_79_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_80(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_81_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_80_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_80_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_80_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_80_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_80_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_81(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_0_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_81_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_81_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_81_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_81_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_81_ctrl_stealReq_ready)
	);
endmodule
module SchedulerClient_64 (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_ctrl_stealReq_valid,
	io_connNetwork_ctrl_stealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_connQ_currLength,
	io_connQ_push_ready,
	io_connQ_push_valid,
	io_connQ_push_bits,
	io_connQ_pop_ready,
	io_connQ_pop_valid,
	io_connQ_pop_bits
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_ctrl_stealReq_valid;
	input io_connNetwork_ctrl_stealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [255:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [255:0] io_connNetwork_data_qOutTask_bits;
	input [3:0] io_connQ_currLength;
	input io_connQ_push_ready;
	output wire io_connQ_push_valid;
	output wire [255:0] io_connQ_push_bits;
	output wire io_connQ_pop_ready;
	input io_connQ_pop_valid;
	input [255:0] io_connQ_pop_bits;
	reg [2:0] stateReg;
	reg [255:0] stolenTaskReg;
	reg [255:0] giveTaskReg;
	reg [31:0] requestKilledCount;
	reg [31:0] requestTaskCount;
	wire _GEN = stateReg == 3'h0;
	wire _GEN_0 = io_connQ_currLength < 4'h6;
	wire _GEN_1 = stateReg == 3'h2;
	wire _GEN_2 = requestKilledCount == 32'h00000000;
	wire _GEN_3 = stateReg == 3'h3;
	wire _GEN_4 = _GEN | _GEN_1;
	wire _GEN_5 = stateReg == 3'h4;
	wire _GEN_6 = io_connQ_currLength == 4'h0;
	wire _GEN_7 = stateReg == 3'h5;
	wire _GEN_8 = ((_GEN | _GEN_1) | _GEN_3) | _GEN_5;
	wire _GEN_9 = stateReg == 3'h6;
	wire io_connNetwork_ctrl_stealReq_valid_0 = ((|requestTaskCount & ~(_GEN_9 & _GEN_0)) & ~(_GEN_5 & _GEN_6)) & ~(_GEN_1 & _GEN_2);
	always @(posedge clock)
		if (reset) begin
			stateReg <= 3'h0;
			stolenTaskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			giveTaskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			requestKilledCount <= 32'h00000052;
			requestTaskCount <= 32'h00000000;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_10;
			reg _GEN_11;
			reg _GEN_12;
			reg _GEN_13;
			reg _GEN_14;
			reg _GEN_15;
			reg [23:0] _GEN_16;
			_GEN_10 = io_connQ_currLength > 4'h6;
			_GEN_11 = io_connQ_currLength > 4'h5;
			_GEN_12 = io_connQ_pop_valid | ~_GEN_6;
			_GEN_13 = io_connQ_currLength[3] | (io_connNetwork_ctrl_serveStealReq_ready & _GEN_11);
			_GEN_14 = _GEN_0 & io_connNetwork_ctrl_serveStealReq_ready;
			_GEN_15 = _GEN_14 | _GEN_0;
			_GEN_16 = {stateReg, (_GEN_13 ? 3'h4 : {~_GEN_15, 2'h2}), (io_connNetwork_data_qOutTask_ready ? 3'h0 : 3'h5), (io_connQ_pop_valid ? 3'h5 : (_GEN_6 ? 3'h2 : 3'h4)), (io_connQ_push_ready ? 3'h0 : (_GEN_10 ? 3'h5 : 3'h3)), (io_connNetwork_data_availableTask_valid ? 3'h3 : (_GEN_11 ? 3'h0 : (_GEN_2 ? stateReg : 3'h2))), stateReg, (_GEN_0 ? 3'h2 : (io_connQ_currLength[3] ? 3'h4 : (_GEN_10 ? 3'h6 : 3'h0)))};
			stateReg <= _GEN_16[stateReg * 3+:3];
			if (_GEN | ~(_GEN_1 & io_connNetwork_data_availableTask_valid))
				;
			else
				stolenTaskReg <= io_connNetwork_data_availableTask_bits;
			if (~_GEN_4) begin
				if (_GEN_3) begin
					if (io_connQ_push_ready | ~_GEN_10)
						;
					else
						giveTaskReg <= stolenTaskReg;
				end
				else if (_GEN_5 & io_connQ_pop_valid)
					giveTaskReg <= io_connQ_pop_bits;
			end
			if (_GEN) begin
				if (_GEN_0)
					requestKilledCount <= 32'h00000054;
			end
			else if (_GEN_1) begin
				if (io_connNetwork_ctrl_serveStealReq_ready)
					requestKilledCount <= 32'h00000054;
				else
					requestKilledCount <= requestKilledCount - 32'h00000001;
			end
			else if (_GEN_3 | (_GEN_5 ? _GEN_12 : ((_GEN_7 | ~_GEN_9) | _GEN_13) | ~_GEN_15))
				;
			else
				requestKilledCount <= 32'h00000054;
			if (io_connNetwork_ctrl_stealReq_valid_0 & io_connNetwork_ctrl_stealReq_ready)
				requestTaskCount <= requestTaskCount - 32'h00000001;
			else begin : sv2v_autoblock_2
				reg [31:0] _GEN_17;
				reg [255:0] _GEN_18;
				_GEN_17 = ((_GEN_7 | ~_GEN_9) | _GEN_13 ? requestTaskCount : (_GEN_14 ? requestTaskCount + 32'h00000002 : (_GEN_0 ? requestTaskCount + 32'h00000001 : requestTaskCount)));
				_GEN_18 = {_GEN_17, _GEN_17, requestTaskCount, (_GEN_12 ? requestTaskCount : requestTaskCount + 32'h00000001), requestTaskCount, ((io_connNetwork_data_availableTask_valid | _GEN_11) | ~_GEN_2 ? requestTaskCount : requestTaskCount + 32'h00000001), _GEN_17, (_GEN_0 ? requestTaskCount + 32'h00000001 : requestTaskCount)};
				requestTaskCount <= _GEN_18[stateReg * 32+:32];
			end
		end
	assign io_connNetwork_ctrl_serveStealReq_valid = ~((((_GEN | _GEN_1) | _GEN_3) | _GEN_5) | _GEN_7) & _GEN_9;
	assign io_connNetwork_ctrl_stealReq_valid = io_connNetwork_ctrl_stealReq_valid_0;
	assign io_connNetwork_data_availableTask_ready = ~_GEN & _GEN_1;
	assign io_connNetwork_data_qOutTask_valid = ~_GEN_8 & _GEN_7;
	assign io_connNetwork_data_qOutTask_bits = (_GEN_8 | ~_GEN_7 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : giveTaskReg);
	assign io_connQ_push_valid = ~_GEN_4 & _GEN_3;
	assign io_connQ_push_bits = (_GEN_4 | ~_GEN_3 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : stolenTaskReg);
	assign io_connQ_pop_ready = ~((_GEN | _GEN_1) | _GEN_3) & _GEN_5;
endmodule
module hw_deque_64 (
	clock,
	reset,
	io_connVec_0_pop_ready,
	io_connVec_0_pop_valid,
	io_connVec_0_pop_bits,
	io_connVec_1_currLength,
	io_connVec_1_push_ready,
	io_connVec_1_push_valid,
	io_connVec_1_push_bits,
	io_connVec_1_pop_ready,
	io_connVec_1_pop_valid,
	io_connVec_1_pop_bits
);
	input clock;
	input reset;
	input io_connVec_0_pop_ready;
	output wire io_connVec_0_pop_valid;
	output wire [255:0] io_connVec_0_pop_bits;
	output wire [4:0] io_connVec_1_currLength;
	output wire io_connVec_1_push_ready;
	input io_connVec_1_push_valid;
	input [255:0] io_connVec_1_push_bits;
	input io_connVec_1_pop_ready;
	output wire io_connVec_1_pop_valid;
	output wire [255:0] io_connVec_1_pop_bits;
	wire [255:0] _bramMem_a_dout;
	wire [255:0] _bramMem_b_dout;
	reg [4:0] sideReg_0;
	reg [4:0] sideReg_1;
	reg readLatency_0;
	reg readLatency_1;
	reg writeLatency_0;
	reg writeLatency_1;
	reg [2:0] stateRegs_0;
	reg [2:0] stateRegs_1;
	wire _GEN = stateRegs_0 == 3'h0;
	wire _GEN_0 = stateRegs_1 == 3'h0;
	wire _GEN_1 = stateRegs_0 == 3'h1;
	wire _GEN_2 = stateRegs_0 == 3'h2;
	wire _GEN_3 = sideReg_0 == 5'h09;
	wire _GEN_4 = stateRegs_0 == 3'h4;
	wire [4:0] _bramMem_io_a_addr_T_2 = sideReg_0 + 5'h01;
	wire _GEN_5 = (_GEN | _GEN_1) | _GEN_2;
	wire _GEN_6 = stateRegs_1 == 3'h1;
	wire _GEN_7 = stateRegs_1 == 3'h2;
	wire _GEN_8 = sideReg_1 == 5'h00;
	wire _GEN_9 = stateRegs_1 == 3'h4;
	wire [4:0] _bramMem_io_b_addr_T_6 = sideReg_1 - 5'h01;
	wire _GEN_10 = (_GEN_0 | _GEN_6) | _GEN_7;
	wire _GEN_11 = stateRegs_1 == 3'h3;
	wire [4:0] currLen = (sideReg_0 > sideReg_1 ? ((sideReg_1 + 5'h0a) - sideReg_0) - 5'h01 : (sideReg_1 - sideReg_0) - 5'h01);
	always @(posedge clock)
		if (reset) begin
			sideReg_0 <= 5'h00;
			sideReg_1 <= 5'h01;
			readLatency_0 <= 1'h0;
			readLatency_1 <= 1'h0;
			writeLatency_0 <= 1'h0;
			writeLatency_1 <= 1'h0;
			stateRegs_0 <= 3'h0;
			stateRegs_1 <= 3'h0;
		end
		else begin : sv2v_autoblock_1
			reg [23:0] _GEN_12;
			reg [23:0] _GEN_13;
			_GEN_12 = {stateRegs_0, stateRegs_0, stateRegs_0, 6'h00, (readLatency_0 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_0, 2'h2, (io_connVec_0_pop_ready & |currLen[4:1]) | ((io_connVec_0_pop_ready & _GEN_0) & |currLen), 1'h0};
			_GEN_13 = {stateRegs_1, stateRegs_1, stateRegs_1, 6'h00, (readLatency_1 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_1, 1'h1, (io_connVec_1_push_valid & (currLen < 5'h09) ? 3'h1 : {1'h0, (io_connVec_1_pop_ready & |currLen[4:1]) | (((io_connVec_1_pop_ready & ~io_connVec_0_pop_ready) & |currLen) & (stateRegs_0 != 3'h4)), 1'h0})};
			if (~_GEN_5) begin
				if (_GEN_4) begin
					if (_GEN_3)
						sideReg_0 <= 5'h00;
					else
						sideReg_0 <= _bramMem_io_a_addr_T_2;
				end
				else if (stateRegs_0 == 3'h3) begin
					if (sideReg_0 == 5'h00)
						sideReg_0 <= 5'h09;
					else
						sideReg_0 <= sideReg_0 - 5'h01;
				end
			end
			if (~_GEN_10) begin
				if (_GEN_9) begin
					if (_GEN_8)
						sideReg_1 <= 5'h09;
					else
						sideReg_1 <= _bramMem_io_b_addr_T_6;
				end
				else if (_GEN_11) begin
					if (sideReg_1 == 5'h09)
						sideReg_1 <= 5'h00;
					else
						sideReg_1 <= sideReg_1 + 5'h01;
				end
			end
			readLatency_0 <= (((_GEN | _GEN_1) | ~_GEN_2) | (readLatency_0 - 1'h1)) & readLatency_0;
			readLatency_1 <= (((_GEN_0 | _GEN_6) | ~_GEN_7) | (readLatency_1 - 1'h1)) & readLatency_1;
			writeLatency_0 <= ((_GEN | ~_GEN_1) | (writeLatency_0 - 1'h1)) & writeLatency_0;
			writeLatency_1 <= ((_GEN_0 | ~_GEN_6) | (writeLatency_1 - 1'h1)) & writeLatency_1;
			stateRegs_0 <= _GEN_12[stateRegs_0 * 3+:3];
			stateRegs_1 <= _GEN_13[stateRegs_1 * 3+:3];
		end
	DualPortBRAM #(
		.ADDR(7),
		.DATA(256)
	) bramMem(
		.clk(clock),
		.rst(reset),
		.a_addr((_GEN ? 7'h7f : (_GEN_1 ? {2'h0, sideReg_0} : (_GEN_2 ? (_GEN_3 ? 7'h00 : {2'h0, sideReg_0 + 5'h01}) : (_GEN_4 ? (_GEN_3 ? 7'h00 : {2'h0, _bramMem_io_a_addr_T_2}) : 7'h7f))))),
		.a_din(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.a_wr(~_GEN & _GEN_1),
		.a_dout(_bramMem_a_dout),
		.b_addr((_GEN_0 ? 7'h7f : (_GEN_6 ? {2'h0, sideReg_1} : (_GEN_7 ? (_GEN_8 ? 7'h09 : {2'h0, sideReg_1 - 5'h01}) : (_GEN_9 ? (_GEN_8 ? 7'h09 : {2'h0, _bramMem_io_b_addr_T_6}) : 7'h7f))))),
		.b_din(io_connVec_1_push_bits),
		.b_wr(~_GEN_0 & _GEN_6),
		.b_dout(_bramMem_b_dout)
	);
	assign io_connVec_0_pop_valid = ~_GEN_5 & _GEN_4;
	assign io_connVec_0_pop_bits = (_GEN_5 | ~_GEN_4 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : _bramMem_a_dout);
	assign io_connVec_1_currLength = currLen;
	assign io_connVec_1_push_ready = ~(((_GEN_0 | _GEN_6) | _GEN_7) | _GEN_9) & _GEN_11;
	assign io_connVec_1_pop_valid = ~_GEN_10 & _GEN_9;
	assign io_connVec_1_pop_bits = (_GEN_10 | ~_GEN_9 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : _bramMem_b_dout);
endmodule
module SchedulerLocalNetwork_1 (
	clock,
	reset,
	io_connPE_0_pop_ready,
	io_connPE_0_pop_valid,
	io_connPE_0_pop_bits,
	io_connPE_1_pop_ready,
	io_connPE_1_pop_valid,
	io_connPE_1_pop_bits,
	io_connPE_2_pop_ready,
	io_connPE_2_pop_valid,
	io_connPE_2_pop_bits,
	io_connPE_3_pop_ready,
	io_connPE_3_pop_valid,
	io_connPE_3_pop_bits,
	io_connPE_4_pop_ready,
	io_connPE_4_pop_valid,
	io_connPE_4_pop_bits,
	io_connPE_5_pop_ready,
	io_connPE_5_pop_valid,
	io_connPE_5_pop_bits,
	io_connPE_6_pop_ready,
	io_connPE_6_pop_valid,
	io_connPE_6_pop_bits,
	io_connPE_7_pop_ready,
	io_connPE_7_pop_valid,
	io_connPE_7_pop_bits,
	io_connPE_8_pop_ready,
	io_connPE_8_pop_valid,
	io_connPE_8_pop_bits,
	io_connPE_9_pop_ready,
	io_connPE_9_pop_valid,
	io_connPE_9_pop_bits,
	io_connPE_10_pop_ready,
	io_connPE_10_pop_valid,
	io_connPE_10_pop_bits,
	io_connPE_11_pop_ready,
	io_connPE_11_pop_valid,
	io_connPE_11_pop_bits,
	io_connPE_12_pop_ready,
	io_connPE_12_pop_valid,
	io_connPE_12_pop_bits,
	io_connPE_13_pop_ready,
	io_connPE_13_pop_valid,
	io_connPE_13_pop_bits,
	io_connPE_14_pop_ready,
	io_connPE_14_pop_valid,
	io_connPE_14_pop_bits,
	io_connPE_15_pop_ready,
	io_connPE_15_pop_valid,
	io_connPE_15_pop_bits,
	io_connPE_16_pop_ready,
	io_connPE_16_pop_valid,
	io_connPE_16_pop_bits,
	io_connPE_17_pop_ready,
	io_connPE_17_pop_valid,
	io_connPE_17_pop_bits,
	io_connPE_18_pop_ready,
	io_connPE_18_pop_valid,
	io_connPE_18_pop_bits,
	io_connPE_19_pop_ready,
	io_connPE_19_pop_valid,
	io_connPE_19_pop_bits,
	io_connPE_20_pop_ready,
	io_connPE_20_pop_valid,
	io_connPE_20_pop_bits,
	io_connPE_21_pop_ready,
	io_connPE_21_pop_valid,
	io_connPE_21_pop_bits,
	io_connPE_22_pop_ready,
	io_connPE_22_pop_valid,
	io_connPE_22_pop_bits,
	io_connPE_23_pop_ready,
	io_connPE_23_pop_valid,
	io_connPE_23_pop_bits,
	io_connPE_24_pop_ready,
	io_connPE_24_pop_valid,
	io_connPE_24_pop_bits,
	io_connPE_25_pop_ready,
	io_connPE_25_pop_valid,
	io_connPE_25_pop_bits,
	io_connPE_26_pop_ready,
	io_connPE_26_pop_valid,
	io_connPE_26_pop_bits,
	io_connPE_27_pop_ready,
	io_connPE_27_pop_valid,
	io_connPE_27_pop_bits,
	io_connPE_28_pop_ready,
	io_connPE_28_pop_valid,
	io_connPE_28_pop_bits,
	io_connPE_29_pop_ready,
	io_connPE_29_pop_valid,
	io_connPE_29_pop_bits,
	io_connPE_30_pop_ready,
	io_connPE_30_pop_valid,
	io_connPE_30_pop_bits,
	io_connPE_31_pop_ready,
	io_connPE_31_pop_valid,
	io_connPE_31_pop_bits,
	io_connPE_32_pop_ready,
	io_connPE_32_pop_valid,
	io_connPE_32_pop_bits,
	io_connPE_33_pop_ready,
	io_connPE_33_pop_valid,
	io_connPE_33_pop_bits,
	io_connPE_34_pop_ready,
	io_connPE_34_pop_valid,
	io_connPE_34_pop_bits,
	io_connPE_35_pop_ready,
	io_connPE_35_pop_valid,
	io_connPE_35_pop_bits,
	io_connPE_36_pop_ready,
	io_connPE_36_pop_valid,
	io_connPE_36_pop_bits,
	io_connPE_37_pop_ready,
	io_connPE_37_pop_valid,
	io_connPE_37_pop_bits,
	io_connPE_38_pop_ready,
	io_connPE_38_pop_valid,
	io_connPE_38_pop_bits,
	io_connPE_39_pop_ready,
	io_connPE_39_pop_valid,
	io_connPE_39_pop_bits,
	io_connPE_40_pop_ready,
	io_connPE_40_pop_valid,
	io_connPE_40_pop_bits,
	io_connPE_41_pop_ready,
	io_connPE_41_pop_valid,
	io_connPE_41_pop_bits,
	io_connPE_42_pop_ready,
	io_connPE_42_pop_valid,
	io_connPE_42_pop_bits,
	io_connPE_43_pop_ready,
	io_connPE_43_pop_valid,
	io_connPE_43_pop_bits,
	io_connPE_44_pop_ready,
	io_connPE_44_pop_valid,
	io_connPE_44_pop_bits,
	io_connPE_45_pop_ready,
	io_connPE_45_pop_valid,
	io_connPE_45_pop_bits,
	io_connPE_46_pop_ready,
	io_connPE_46_pop_valid,
	io_connPE_46_pop_bits,
	io_connPE_47_pop_ready,
	io_connPE_47_pop_valid,
	io_connPE_47_pop_bits,
	io_connPE_48_pop_ready,
	io_connPE_48_pop_valid,
	io_connPE_48_pop_bits,
	io_connPE_49_pop_ready,
	io_connPE_49_pop_valid,
	io_connPE_49_pop_bits,
	io_connPE_50_pop_ready,
	io_connPE_50_pop_valid,
	io_connPE_50_pop_bits,
	io_connPE_51_pop_ready,
	io_connPE_51_pop_valid,
	io_connPE_51_pop_bits,
	io_connPE_52_pop_ready,
	io_connPE_52_pop_valid,
	io_connPE_52_pop_bits,
	io_connPE_53_pop_ready,
	io_connPE_53_pop_valid,
	io_connPE_53_pop_bits,
	io_connPE_54_pop_ready,
	io_connPE_54_pop_valid,
	io_connPE_54_pop_bits,
	io_connPE_55_pop_ready,
	io_connPE_55_pop_valid,
	io_connPE_55_pop_bits,
	io_connPE_56_pop_ready,
	io_connPE_56_pop_valid,
	io_connPE_56_pop_bits,
	io_connPE_57_pop_ready,
	io_connPE_57_pop_valid,
	io_connPE_57_pop_bits,
	io_connPE_58_pop_ready,
	io_connPE_58_pop_valid,
	io_connPE_58_pop_bits,
	io_connPE_59_pop_ready,
	io_connPE_59_pop_valid,
	io_connPE_59_pop_bits,
	io_connPE_60_pop_ready,
	io_connPE_60_pop_valid,
	io_connPE_60_pop_bits,
	io_connPE_61_pop_ready,
	io_connPE_61_pop_valid,
	io_connPE_61_pop_bits,
	io_connPE_62_pop_ready,
	io_connPE_62_pop_valid,
	io_connPE_62_pop_bits,
	io_connPE_63_pop_ready,
	io_connPE_63_pop_valid,
	io_connPE_63_pop_bits,
	io_connVSS_0_ctrl_serveStealReq_valid,
	io_connVSS_0_ctrl_serveStealReq_ready,
	io_connVSS_0_data_availableTask_ready,
	io_connVSS_0_data_availableTask_valid,
	io_connVSS_0_data_availableTask_bits,
	io_connVSS_0_data_qOutTask_ready,
	io_connVSS_0_data_qOutTask_valid,
	io_connVSS_0_data_qOutTask_bits,
	io_connVSS_1_ctrl_serveStealReq_valid,
	io_connVSS_1_ctrl_serveStealReq_ready,
	io_connVSS_1_data_availableTask_ready,
	io_connVSS_1_data_availableTask_valid,
	io_connVSS_1_data_availableTask_bits,
	io_connVSS_1_data_qOutTask_ready,
	io_connVSS_1_data_qOutTask_valid,
	io_connVSS_1_data_qOutTask_bits,
	io_connVAS_0_ctrl_serveStealReq_valid,
	io_connVAS_0_ctrl_serveStealReq_ready,
	io_connVAS_0_data_qOutTask_ready,
	io_connVAS_0_data_qOutTask_valid,
	io_connVAS_0_data_qOutTask_bits,
	io_connVAS_1_ctrl_serveStealReq_valid,
	io_connVAS_1_ctrl_serveStealReq_ready,
	io_connVAS_1_data_qOutTask_ready,
	io_connVAS_1_data_qOutTask_valid,
	io_connVAS_1_data_qOutTask_bits,
	io_connVAS_2_ctrl_serveStealReq_valid,
	io_connVAS_2_ctrl_serveStealReq_ready,
	io_connVAS_2_data_qOutTask_ready,
	io_connVAS_2_data_qOutTask_valid,
	io_connVAS_2_data_qOutTask_bits,
	io_connVAS_3_ctrl_serveStealReq_valid,
	io_connVAS_3_ctrl_serveStealReq_ready,
	io_connVAS_3_data_qOutTask_ready,
	io_connVAS_3_data_qOutTask_valid,
	io_connVAS_3_data_qOutTask_bits,
	io_connVAS_4_ctrl_serveStealReq_valid,
	io_connVAS_4_ctrl_serveStealReq_ready,
	io_connVAS_4_data_qOutTask_ready,
	io_connVAS_4_data_qOutTask_valid,
	io_connVAS_4_data_qOutTask_bits,
	io_connVAS_5_ctrl_serveStealReq_valid,
	io_connVAS_5_ctrl_serveStealReq_ready,
	io_connVAS_5_data_qOutTask_ready,
	io_connVAS_5_data_qOutTask_valid,
	io_connVAS_5_data_qOutTask_bits,
	io_connVAS_6_ctrl_serveStealReq_valid,
	io_connVAS_6_ctrl_serveStealReq_ready,
	io_connVAS_6_data_qOutTask_ready,
	io_connVAS_6_data_qOutTask_valid,
	io_connVAS_6_data_qOutTask_bits,
	io_connVAS_7_ctrl_serveStealReq_valid,
	io_connVAS_7_ctrl_serveStealReq_ready,
	io_connVAS_7_data_qOutTask_ready,
	io_connVAS_7_data_qOutTask_valid,
	io_connVAS_7_data_qOutTask_bits,
	io_connVAS_8_ctrl_serveStealReq_valid,
	io_connVAS_8_ctrl_serveStealReq_ready,
	io_connVAS_8_data_qOutTask_ready,
	io_connVAS_8_data_qOutTask_valid,
	io_connVAS_8_data_qOutTask_bits,
	io_connVAS_9_ctrl_serveStealReq_valid,
	io_connVAS_9_ctrl_serveStealReq_ready,
	io_connVAS_9_data_qOutTask_ready,
	io_connVAS_9_data_qOutTask_valid,
	io_connVAS_9_data_qOutTask_bits,
	io_connVAS_10_ctrl_serveStealReq_valid,
	io_connVAS_10_ctrl_serveStealReq_ready,
	io_connVAS_10_data_qOutTask_ready,
	io_connVAS_10_data_qOutTask_valid,
	io_connVAS_10_data_qOutTask_bits,
	io_connVAS_11_ctrl_serveStealReq_valid,
	io_connVAS_11_ctrl_serveStealReq_ready,
	io_connVAS_11_data_qOutTask_ready,
	io_connVAS_11_data_qOutTask_valid,
	io_connVAS_11_data_qOutTask_bits,
	io_connVAS_12_ctrl_serveStealReq_valid,
	io_connVAS_12_ctrl_serveStealReq_ready,
	io_connVAS_12_data_qOutTask_ready,
	io_connVAS_12_data_qOutTask_valid,
	io_connVAS_12_data_qOutTask_bits,
	io_connVAS_13_ctrl_serveStealReq_valid,
	io_connVAS_13_ctrl_serveStealReq_ready,
	io_connVAS_13_data_qOutTask_ready,
	io_connVAS_13_data_qOutTask_valid,
	io_connVAS_13_data_qOutTask_bits,
	io_connVAS_14_ctrl_serveStealReq_valid,
	io_connVAS_14_ctrl_serveStealReq_ready,
	io_connVAS_14_data_qOutTask_ready,
	io_connVAS_14_data_qOutTask_valid,
	io_connVAS_14_data_qOutTask_bits,
	io_connVAS_15_ctrl_serveStealReq_valid,
	io_connVAS_15_ctrl_serveStealReq_ready,
	io_connVAS_15_data_qOutTask_ready,
	io_connVAS_15_data_qOutTask_valid,
	io_connVAS_15_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0,
	io_ntwDataUnitOccupancyVSS_1
);
	input clock;
	input reset;
	input io_connPE_0_pop_ready;
	output wire io_connPE_0_pop_valid;
	output wire [255:0] io_connPE_0_pop_bits;
	input io_connPE_1_pop_ready;
	output wire io_connPE_1_pop_valid;
	output wire [255:0] io_connPE_1_pop_bits;
	input io_connPE_2_pop_ready;
	output wire io_connPE_2_pop_valid;
	output wire [255:0] io_connPE_2_pop_bits;
	input io_connPE_3_pop_ready;
	output wire io_connPE_3_pop_valid;
	output wire [255:0] io_connPE_3_pop_bits;
	input io_connPE_4_pop_ready;
	output wire io_connPE_4_pop_valid;
	output wire [255:0] io_connPE_4_pop_bits;
	input io_connPE_5_pop_ready;
	output wire io_connPE_5_pop_valid;
	output wire [255:0] io_connPE_5_pop_bits;
	input io_connPE_6_pop_ready;
	output wire io_connPE_6_pop_valid;
	output wire [255:0] io_connPE_6_pop_bits;
	input io_connPE_7_pop_ready;
	output wire io_connPE_7_pop_valid;
	output wire [255:0] io_connPE_7_pop_bits;
	input io_connPE_8_pop_ready;
	output wire io_connPE_8_pop_valid;
	output wire [255:0] io_connPE_8_pop_bits;
	input io_connPE_9_pop_ready;
	output wire io_connPE_9_pop_valid;
	output wire [255:0] io_connPE_9_pop_bits;
	input io_connPE_10_pop_ready;
	output wire io_connPE_10_pop_valid;
	output wire [255:0] io_connPE_10_pop_bits;
	input io_connPE_11_pop_ready;
	output wire io_connPE_11_pop_valid;
	output wire [255:0] io_connPE_11_pop_bits;
	input io_connPE_12_pop_ready;
	output wire io_connPE_12_pop_valid;
	output wire [255:0] io_connPE_12_pop_bits;
	input io_connPE_13_pop_ready;
	output wire io_connPE_13_pop_valid;
	output wire [255:0] io_connPE_13_pop_bits;
	input io_connPE_14_pop_ready;
	output wire io_connPE_14_pop_valid;
	output wire [255:0] io_connPE_14_pop_bits;
	input io_connPE_15_pop_ready;
	output wire io_connPE_15_pop_valid;
	output wire [255:0] io_connPE_15_pop_bits;
	input io_connPE_16_pop_ready;
	output wire io_connPE_16_pop_valid;
	output wire [255:0] io_connPE_16_pop_bits;
	input io_connPE_17_pop_ready;
	output wire io_connPE_17_pop_valid;
	output wire [255:0] io_connPE_17_pop_bits;
	input io_connPE_18_pop_ready;
	output wire io_connPE_18_pop_valid;
	output wire [255:0] io_connPE_18_pop_bits;
	input io_connPE_19_pop_ready;
	output wire io_connPE_19_pop_valid;
	output wire [255:0] io_connPE_19_pop_bits;
	input io_connPE_20_pop_ready;
	output wire io_connPE_20_pop_valid;
	output wire [255:0] io_connPE_20_pop_bits;
	input io_connPE_21_pop_ready;
	output wire io_connPE_21_pop_valid;
	output wire [255:0] io_connPE_21_pop_bits;
	input io_connPE_22_pop_ready;
	output wire io_connPE_22_pop_valid;
	output wire [255:0] io_connPE_22_pop_bits;
	input io_connPE_23_pop_ready;
	output wire io_connPE_23_pop_valid;
	output wire [255:0] io_connPE_23_pop_bits;
	input io_connPE_24_pop_ready;
	output wire io_connPE_24_pop_valid;
	output wire [255:0] io_connPE_24_pop_bits;
	input io_connPE_25_pop_ready;
	output wire io_connPE_25_pop_valid;
	output wire [255:0] io_connPE_25_pop_bits;
	input io_connPE_26_pop_ready;
	output wire io_connPE_26_pop_valid;
	output wire [255:0] io_connPE_26_pop_bits;
	input io_connPE_27_pop_ready;
	output wire io_connPE_27_pop_valid;
	output wire [255:0] io_connPE_27_pop_bits;
	input io_connPE_28_pop_ready;
	output wire io_connPE_28_pop_valid;
	output wire [255:0] io_connPE_28_pop_bits;
	input io_connPE_29_pop_ready;
	output wire io_connPE_29_pop_valid;
	output wire [255:0] io_connPE_29_pop_bits;
	input io_connPE_30_pop_ready;
	output wire io_connPE_30_pop_valid;
	output wire [255:0] io_connPE_30_pop_bits;
	input io_connPE_31_pop_ready;
	output wire io_connPE_31_pop_valid;
	output wire [255:0] io_connPE_31_pop_bits;
	input io_connPE_32_pop_ready;
	output wire io_connPE_32_pop_valid;
	output wire [255:0] io_connPE_32_pop_bits;
	input io_connPE_33_pop_ready;
	output wire io_connPE_33_pop_valid;
	output wire [255:0] io_connPE_33_pop_bits;
	input io_connPE_34_pop_ready;
	output wire io_connPE_34_pop_valid;
	output wire [255:0] io_connPE_34_pop_bits;
	input io_connPE_35_pop_ready;
	output wire io_connPE_35_pop_valid;
	output wire [255:0] io_connPE_35_pop_bits;
	input io_connPE_36_pop_ready;
	output wire io_connPE_36_pop_valid;
	output wire [255:0] io_connPE_36_pop_bits;
	input io_connPE_37_pop_ready;
	output wire io_connPE_37_pop_valid;
	output wire [255:0] io_connPE_37_pop_bits;
	input io_connPE_38_pop_ready;
	output wire io_connPE_38_pop_valid;
	output wire [255:0] io_connPE_38_pop_bits;
	input io_connPE_39_pop_ready;
	output wire io_connPE_39_pop_valid;
	output wire [255:0] io_connPE_39_pop_bits;
	input io_connPE_40_pop_ready;
	output wire io_connPE_40_pop_valid;
	output wire [255:0] io_connPE_40_pop_bits;
	input io_connPE_41_pop_ready;
	output wire io_connPE_41_pop_valid;
	output wire [255:0] io_connPE_41_pop_bits;
	input io_connPE_42_pop_ready;
	output wire io_connPE_42_pop_valid;
	output wire [255:0] io_connPE_42_pop_bits;
	input io_connPE_43_pop_ready;
	output wire io_connPE_43_pop_valid;
	output wire [255:0] io_connPE_43_pop_bits;
	input io_connPE_44_pop_ready;
	output wire io_connPE_44_pop_valid;
	output wire [255:0] io_connPE_44_pop_bits;
	input io_connPE_45_pop_ready;
	output wire io_connPE_45_pop_valid;
	output wire [255:0] io_connPE_45_pop_bits;
	input io_connPE_46_pop_ready;
	output wire io_connPE_46_pop_valid;
	output wire [255:0] io_connPE_46_pop_bits;
	input io_connPE_47_pop_ready;
	output wire io_connPE_47_pop_valid;
	output wire [255:0] io_connPE_47_pop_bits;
	input io_connPE_48_pop_ready;
	output wire io_connPE_48_pop_valid;
	output wire [255:0] io_connPE_48_pop_bits;
	input io_connPE_49_pop_ready;
	output wire io_connPE_49_pop_valid;
	output wire [255:0] io_connPE_49_pop_bits;
	input io_connPE_50_pop_ready;
	output wire io_connPE_50_pop_valid;
	output wire [255:0] io_connPE_50_pop_bits;
	input io_connPE_51_pop_ready;
	output wire io_connPE_51_pop_valid;
	output wire [255:0] io_connPE_51_pop_bits;
	input io_connPE_52_pop_ready;
	output wire io_connPE_52_pop_valid;
	output wire [255:0] io_connPE_52_pop_bits;
	input io_connPE_53_pop_ready;
	output wire io_connPE_53_pop_valid;
	output wire [255:0] io_connPE_53_pop_bits;
	input io_connPE_54_pop_ready;
	output wire io_connPE_54_pop_valid;
	output wire [255:0] io_connPE_54_pop_bits;
	input io_connPE_55_pop_ready;
	output wire io_connPE_55_pop_valid;
	output wire [255:0] io_connPE_55_pop_bits;
	input io_connPE_56_pop_ready;
	output wire io_connPE_56_pop_valid;
	output wire [255:0] io_connPE_56_pop_bits;
	input io_connPE_57_pop_ready;
	output wire io_connPE_57_pop_valid;
	output wire [255:0] io_connPE_57_pop_bits;
	input io_connPE_58_pop_ready;
	output wire io_connPE_58_pop_valid;
	output wire [255:0] io_connPE_58_pop_bits;
	input io_connPE_59_pop_ready;
	output wire io_connPE_59_pop_valid;
	output wire [255:0] io_connPE_59_pop_bits;
	input io_connPE_60_pop_ready;
	output wire io_connPE_60_pop_valid;
	output wire [255:0] io_connPE_60_pop_bits;
	input io_connPE_61_pop_ready;
	output wire io_connPE_61_pop_valid;
	output wire [255:0] io_connPE_61_pop_bits;
	input io_connPE_62_pop_ready;
	output wire io_connPE_62_pop_valid;
	output wire [255:0] io_connPE_62_pop_bits;
	input io_connPE_63_pop_ready;
	output wire io_connPE_63_pop_valid;
	output wire [255:0] io_connPE_63_pop_bits;
	input io_connVSS_0_ctrl_serveStealReq_valid;
	output wire io_connVSS_0_ctrl_serveStealReq_ready;
	input io_connVSS_0_data_availableTask_ready;
	output wire io_connVSS_0_data_availableTask_valid;
	output wire [255:0] io_connVSS_0_data_availableTask_bits;
	output wire io_connVSS_0_data_qOutTask_ready;
	input io_connVSS_0_data_qOutTask_valid;
	input [255:0] io_connVSS_0_data_qOutTask_bits;
	input io_connVSS_1_ctrl_serveStealReq_valid;
	output wire io_connVSS_1_ctrl_serveStealReq_ready;
	input io_connVSS_1_data_availableTask_ready;
	output wire io_connVSS_1_data_availableTask_valid;
	output wire [255:0] io_connVSS_1_data_availableTask_bits;
	output wire io_connVSS_1_data_qOutTask_ready;
	input io_connVSS_1_data_qOutTask_valid;
	input [255:0] io_connVSS_1_data_qOutTask_bits;
	input io_connVAS_0_ctrl_serveStealReq_valid;
	output wire io_connVAS_0_ctrl_serveStealReq_ready;
	output wire io_connVAS_0_data_qOutTask_ready;
	input io_connVAS_0_data_qOutTask_valid;
	input [255:0] io_connVAS_0_data_qOutTask_bits;
	input io_connVAS_1_ctrl_serveStealReq_valid;
	output wire io_connVAS_1_ctrl_serveStealReq_ready;
	output wire io_connVAS_1_data_qOutTask_ready;
	input io_connVAS_1_data_qOutTask_valid;
	input [255:0] io_connVAS_1_data_qOutTask_bits;
	input io_connVAS_2_ctrl_serveStealReq_valid;
	output wire io_connVAS_2_ctrl_serveStealReq_ready;
	output wire io_connVAS_2_data_qOutTask_ready;
	input io_connVAS_2_data_qOutTask_valid;
	input [255:0] io_connVAS_2_data_qOutTask_bits;
	input io_connVAS_3_ctrl_serveStealReq_valid;
	output wire io_connVAS_3_ctrl_serveStealReq_ready;
	output wire io_connVAS_3_data_qOutTask_ready;
	input io_connVAS_3_data_qOutTask_valid;
	input [255:0] io_connVAS_3_data_qOutTask_bits;
	input io_connVAS_4_ctrl_serveStealReq_valid;
	output wire io_connVAS_4_ctrl_serveStealReq_ready;
	output wire io_connVAS_4_data_qOutTask_ready;
	input io_connVAS_4_data_qOutTask_valid;
	input [255:0] io_connVAS_4_data_qOutTask_bits;
	input io_connVAS_5_ctrl_serveStealReq_valid;
	output wire io_connVAS_5_ctrl_serveStealReq_ready;
	output wire io_connVAS_5_data_qOutTask_ready;
	input io_connVAS_5_data_qOutTask_valid;
	input [255:0] io_connVAS_5_data_qOutTask_bits;
	input io_connVAS_6_ctrl_serveStealReq_valid;
	output wire io_connVAS_6_ctrl_serveStealReq_ready;
	output wire io_connVAS_6_data_qOutTask_ready;
	input io_connVAS_6_data_qOutTask_valid;
	input [255:0] io_connVAS_6_data_qOutTask_bits;
	input io_connVAS_7_ctrl_serveStealReq_valid;
	output wire io_connVAS_7_ctrl_serveStealReq_ready;
	output wire io_connVAS_7_data_qOutTask_ready;
	input io_connVAS_7_data_qOutTask_valid;
	input [255:0] io_connVAS_7_data_qOutTask_bits;
	input io_connVAS_8_ctrl_serveStealReq_valid;
	output wire io_connVAS_8_ctrl_serveStealReq_ready;
	output wire io_connVAS_8_data_qOutTask_ready;
	input io_connVAS_8_data_qOutTask_valid;
	input [255:0] io_connVAS_8_data_qOutTask_bits;
	input io_connVAS_9_ctrl_serveStealReq_valid;
	output wire io_connVAS_9_ctrl_serveStealReq_ready;
	output wire io_connVAS_9_data_qOutTask_ready;
	input io_connVAS_9_data_qOutTask_valid;
	input [255:0] io_connVAS_9_data_qOutTask_bits;
	input io_connVAS_10_ctrl_serveStealReq_valid;
	output wire io_connVAS_10_ctrl_serveStealReq_ready;
	output wire io_connVAS_10_data_qOutTask_ready;
	input io_connVAS_10_data_qOutTask_valid;
	input [255:0] io_connVAS_10_data_qOutTask_bits;
	input io_connVAS_11_ctrl_serveStealReq_valid;
	output wire io_connVAS_11_ctrl_serveStealReq_ready;
	output wire io_connVAS_11_data_qOutTask_ready;
	input io_connVAS_11_data_qOutTask_valid;
	input [255:0] io_connVAS_11_data_qOutTask_bits;
	input io_connVAS_12_ctrl_serveStealReq_valid;
	output wire io_connVAS_12_ctrl_serveStealReq_ready;
	output wire io_connVAS_12_data_qOutTask_ready;
	input io_connVAS_12_data_qOutTask_valid;
	input [255:0] io_connVAS_12_data_qOutTask_bits;
	input io_connVAS_13_ctrl_serveStealReq_valid;
	output wire io_connVAS_13_ctrl_serveStealReq_ready;
	output wire io_connVAS_13_data_qOutTask_ready;
	input io_connVAS_13_data_qOutTask_valid;
	input [255:0] io_connVAS_13_data_qOutTask_bits;
	input io_connVAS_14_ctrl_serveStealReq_valid;
	output wire io_connVAS_14_ctrl_serveStealReq_ready;
	output wire io_connVAS_14_data_qOutTask_ready;
	input io_connVAS_14_data_qOutTask_valid;
	input [255:0] io_connVAS_14_data_qOutTask_bits;
	input io_connVAS_15_ctrl_serveStealReq_valid;
	output wire io_connVAS_15_ctrl_serveStealReq_ready;
	output wire io_connVAS_15_data_qOutTask_ready;
	input io_connVAS_15_data_qOutTask_valid;
	input [255:0] io_connVAS_15_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	output wire io_ntwDataUnitOccupancyVSS_1;
	wire [4:0] _taskQueues_63_io_connVec_1_currLength;
	wire _taskQueues_63_io_connVec_1_push_ready;
	wire _taskQueues_63_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_63_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_62_io_connVec_1_currLength;
	wire _taskQueues_62_io_connVec_1_push_ready;
	wire _taskQueues_62_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_62_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_61_io_connVec_1_currLength;
	wire _taskQueues_61_io_connVec_1_push_ready;
	wire _taskQueues_61_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_61_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_60_io_connVec_1_currLength;
	wire _taskQueues_60_io_connVec_1_push_ready;
	wire _taskQueues_60_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_60_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_59_io_connVec_1_currLength;
	wire _taskQueues_59_io_connVec_1_push_ready;
	wire _taskQueues_59_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_59_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_58_io_connVec_1_currLength;
	wire _taskQueues_58_io_connVec_1_push_ready;
	wire _taskQueues_58_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_58_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_57_io_connVec_1_currLength;
	wire _taskQueues_57_io_connVec_1_push_ready;
	wire _taskQueues_57_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_57_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_56_io_connVec_1_currLength;
	wire _taskQueues_56_io_connVec_1_push_ready;
	wire _taskQueues_56_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_56_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_55_io_connVec_1_currLength;
	wire _taskQueues_55_io_connVec_1_push_ready;
	wire _taskQueues_55_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_55_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_54_io_connVec_1_currLength;
	wire _taskQueues_54_io_connVec_1_push_ready;
	wire _taskQueues_54_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_54_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_53_io_connVec_1_currLength;
	wire _taskQueues_53_io_connVec_1_push_ready;
	wire _taskQueues_53_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_53_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_52_io_connVec_1_currLength;
	wire _taskQueues_52_io_connVec_1_push_ready;
	wire _taskQueues_52_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_52_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_51_io_connVec_1_currLength;
	wire _taskQueues_51_io_connVec_1_push_ready;
	wire _taskQueues_51_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_51_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_50_io_connVec_1_currLength;
	wire _taskQueues_50_io_connVec_1_push_ready;
	wire _taskQueues_50_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_50_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_49_io_connVec_1_currLength;
	wire _taskQueues_49_io_connVec_1_push_ready;
	wire _taskQueues_49_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_49_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_48_io_connVec_1_currLength;
	wire _taskQueues_48_io_connVec_1_push_ready;
	wire _taskQueues_48_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_48_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_47_io_connVec_1_currLength;
	wire _taskQueues_47_io_connVec_1_push_ready;
	wire _taskQueues_47_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_47_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_46_io_connVec_1_currLength;
	wire _taskQueues_46_io_connVec_1_push_ready;
	wire _taskQueues_46_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_46_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_45_io_connVec_1_currLength;
	wire _taskQueues_45_io_connVec_1_push_ready;
	wire _taskQueues_45_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_45_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_44_io_connVec_1_currLength;
	wire _taskQueues_44_io_connVec_1_push_ready;
	wire _taskQueues_44_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_44_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_43_io_connVec_1_currLength;
	wire _taskQueues_43_io_connVec_1_push_ready;
	wire _taskQueues_43_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_43_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_42_io_connVec_1_currLength;
	wire _taskQueues_42_io_connVec_1_push_ready;
	wire _taskQueues_42_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_42_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_41_io_connVec_1_currLength;
	wire _taskQueues_41_io_connVec_1_push_ready;
	wire _taskQueues_41_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_41_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_40_io_connVec_1_currLength;
	wire _taskQueues_40_io_connVec_1_push_ready;
	wire _taskQueues_40_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_40_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_39_io_connVec_1_currLength;
	wire _taskQueues_39_io_connVec_1_push_ready;
	wire _taskQueues_39_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_39_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_38_io_connVec_1_currLength;
	wire _taskQueues_38_io_connVec_1_push_ready;
	wire _taskQueues_38_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_38_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_37_io_connVec_1_currLength;
	wire _taskQueues_37_io_connVec_1_push_ready;
	wire _taskQueues_37_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_37_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_36_io_connVec_1_currLength;
	wire _taskQueues_36_io_connVec_1_push_ready;
	wire _taskQueues_36_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_36_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_35_io_connVec_1_currLength;
	wire _taskQueues_35_io_connVec_1_push_ready;
	wire _taskQueues_35_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_35_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_34_io_connVec_1_currLength;
	wire _taskQueues_34_io_connVec_1_push_ready;
	wire _taskQueues_34_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_34_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_33_io_connVec_1_currLength;
	wire _taskQueues_33_io_connVec_1_push_ready;
	wire _taskQueues_33_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_33_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_32_io_connVec_1_currLength;
	wire _taskQueues_32_io_connVec_1_push_ready;
	wire _taskQueues_32_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_32_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_31_io_connVec_1_currLength;
	wire _taskQueues_31_io_connVec_1_push_ready;
	wire _taskQueues_31_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_31_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_30_io_connVec_1_currLength;
	wire _taskQueues_30_io_connVec_1_push_ready;
	wire _taskQueues_30_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_30_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_29_io_connVec_1_currLength;
	wire _taskQueues_29_io_connVec_1_push_ready;
	wire _taskQueues_29_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_29_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_28_io_connVec_1_currLength;
	wire _taskQueues_28_io_connVec_1_push_ready;
	wire _taskQueues_28_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_28_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_27_io_connVec_1_currLength;
	wire _taskQueues_27_io_connVec_1_push_ready;
	wire _taskQueues_27_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_27_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_26_io_connVec_1_currLength;
	wire _taskQueues_26_io_connVec_1_push_ready;
	wire _taskQueues_26_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_26_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_25_io_connVec_1_currLength;
	wire _taskQueues_25_io_connVec_1_push_ready;
	wire _taskQueues_25_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_25_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_24_io_connVec_1_currLength;
	wire _taskQueues_24_io_connVec_1_push_ready;
	wire _taskQueues_24_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_24_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_23_io_connVec_1_currLength;
	wire _taskQueues_23_io_connVec_1_push_ready;
	wire _taskQueues_23_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_23_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_22_io_connVec_1_currLength;
	wire _taskQueues_22_io_connVec_1_push_ready;
	wire _taskQueues_22_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_22_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_21_io_connVec_1_currLength;
	wire _taskQueues_21_io_connVec_1_push_ready;
	wire _taskQueues_21_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_21_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_20_io_connVec_1_currLength;
	wire _taskQueues_20_io_connVec_1_push_ready;
	wire _taskQueues_20_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_20_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_19_io_connVec_1_currLength;
	wire _taskQueues_19_io_connVec_1_push_ready;
	wire _taskQueues_19_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_19_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_18_io_connVec_1_currLength;
	wire _taskQueues_18_io_connVec_1_push_ready;
	wire _taskQueues_18_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_18_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_17_io_connVec_1_currLength;
	wire _taskQueues_17_io_connVec_1_push_ready;
	wire _taskQueues_17_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_17_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_16_io_connVec_1_currLength;
	wire _taskQueues_16_io_connVec_1_push_ready;
	wire _taskQueues_16_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_16_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_15_io_connVec_1_currLength;
	wire _taskQueues_15_io_connVec_1_push_ready;
	wire _taskQueues_15_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_15_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_14_io_connVec_1_currLength;
	wire _taskQueues_14_io_connVec_1_push_ready;
	wire _taskQueues_14_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_14_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_13_io_connVec_1_currLength;
	wire _taskQueues_13_io_connVec_1_push_ready;
	wire _taskQueues_13_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_13_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_12_io_connVec_1_currLength;
	wire _taskQueues_12_io_connVec_1_push_ready;
	wire _taskQueues_12_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_12_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_11_io_connVec_1_currLength;
	wire _taskQueues_11_io_connVec_1_push_ready;
	wire _taskQueues_11_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_11_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_10_io_connVec_1_currLength;
	wire _taskQueues_10_io_connVec_1_push_ready;
	wire _taskQueues_10_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_10_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_9_io_connVec_1_currLength;
	wire _taskQueues_9_io_connVec_1_push_ready;
	wire _taskQueues_9_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_9_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_8_io_connVec_1_currLength;
	wire _taskQueues_8_io_connVec_1_push_ready;
	wire _taskQueues_8_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_8_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_7_io_connVec_1_currLength;
	wire _taskQueues_7_io_connVec_1_push_ready;
	wire _taskQueues_7_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_7_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_6_io_connVec_1_currLength;
	wire _taskQueues_6_io_connVec_1_push_ready;
	wire _taskQueues_6_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_6_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_5_io_connVec_1_currLength;
	wire _taskQueues_5_io_connVec_1_push_ready;
	wire _taskQueues_5_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_5_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_4_io_connVec_1_currLength;
	wire _taskQueues_4_io_connVec_1_push_ready;
	wire _taskQueues_4_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_4_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_3_io_connVec_1_currLength;
	wire _taskQueues_3_io_connVec_1_push_ready;
	wire _taskQueues_3_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_3_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_2_io_connVec_1_currLength;
	wire _taskQueues_2_io_connVec_1_push_ready;
	wire _taskQueues_2_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_2_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_1_io_connVec_1_currLength;
	wire _taskQueues_1_io_connVec_1_push_ready;
	wire _taskQueues_1_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_1_io_connVec_1_pop_bits;
	wire [4:0] _taskQueues_0_io_connVec_1_currLength;
	wire _taskQueues_0_io_connVec_1_push_ready;
	wire _taskQueues_0_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_0_io_connVec_1_pop_bits;
	wire _stealServers_63_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_63_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_63_io_connNetwork_data_availableTask_ready;
	wire _stealServers_63_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_63_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_63_io_connQ_push_valid;
	wire [255:0] _stealServers_63_io_connQ_push_bits;
	wire _stealServers_63_io_connQ_pop_ready;
	wire _stealServers_62_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_62_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_62_io_connNetwork_data_availableTask_ready;
	wire _stealServers_62_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_62_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_62_io_connQ_push_valid;
	wire [255:0] _stealServers_62_io_connQ_push_bits;
	wire _stealServers_62_io_connQ_pop_ready;
	wire _stealServers_61_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_61_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_61_io_connNetwork_data_availableTask_ready;
	wire _stealServers_61_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_61_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_61_io_connQ_push_valid;
	wire [255:0] _stealServers_61_io_connQ_push_bits;
	wire _stealServers_61_io_connQ_pop_ready;
	wire _stealServers_60_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_60_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_60_io_connNetwork_data_availableTask_ready;
	wire _stealServers_60_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_60_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_60_io_connQ_push_valid;
	wire [255:0] _stealServers_60_io_connQ_push_bits;
	wire _stealServers_60_io_connQ_pop_ready;
	wire _stealServers_59_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_59_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_59_io_connNetwork_data_availableTask_ready;
	wire _stealServers_59_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_59_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_59_io_connQ_push_valid;
	wire [255:0] _stealServers_59_io_connQ_push_bits;
	wire _stealServers_59_io_connQ_pop_ready;
	wire _stealServers_58_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_58_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_58_io_connNetwork_data_availableTask_ready;
	wire _stealServers_58_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_58_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_58_io_connQ_push_valid;
	wire [255:0] _stealServers_58_io_connQ_push_bits;
	wire _stealServers_58_io_connQ_pop_ready;
	wire _stealServers_57_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_57_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_57_io_connNetwork_data_availableTask_ready;
	wire _stealServers_57_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_57_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_57_io_connQ_push_valid;
	wire [255:0] _stealServers_57_io_connQ_push_bits;
	wire _stealServers_57_io_connQ_pop_ready;
	wire _stealServers_56_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_56_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_56_io_connNetwork_data_availableTask_ready;
	wire _stealServers_56_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_56_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_56_io_connQ_push_valid;
	wire [255:0] _stealServers_56_io_connQ_push_bits;
	wire _stealServers_56_io_connQ_pop_ready;
	wire _stealServers_55_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_55_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_55_io_connNetwork_data_availableTask_ready;
	wire _stealServers_55_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_55_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_55_io_connQ_push_valid;
	wire [255:0] _stealServers_55_io_connQ_push_bits;
	wire _stealServers_55_io_connQ_pop_ready;
	wire _stealServers_54_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_54_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_54_io_connNetwork_data_availableTask_ready;
	wire _stealServers_54_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_54_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_54_io_connQ_push_valid;
	wire [255:0] _stealServers_54_io_connQ_push_bits;
	wire _stealServers_54_io_connQ_pop_ready;
	wire _stealServers_53_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_53_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_53_io_connNetwork_data_availableTask_ready;
	wire _stealServers_53_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_53_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_53_io_connQ_push_valid;
	wire [255:0] _stealServers_53_io_connQ_push_bits;
	wire _stealServers_53_io_connQ_pop_ready;
	wire _stealServers_52_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_52_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_52_io_connNetwork_data_availableTask_ready;
	wire _stealServers_52_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_52_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_52_io_connQ_push_valid;
	wire [255:0] _stealServers_52_io_connQ_push_bits;
	wire _stealServers_52_io_connQ_pop_ready;
	wire _stealServers_51_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_51_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_51_io_connNetwork_data_availableTask_ready;
	wire _stealServers_51_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_51_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_51_io_connQ_push_valid;
	wire [255:0] _stealServers_51_io_connQ_push_bits;
	wire _stealServers_51_io_connQ_pop_ready;
	wire _stealServers_50_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_50_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_50_io_connNetwork_data_availableTask_ready;
	wire _stealServers_50_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_50_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_50_io_connQ_push_valid;
	wire [255:0] _stealServers_50_io_connQ_push_bits;
	wire _stealServers_50_io_connQ_pop_ready;
	wire _stealServers_49_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_49_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_49_io_connNetwork_data_availableTask_ready;
	wire _stealServers_49_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_49_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_49_io_connQ_push_valid;
	wire [255:0] _stealServers_49_io_connQ_push_bits;
	wire _stealServers_49_io_connQ_pop_ready;
	wire _stealServers_48_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_48_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_48_io_connNetwork_data_availableTask_ready;
	wire _stealServers_48_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_48_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_48_io_connQ_push_valid;
	wire [255:0] _stealServers_48_io_connQ_push_bits;
	wire _stealServers_48_io_connQ_pop_ready;
	wire _stealServers_47_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_47_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_47_io_connNetwork_data_availableTask_ready;
	wire _stealServers_47_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_47_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_47_io_connQ_push_valid;
	wire [255:0] _stealServers_47_io_connQ_push_bits;
	wire _stealServers_47_io_connQ_pop_ready;
	wire _stealServers_46_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_46_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_46_io_connNetwork_data_availableTask_ready;
	wire _stealServers_46_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_46_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_46_io_connQ_push_valid;
	wire [255:0] _stealServers_46_io_connQ_push_bits;
	wire _stealServers_46_io_connQ_pop_ready;
	wire _stealServers_45_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_45_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_45_io_connNetwork_data_availableTask_ready;
	wire _stealServers_45_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_45_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_45_io_connQ_push_valid;
	wire [255:0] _stealServers_45_io_connQ_push_bits;
	wire _stealServers_45_io_connQ_pop_ready;
	wire _stealServers_44_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_44_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_44_io_connNetwork_data_availableTask_ready;
	wire _stealServers_44_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_44_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_44_io_connQ_push_valid;
	wire [255:0] _stealServers_44_io_connQ_push_bits;
	wire _stealServers_44_io_connQ_pop_ready;
	wire _stealServers_43_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_43_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_43_io_connNetwork_data_availableTask_ready;
	wire _stealServers_43_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_43_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_43_io_connQ_push_valid;
	wire [255:0] _stealServers_43_io_connQ_push_bits;
	wire _stealServers_43_io_connQ_pop_ready;
	wire _stealServers_42_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_42_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_42_io_connNetwork_data_availableTask_ready;
	wire _stealServers_42_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_42_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_42_io_connQ_push_valid;
	wire [255:0] _stealServers_42_io_connQ_push_bits;
	wire _stealServers_42_io_connQ_pop_ready;
	wire _stealServers_41_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_41_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_41_io_connNetwork_data_availableTask_ready;
	wire _stealServers_41_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_41_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_41_io_connQ_push_valid;
	wire [255:0] _stealServers_41_io_connQ_push_bits;
	wire _stealServers_41_io_connQ_pop_ready;
	wire _stealServers_40_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_40_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_40_io_connNetwork_data_availableTask_ready;
	wire _stealServers_40_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_40_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_40_io_connQ_push_valid;
	wire [255:0] _stealServers_40_io_connQ_push_bits;
	wire _stealServers_40_io_connQ_pop_ready;
	wire _stealServers_39_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_39_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_39_io_connNetwork_data_availableTask_ready;
	wire _stealServers_39_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_39_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_39_io_connQ_push_valid;
	wire [255:0] _stealServers_39_io_connQ_push_bits;
	wire _stealServers_39_io_connQ_pop_ready;
	wire _stealServers_38_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_38_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_38_io_connNetwork_data_availableTask_ready;
	wire _stealServers_38_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_38_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_38_io_connQ_push_valid;
	wire [255:0] _stealServers_38_io_connQ_push_bits;
	wire _stealServers_38_io_connQ_pop_ready;
	wire _stealServers_37_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_37_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_37_io_connNetwork_data_availableTask_ready;
	wire _stealServers_37_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_37_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_37_io_connQ_push_valid;
	wire [255:0] _stealServers_37_io_connQ_push_bits;
	wire _stealServers_37_io_connQ_pop_ready;
	wire _stealServers_36_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_36_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_36_io_connNetwork_data_availableTask_ready;
	wire _stealServers_36_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_36_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_36_io_connQ_push_valid;
	wire [255:0] _stealServers_36_io_connQ_push_bits;
	wire _stealServers_36_io_connQ_pop_ready;
	wire _stealServers_35_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_35_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_35_io_connNetwork_data_availableTask_ready;
	wire _stealServers_35_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_35_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_35_io_connQ_push_valid;
	wire [255:0] _stealServers_35_io_connQ_push_bits;
	wire _stealServers_35_io_connQ_pop_ready;
	wire _stealServers_34_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_34_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_34_io_connNetwork_data_availableTask_ready;
	wire _stealServers_34_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_34_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_34_io_connQ_push_valid;
	wire [255:0] _stealServers_34_io_connQ_push_bits;
	wire _stealServers_34_io_connQ_pop_ready;
	wire _stealServers_33_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_33_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_33_io_connNetwork_data_availableTask_ready;
	wire _stealServers_33_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_33_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_33_io_connQ_push_valid;
	wire [255:0] _stealServers_33_io_connQ_push_bits;
	wire _stealServers_33_io_connQ_pop_ready;
	wire _stealServers_32_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_32_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_32_io_connNetwork_data_availableTask_ready;
	wire _stealServers_32_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_32_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_32_io_connQ_push_valid;
	wire [255:0] _stealServers_32_io_connQ_push_bits;
	wire _stealServers_32_io_connQ_pop_ready;
	wire _stealServers_31_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_31_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_31_io_connNetwork_data_availableTask_ready;
	wire _stealServers_31_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_31_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_31_io_connQ_push_valid;
	wire [255:0] _stealServers_31_io_connQ_push_bits;
	wire _stealServers_31_io_connQ_pop_ready;
	wire _stealServers_30_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_30_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_30_io_connNetwork_data_availableTask_ready;
	wire _stealServers_30_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_30_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_30_io_connQ_push_valid;
	wire [255:0] _stealServers_30_io_connQ_push_bits;
	wire _stealServers_30_io_connQ_pop_ready;
	wire _stealServers_29_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_29_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_29_io_connNetwork_data_availableTask_ready;
	wire _stealServers_29_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_29_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_29_io_connQ_push_valid;
	wire [255:0] _stealServers_29_io_connQ_push_bits;
	wire _stealServers_29_io_connQ_pop_ready;
	wire _stealServers_28_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_28_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_28_io_connNetwork_data_availableTask_ready;
	wire _stealServers_28_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_28_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_28_io_connQ_push_valid;
	wire [255:0] _stealServers_28_io_connQ_push_bits;
	wire _stealServers_28_io_connQ_pop_ready;
	wire _stealServers_27_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_27_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_27_io_connNetwork_data_availableTask_ready;
	wire _stealServers_27_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_27_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_27_io_connQ_push_valid;
	wire [255:0] _stealServers_27_io_connQ_push_bits;
	wire _stealServers_27_io_connQ_pop_ready;
	wire _stealServers_26_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_26_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_26_io_connNetwork_data_availableTask_ready;
	wire _stealServers_26_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_26_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_26_io_connQ_push_valid;
	wire [255:0] _stealServers_26_io_connQ_push_bits;
	wire _stealServers_26_io_connQ_pop_ready;
	wire _stealServers_25_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_25_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_25_io_connNetwork_data_availableTask_ready;
	wire _stealServers_25_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_25_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_25_io_connQ_push_valid;
	wire [255:0] _stealServers_25_io_connQ_push_bits;
	wire _stealServers_25_io_connQ_pop_ready;
	wire _stealServers_24_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_24_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_24_io_connNetwork_data_availableTask_ready;
	wire _stealServers_24_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_24_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_24_io_connQ_push_valid;
	wire [255:0] _stealServers_24_io_connQ_push_bits;
	wire _stealServers_24_io_connQ_pop_ready;
	wire _stealServers_23_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_23_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_23_io_connNetwork_data_availableTask_ready;
	wire _stealServers_23_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_23_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_23_io_connQ_push_valid;
	wire [255:0] _stealServers_23_io_connQ_push_bits;
	wire _stealServers_23_io_connQ_pop_ready;
	wire _stealServers_22_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_22_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_22_io_connNetwork_data_availableTask_ready;
	wire _stealServers_22_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_22_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_22_io_connQ_push_valid;
	wire [255:0] _stealServers_22_io_connQ_push_bits;
	wire _stealServers_22_io_connQ_pop_ready;
	wire _stealServers_21_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_21_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_21_io_connNetwork_data_availableTask_ready;
	wire _stealServers_21_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_21_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_21_io_connQ_push_valid;
	wire [255:0] _stealServers_21_io_connQ_push_bits;
	wire _stealServers_21_io_connQ_pop_ready;
	wire _stealServers_20_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_20_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_20_io_connNetwork_data_availableTask_ready;
	wire _stealServers_20_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_20_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_20_io_connQ_push_valid;
	wire [255:0] _stealServers_20_io_connQ_push_bits;
	wire _stealServers_20_io_connQ_pop_ready;
	wire _stealServers_19_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_19_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_19_io_connNetwork_data_availableTask_ready;
	wire _stealServers_19_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_19_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_19_io_connQ_push_valid;
	wire [255:0] _stealServers_19_io_connQ_push_bits;
	wire _stealServers_19_io_connQ_pop_ready;
	wire _stealServers_18_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_18_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_18_io_connNetwork_data_availableTask_ready;
	wire _stealServers_18_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_18_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_18_io_connQ_push_valid;
	wire [255:0] _stealServers_18_io_connQ_push_bits;
	wire _stealServers_18_io_connQ_pop_ready;
	wire _stealServers_17_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_17_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_17_io_connNetwork_data_availableTask_ready;
	wire _stealServers_17_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_17_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_17_io_connQ_push_valid;
	wire [255:0] _stealServers_17_io_connQ_push_bits;
	wire _stealServers_17_io_connQ_pop_ready;
	wire _stealServers_16_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_16_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_16_io_connNetwork_data_availableTask_ready;
	wire _stealServers_16_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_16_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_16_io_connQ_push_valid;
	wire [255:0] _stealServers_16_io_connQ_push_bits;
	wire _stealServers_16_io_connQ_pop_ready;
	wire _stealServers_15_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_15_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_15_io_connNetwork_data_availableTask_ready;
	wire _stealServers_15_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_15_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_15_io_connQ_push_valid;
	wire [255:0] _stealServers_15_io_connQ_push_bits;
	wire _stealServers_15_io_connQ_pop_ready;
	wire _stealServers_14_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_14_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_14_io_connNetwork_data_availableTask_ready;
	wire _stealServers_14_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_14_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_14_io_connQ_push_valid;
	wire [255:0] _stealServers_14_io_connQ_push_bits;
	wire _stealServers_14_io_connQ_pop_ready;
	wire _stealServers_13_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_13_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_13_io_connNetwork_data_availableTask_ready;
	wire _stealServers_13_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_13_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_13_io_connQ_push_valid;
	wire [255:0] _stealServers_13_io_connQ_push_bits;
	wire _stealServers_13_io_connQ_pop_ready;
	wire _stealServers_12_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_12_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_12_io_connNetwork_data_availableTask_ready;
	wire _stealServers_12_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_12_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_12_io_connQ_push_valid;
	wire [255:0] _stealServers_12_io_connQ_push_bits;
	wire _stealServers_12_io_connQ_pop_ready;
	wire _stealServers_11_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_11_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_11_io_connNetwork_data_availableTask_ready;
	wire _stealServers_11_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_11_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_11_io_connQ_push_valid;
	wire [255:0] _stealServers_11_io_connQ_push_bits;
	wire _stealServers_11_io_connQ_pop_ready;
	wire _stealServers_10_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_10_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_10_io_connNetwork_data_availableTask_ready;
	wire _stealServers_10_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_10_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_10_io_connQ_push_valid;
	wire [255:0] _stealServers_10_io_connQ_push_bits;
	wire _stealServers_10_io_connQ_pop_ready;
	wire _stealServers_9_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_9_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_9_io_connNetwork_data_availableTask_ready;
	wire _stealServers_9_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_9_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_9_io_connQ_push_valid;
	wire [255:0] _stealServers_9_io_connQ_push_bits;
	wire _stealServers_9_io_connQ_pop_ready;
	wire _stealServers_8_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_8_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_8_io_connNetwork_data_availableTask_ready;
	wire _stealServers_8_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_8_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_8_io_connQ_push_valid;
	wire [255:0] _stealServers_8_io_connQ_push_bits;
	wire _stealServers_8_io_connQ_pop_ready;
	wire _stealServers_7_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_7_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_7_io_connNetwork_data_availableTask_ready;
	wire _stealServers_7_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_7_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_7_io_connQ_push_valid;
	wire [255:0] _stealServers_7_io_connQ_push_bits;
	wire _stealServers_7_io_connQ_pop_ready;
	wire _stealServers_6_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_6_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_6_io_connNetwork_data_availableTask_ready;
	wire _stealServers_6_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_6_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_6_io_connQ_push_valid;
	wire [255:0] _stealServers_6_io_connQ_push_bits;
	wire _stealServers_6_io_connQ_pop_ready;
	wire _stealServers_5_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_5_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_5_io_connNetwork_data_availableTask_ready;
	wire _stealServers_5_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_5_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_5_io_connQ_push_valid;
	wire [255:0] _stealServers_5_io_connQ_push_bits;
	wire _stealServers_5_io_connQ_pop_ready;
	wire _stealServers_4_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_4_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_4_io_connNetwork_data_availableTask_ready;
	wire _stealServers_4_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_4_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_4_io_connQ_push_valid;
	wire [255:0] _stealServers_4_io_connQ_push_bits;
	wire _stealServers_4_io_connQ_pop_ready;
	wire _stealServers_3_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_3_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_3_io_connNetwork_data_availableTask_ready;
	wire _stealServers_3_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_3_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_3_io_connQ_push_valid;
	wire [255:0] _stealServers_3_io_connQ_push_bits;
	wire _stealServers_3_io_connQ_pop_ready;
	wire _stealServers_2_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_2_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_2_io_connNetwork_data_availableTask_ready;
	wire _stealServers_2_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_2_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_2_io_connQ_push_valid;
	wire [255:0] _stealServers_2_io_connQ_push_bits;
	wire _stealServers_2_io_connQ_pop_ready;
	wire _stealServers_1_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_1_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_1_io_connNetwork_data_availableTask_ready;
	wire _stealServers_1_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_1_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_1_io_connQ_push_valid;
	wire [255:0] _stealServers_1_io_connQ_push_bits;
	wire _stealServers_1_io_connQ_pop_ready;
	wire _stealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_0_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_0_io_connNetwork_data_availableTask_ready;
	wire _stealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_0_io_connQ_push_valid;
	wire [255:0] _stealServers_0_io_connQ_push_bits;
	wire _stealServers_0_io_connQ_pop_ready;
	wire _stealNet_io_connSS_18_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_18_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_18_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_18_data_availableTask_bits;
	wire _stealNet_io_connSS_18_data_qOutTask_ready;
	wire _stealNet_io_connSS_19_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_19_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_19_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_19_data_availableTask_bits;
	wire _stealNet_io_connSS_19_data_qOutTask_ready;
	wire _stealNet_io_connSS_20_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_20_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_20_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_20_data_availableTask_bits;
	wire _stealNet_io_connSS_20_data_qOutTask_ready;
	wire _stealNet_io_connSS_21_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_21_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_21_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_21_data_availableTask_bits;
	wire _stealNet_io_connSS_21_data_qOutTask_ready;
	wire _stealNet_io_connSS_22_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_22_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_22_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_22_data_availableTask_bits;
	wire _stealNet_io_connSS_22_data_qOutTask_ready;
	wire _stealNet_io_connSS_23_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_23_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_23_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_23_data_availableTask_bits;
	wire _stealNet_io_connSS_23_data_qOutTask_ready;
	wire _stealNet_io_connSS_24_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_24_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_24_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_24_data_availableTask_bits;
	wire _stealNet_io_connSS_24_data_qOutTask_ready;
	wire _stealNet_io_connSS_25_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_25_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_25_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_25_data_availableTask_bits;
	wire _stealNet_io_connSS_25_data_qOutTask_ready;
	wire _stealNet_io_connSS_26_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_26_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_26_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_26_data_availableTask_bits;
	wire _stealNet_io_connSS_26_data_qOutTask_ready;
	wire _stealNet_io_connSS_27_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_27_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_27_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_27_data_availableTask_bits;
	wire _stealNet_io_connSS_27_data_qOutTask_ready;
	wire _stealNet_io_connSS_28_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_28_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_28_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_28_data_availableTask_bits;
	wire _stealNet_io_connSS_28_data_qOutTask_ready;
	wire _stealNet_io_connSS_29_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_29_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_29_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_29_data_availableTask_bits;
	wire _stealNet_io_connSS_29_data_qOutTask_ready;
	wire _stealNet_io_connSS_30_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_30_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_30_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_30_data_availableTask_bits;
	wire _stealNet_io_connSS_30_data_qOutTask_ready;
	wire _stealNet_io_connSS_31_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_31_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_31_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_31_data_availableTask_bits;
	wire _stealNet_io_connSS_31_data_qOutTask_ready;
	wire _stealNet_io_connSS_32_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_32_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_32_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_32_data_availableTask_bits;
	wire _stealNet_io_connSS_32_data_qOutTask_ready;
	wire _stealNet_io_connSS_33_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_33_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_33_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_33_data_availableTask_bits;
	wire _stealNet_io_connSS_33_data_qOutTask_ready;
	wire _stealNet_io_connSS_34_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_34_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_34_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_34_data_availableTask_bits;
	wire _stealNet_io_connSS_34_data_qOutTask_ready;
	wire _stealNet_io_connSS_35_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_35_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_35_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_35_data_availableTask_bits;
	wire _stealNet_io_connSS_35_data_qOutTask_ready;
	wire _stealNet_io_connSS_36_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_36_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_36_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_36_data_availableTask_bits;
	wire _stealNet_io_connSS_36_data_qOutTask_ready;
	wire _stealNet_io_connSS_37_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_37_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_37_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_37_data_availableTask_bits;
	wire _stealNet_io_connSS_37_data_qOutTask_ready;
	wire _stealNet_io_connSS_38_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_38_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_38_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_38_data_availableTask_bits;
	wire _stealNet_io_connSS_38_data_qOutTask_ready;
	wire _stealNet_io_connSS_39_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_39_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_39_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_39_data_availableTask_bits;
	wire _stealNet_io_connSS_39_data_qOutTask_ready;
	wire _stealNet_io_connSS_40_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_40_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_40_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_40_data_availableTask_bits;
	wire _stealNet_io_connSS_40_data_qOutTask_ready;
	wire _stealNet_io_connSS_41_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_41_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_41_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_41_data_availableTask_bits;
	wire _stealNet_io_connSS_41_data_qOutTask_ready;
	wire _stealNet_io_connSS_42_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_42_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_42_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_42_data_availableTask_bits;
	wire _stealNet_io_connSS_42_data_qOutTask_ready;
	wire _stealNet_io_connSS_43_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_43_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_43_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_43_data_availableTask_bits;
	wire _stealNet_io_connSS_43_data_qOutTask_ready;
	wire _stealNet_io_connSS_44_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_44_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_44_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_44_data_availableTask_bits;
	wire _stealNet_io_connSS_44_data_qOutTask_ready;
	wire _stealNet_io_connSS_45_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_45_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_45_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_45_data_availableTask_bits;
	wire _stealNet_io_connSS_45_data_qOutTask_ready;
	wire _stealNet_io_connSS_46_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_46_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_46_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_46_data_availableTask_bits;
	wire _stealNet_io_connSS_46_data_qOutTask_ready;
	wire _stealNet_io_connSS_47_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_47_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_47_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_47_data_availableTask_bits;
	wire _stealNet_io_connSS_47_data_qOutTask_ready;
	wire _stealNet_io_connSS_48_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_48_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_48_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_48_data_availableTask_bits;
	wire _stealNet_io_connSS_48_data_qOutTask_ready;
	wire _stealNet_io_connSS_49_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_49_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_49_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_49_data_availableTask_bits;
	wire _stealNet_io_connSS_49_data_qOutTask_ready;
	wire _stealNet_io_connSS_50_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_50_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_50_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_50_data_availableTask_bits;
	wire _stealNet_io_connSS_50_data_qOutTask_ready;
	wire _stealNet_io_connSS_51_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_51_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_51_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_51_data_availableTask_bits;
	wire _stealNet_io_connSS_51_data_qOutTask_ready;
	wire _stealNet_io_connSS_52_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_52_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_52_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_52_data_availableTask_bits;
	wire _stealNet_io_connSS_52_data_qOutTask_ready;
	wire _stealNet_io_connSS_53_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_53_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_53_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_53_data_availableTask_bits;
	wire _stealNet_io_connSS_53_data_qOutTask_ready;
	wire _stealNet_io_connSS_54_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_54_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_54_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_54_data_availableTask_bits;
	wire _stealNet_io_connSS_54_data_qOutTask_ready;
	wire _stealNet_io_connSS_55_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_55_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_55_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_55_data_availableTask_bits;
	wire _stealNet_io_connSS_55_data_qOutTask_ready;
	wire _stealNet_io_connSS_56_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_56_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_56_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_56_data_availableTask_bits;
	wire _stealNet_io_connSS_56_data_qOutTask_ready;
	wire _stealNet_io_connSS_57_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_57_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_57_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_57_data_availableTask_bits;
	wire _stealNet_io_connSS_57_data_qOutTask_ready;
	wire _stealNet_io_connSS_58_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_58_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_58_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_58_data_availableTask_bits;
	wire _stealNet_io_connSS_58_data_qOutTask_ready;
	wire _stealNet_io_connSS_59_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_59_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_59_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_59_data_availableTask_bits;
	wire _stealNet_io_connSS_59_data_qOutTask_ready;
	wire _stealNet_io_connSS_60_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_60_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_60_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_60_data_availableTask_bits;
	wire _stealNet_io_connSS_60_data_qOutTask_ready;
	wire _stealNet_io_connSS_61_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_61_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_61_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_61_data_availableTask_bits;
	wire _stealNet_io_connSS_61_data_qOutTask_ready;
	wire _stealNet_io_connSS_62_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_62_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_62_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_62_data_availableTask_bits;
	wire _stealNet_io_connSS_62_data_qOutTask_ready;
	wire _stealNet_io_connSS_63_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_63_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_63_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_63_data_availableTask_bits;
	wire _stealNet_io_connSS_63_data_qOutTask_ready;
	wire _stealNet_io_connSS_64_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_64_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_64_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_64_data_availableTask_bits;
	wire _stealNet_io_connSS_64_data_qOutTask_ready;
	wire _stealNet_io_connSS_65_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_65_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_65_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_65_data_availableTask_bits;
	wire _stealNet_io_connSS_65_data_qOutTask_ready;
	wire _stealNet_io_connSS_66_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_66_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_66_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_66_data_availableTask_bits;
	wire _stealNet_io_connSS_66_data_qOutTask_ready;
	wire _stealNet_io_connSS_67_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_67_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_67_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_67_data_availableTask_bits;
	wire _stealNet_io_connSS_67_data_qOutTask_ready;
	wire _stealNet_io_connSS_68_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_68_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_68_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_68_data_availableTask_bits;
	wire _stealNet_io_connSS_68_data_qOutTask_ready;
	wire _stealNet_io_connSS_69_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_69_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_69_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_69_data_availableTask_bits;
	wire _stealNet_io_connSS_69_data_qOutTask_ready;
	wire _stealNet_io_connSS_70_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_70_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_70_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_70_data_availableTask_bits;
	wire _stealNet_io_connSS_70_data_qOutTask_ready;
	wire _stealNet_io_connSS_71_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_71_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_71_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_71_data_availableTask_bits;
	wire _stealNet_io_connSS_71_data_qOutTask_ready;
	wire _stealNet_io_connSS_72_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_72_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_72_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_72_data_availableTask_bits;
	wire _stealNet_io_connSS_72_data_qOutTask_ready;
	wire _stealNet_io_connSS_73_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_73_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_73_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_73_data_availableTask_bits;
	wire _stealNet_io_connSS_73_data_qOutTask_ready;
	wire _stealNet_io_connSS_74_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_74_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_74_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_74_data_availableTask_bits;
	wire _stealNet_io_connSS_74_data_qOutTask_ready;
	wire _stealNet_io_connSS_75_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_75_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_75_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_75_data_availableTask_bits;
	wire _stealNet_io_connSS_75_data_qOutTask_ready;
	wire _stealNet_io_connSS_76_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_76_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_76_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_76_data_availableTask_bits;
	wire _stealNet_io_connSS_76_data_qOutTask_ready;
	wire _stealNet_io_connSS_77_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_77_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_77_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_77_data_availableTask_bits;
	wire _stealNet_io_connSS_77_data_qOutTask_ready;
	wire _stealNet_io_connSS_78_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_78_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_78_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_78_data_availableTask_bits;
	wire _stealNet_io_connSS_78_data_qOutTask_ready;
	wire _stealNet_io_connSS_79_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_79_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_79_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_79_data_availableTask_bits;
	wire _stealNet_io_connSS_79_data_qOutTask_ready;
	wire _stealNet_io_connSS_80_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_80_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_80_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_80_data_availableTask_bits;
	wire _stealNet_io_connSS_80_data_qOutTask_ready;
	wire _stealNet_io_connSS_81_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_81_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_81_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_81_data_availableTask_bits;
	wire _stealNet_io_connSS_81_data_qOutTask_ready;
	SchedulerNetwork_1 stealNet(
		.clock(clock),
		.reset(reset),
		.io_connSS_0_ctrl_serveStealReq_valid(io_connVAS_0_ctrl_serveStealReq_valid),
		.io_connSS_0_ctrl_serveStealReq_ready(io_connVAS_0_ctrl_serveStealReq_ready),
		.io_connSS_0_data_availableTask_ready(io_connVSS_0_data_availableTask_ready),
		.io_connSS_0_data_availableTask_valid(io_connVSS_0_data_availableTask_valid),
		.io_connSS_0_data_availableTask_bits(io_connVSS_0_data_availableTask_bits),
		.io_connSS_0_data_qOutTask_ready(io_connVSS_0_data_qOutTask_ready),
		.io_connSS_0_data_qOutTask_valid(io_connVSS_0_data_qOutTask_valid),
		.io_connSS_0_data_qOutTask_bits(io_connVSS_0_data_qOutTask_bits),
		.io_connSS_1_ctrl_serveStealReq_valid(io_connVAS_1_ctrl_serveStealReq_valid),
		.io_connSS_1_ctrl_serveStealReq_ready(io_connVAS_1_ctrl_serveStealReq_ready),
		.io_connSS_1_data_availableTask_ready(io_connVSS_1_data_availableTask_ready),
		.io_connSS_1_data_availableTask_valid(io_connVSS_1_data_availableTask_valid),
		.io_connSS_1_data_availableTask_bits(io_connVSS_1_data_availableTask_bits),
		.io_connSS_1_data_qOutTask_ready(io_connVSS_1_data_qOutTask_ready),
		.io_connSS_1_data_qOutTask_valid(io_connVSS_1_data_qOutTask_valid),
		.io_connSS_1_data_qOutTask_bits(io_connVSS_1_data_qOutTask_bits),
		.io_connSS_2_ctrl_serveStealReq_valid(io_connVAS_2_ctrl_serveStealReq_valid),
		.io_connSS_2_ctrl_serveStealReq_ready(io_connVAS_2_ctrl_serveStealReq_ready),
		.io_connSS_2_data_qOutTask_ready(io_connVAS_0_data_qOutTask_ready),
		.io_connSS_2_data_qOutTask_valid(io_connVAS_0_data_qOutTask_valid),
		.io_connSS_2_data_qOutTask_bits(io_connVAS_0_data_qOutTask_bits),
		.io_connSS_3_ctrl_serveStealReq_valid(io_connVAS_3_ctrl_serveStealReq_valid),
		.io_connSS_3_ctrl_serveStealReq_ready(io_connVAS_3_ctrl_serveStealReq_ready),
		.io_connSS_3_data_qOutTask_ready(io_connVAS_1_data_qOutTask_ready),
		.io_connSS_3_data_qOutTask_valid(io_connVAS_1_data_qOutTask_valid),
		.io_connSS_3_data_qOutTask_bits(io_connVAS_1_data_qOutTask_bits),
		.io_connSS_4_ctrl_serveStealReq_valid(io_connVAS_4_ctrl_serveStealReq_valid),
		.io_connSS_4_ctrl_serveStealReq_ready(io_connVAS_4_ctrl_serveStealReq_ready),
		.io_connSS_4_data_qOutTask_ready(io_connVAS_2_data_qOutTask_ready),
		.io_connSS_4_data_qOutTask_valid(io_connVAS_2_data_qOutTask_valid),
		.io_connSS_4_data_qOutTask_bits(io_connVAS_2_data_qOutTask_bits),
		.io_connSS_5_ctrl_serveStealReq_valid(io_connVAS_5_ctrl_serveStealReq_valid),
		.io_connSS_5_ctrl_serveStealReq_ready(io_connVAS_5_ctrl_serveStealReq_ready),
		.io_connSS_5_data_qOutTask_ready(io_connVAS_3_data_qOutTask_ready),
		.io_connSS_5_data_qOutTask_valid(io_connVAS_3_data_qOutTask_valid),
		.io_connSS_5_data_qOutTask_bits(io_connVAS_3_data_qOutTask_bits),
		.io_connSS_6_ctrl_serveStealReq_valid(io_connVAS_6_ctrl_serveStealReq_valid),
		.io_connSS_6_ctrl_serveStealReq_ready(io_connVAS_6_ctrl_serveStealReq_ready),
		.io_connSS_6_data_qOutTask_ready(io_connVAS_4_data_qOutTask_ready),
		.io_connSS_6_data_qOutTask_valid(io_connVAS_4_data_qOutTask_valid),
		.io_connSS_6_data_qOutTask_bits(io_connVAS_4_data_qOutTask_bits),
		.io_connSS_7_ctrl_serveStealReq_valid(io_connVAS_7_ctrl_serveStealReq_valid),
		.io_connSS_7_ctrl_serveStealReq_ready(io_connVAS_7_ctrl_serveStealReq_ready),
		.io_connSS_7_data_qOutTask_ready(io_connVAS_5_data_qOutTask_ready),
		.io_connSS_7_data_qOutTask_valid(io_connVAS_5_data_qOutTask_valid),
		.io_connSS_7_data_qOutTask_bits(io_connVAS_5_data_qOutTask_bits),
		.io_connSS_8_ctrl_serveStealReq_valid(io_connVAS_8_ctrl_serveStealReq_valid),
		.io_connSS_8_ctrl_serveStealReq_ready(io_connVAS_8_ctrl_serveStealReq_ready),
		.io_connSS_8_data_qOutTask_ready(io_connVAS_6_data_qOutTask_ready),
		.io_connSS_8_data_qOutTask_valid(io_connVAS_6_data_qOutTask_valid),
		.io_connSS_8_data_qOutTask_bits(io_connVAS_6_data_qOutTask_bits),
		.io_connSS_9_ctrl_serveStealReq_valid(io_connVAS_9_ctrl_serveStealReq_valid),
		.io_connSS_9_ctrl_serveStealReq_ready(io_connVAS_9_ctrl_serveStealReq_ready),
		.io_connSS_9_data_qOutTask_ready(io_connVAS_7_data_qOutTask_ready),
		.io_connSS_9_data_qOutTask_valid(io_connVAS_7_data_qOutTask_valid),
		.io_connSS_9_data_qOutTask_bits(io_connVAS_7_data_qOutTask_bits),
		.io_connSS_10_ctrl_serveStealReq_valid(io_connVAS_10_ctrl_serveStealReq_valid),
		.io_connSS_10_ctrl_serveStealReq_ready(io_connVAS_10_ctrl_serveStealReq_ready),
		.io_connSS_10_data_qOutTask_ready(io_connVAS_8_data_qOutTask_ready),
		.io_connSS_10_data_qOutTask_valid(io_connVAS_8_data_qOutTask_valid),
		.io_connSS_10_data_qOutTask_bits(io_connVAS_8_data_qOutTask_bits),
		.io_connSS_11_ctrl_serveStealReq_valid(io_connVAS_11_ctrl_serveStealReq_valid),
		.io_connSS_11_ctrl_serveStealReq_ready(io_connVAS_11_ctrl_serveStealReq_ready),
		.io_connSS_11_data_qOutTask_ready(io_connVAS_9_data_qOutTask_ready),
		.io_connSS_11_data_qOutTask_valid(io_connVAS_9_data_qOutTask_valid),
		.io_connSS_11_data_qOutTask_bits(io_connVAS_9_data_qOutTask_bits),
		.io_connSS_12_ctrl_serveStealReq_valid(io_connVAS_12_ctrl_serveStealReq_valid),
		.io_connSS_12_ctrl_serveStealReq_ready(io_connVAS_12_ctrl_serveStealReq_ready),
		.io_connSS_12_data_qOutTask_ready(io_connVAS_10_data_qOutTask_ready),
		.io_connSS_12_data_qOutTask_valid(io_connVAS_10_data_qOutTask_valid),
		.io_connSS_12_data_qOutTask_bits(io_connVAS_10_data_qOutTask_bits),
		.io_connSS_13_ctrl_serveStealReq_valid(io_connVAS_13_ctrl_serveStealReq_valid),
		.io_connSS_13_ctrl_serveStealReq_ready(io_connVAS_13_ctrl_serveStealReq_ready),
		.io_connSS_13_data_qOutTask_ready(io_connVAS_11_data_qOutTask_ready),
		.io_connSS_13_data_qOutTask_valid(io_connVAS_11_data_qOutTask_valid),
		.io_connSS_13_data_qOutTask_bits(io_connVAS_11_data_qOutTask_bits),
		.io_connSS_14_ctrl_serveStealReq_valid(io_connVAS_14_ctrl_serveStealReq_valid),
		.io_connSS_14_ctrl_serveStealReq_ready(io_connVAS_14_ctrl_serveStealReq_ready),
		.io_connSS_14_data_qOutTask_ready(io_connVAS_12_data_qOutTask_ready),
		.io_connSS_14_data_qOutTask_valid(io_connVAS_12_data_qOutTask_valid),
		.io_connSS_14_data_qOutTask_bits(io_connVAS_12_data_qOutTask_bits),
		.io_connSS_15_ctrl_serveStealReq_valid(io_connVAS_15_ctrl_serveStealReq_valid),
		.io_connSS_15_ctrl_serveStealReq_ready(io_connVAS_15_ctrl_serveStealReq_ready),
		.io_connSS_15_data_qOutTask_ready(io_connVAS_13_data_qOutTask_ready),
		.io_connSS_15_data_qOutTask_valid(io_connVAS_13_data_qOutTask_valid),
		.io_connSS_15_data_qOutTask_bits(io_connVAS_13_data_qOutTask_bits),
		.io_connSS_16_ctrl_serveStealReq_valid(io_connVSS_0_ctrl_serveStealReq_valid),
		.io_connSS_16_ctrl_serveStealReq_ready(io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connSS_16_data_qOutTask_ready(io_connVAS_14_data_qOutTask_ready),
		.io_connSS_16_data_qOutTask_valid(io_connVAS_14_data_qOutTask_valid),
		.io_connSS_16_data_qOutTask_bits(io_connVAS_14_data_qOutTask_bits),
		.io_connSS_17_ctrl_serveStealReq_valid(io_connVSS_1_ctrl_serveStealReq_valid),
		.io_connSS_17_ctrl_serveStealReq_ready(io_connVSS_1_ctrl_serveStealReq_ready),
		.io_connSS_17_data_qOutTask_ready(io_connVAS_15_data_qOutTask_ready),
		.io_connSS_17_data_qOutTask_valid(io_connVAS_15_data_qOutTask_valid),
		.io_connSS_17_data_qOutTask_bits(io_connVAS_15_data_qOutTask_bits),
		.io_connSS_18_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_18_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_18_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_18_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connSS_18_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connSS_18_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connSS_18_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connSS_18_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connSS_18_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connSS_18_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connSS_19_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_19_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_19_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_19_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connSS_19_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connSS_19_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connSS_19_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connSS_19_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connSS_19_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connSS_19_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connSS_20_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_20_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_20_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_20_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connSS_20_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connSS_20_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connSS_20_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connSS_20_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connSS_20_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connSS_20_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connSS_21_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_21_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_21_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_21_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connSS_21_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connSS_21_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connSS_21_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connSS_21_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connSS_21_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connSS_21_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connSS_22_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_22_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_22_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_22_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connSS_22_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connSS_22_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connSS_22_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connSS_22_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connSS_22_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connSS_22_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connSS_23_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_23_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_23_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_23_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connSS_23_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connSS_23_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connSS_23_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connSS_23_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connSS_23_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connSS_23_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connSS_24_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_24_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_24_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_24_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connSS_24_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connSS_24_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connSS_24_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connSS_24_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connSS_24_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connSS_24_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connSS_25_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_25_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_25_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_25_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connSS_25_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connSS_25_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connSS_25_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connSS_25_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connSS_25_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connSS_25_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connSS_26_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_26_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_26_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_26_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connSS_26_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connSS_26_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connSS_26_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connSS_26_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connSS_26_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connSS_26_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connSS_27_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_27_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_27_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_27_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connSS_27_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connSS_27_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connSS_27_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connSS_27_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connSS_27_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connSS_27_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connSS_28_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_28_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_28_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_28_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connSS_28_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connSS_28_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connSS_28_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connSS_28_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connSS_28_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connSS_28_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connSS_29_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_29_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_29_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_29_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connSS_29_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connSS_29_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connSS_29_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connSS_29_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connSS_29_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connSS_29_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connSS_30_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_30_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_30_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_30_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connSS_30_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connSS_30_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connSS_30_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connSS_30_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connSS_30_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connSS_30_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connSS_31_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_31_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_31_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_31_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connSS_31_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connSS_31_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connSS_31_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connSS_31_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connSS_31_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connSS_31_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connSS_32_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_32_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_32_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_32_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connSS_32_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connSS_32_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connSS_32_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connSS_32_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connSS_32_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connSS_32_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connSS_33_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_33_ctrl_serveStealReq_ready(_stealNet_io_connSS_33_ctrl_serveStealReq_ready),
		.io_connSS_33_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_33_ctrl_stealReq_ready(_stealNet_io_connSS_33_ctrl_stealReq_ready),
		.io_connSS_33_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connSS_33_data_availableTask_valid(_stealNet_io_connSS_33_data_availableTask_valid),
		.io_connSS_33_data_availableTask_bits(_stealNet_io_connSS_33_data_availableTask_bits),
		.io_connSS_33_data_qOutTask_ready(_stealNet_io_connSS_33_data_qOutTask_ready),
		.io_connSS_33_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connSS_33_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connSS_34_ctrl_serveStealReq_valid(_stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_34_ctrl_serveStealReq_ready(_stealNet_io_connSS_34_ctrl_serveStealReq_ready),
		.io_connSS_34_ctrl_stealReq_valid(_stealServers_16_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_34_ctrl_stealReq_ready(_stealNet_io_connSS_34_ctrl_stealReq_ready),
		.io_connSS_34_data_availableTask_ready(_stealServers_16_io_connNetwork_data_availableTask_ready),
		.io_connSS_34_data_availableTask_valid(_stealNet_io_connSS_34_data_availableTask_valid),
		.io_connSS_34_data_availableTask_bits(_stealNet_io_connSS_34_data_availableTask_bits),
		.io_connSS_34_data_qOutTask_ready(_stealNet_io_connSS_34_data_qOutTask_ready),
		.io_connSS_34_data_qOutTask_valid(_stealServers_16_io_connNetwork_data_qOutTask_valid),
		.io_connSS_34_data_qOutTask_bits(_stealServers_16_io_connNetwork_data_qOutTask_bits),
		.io_connSS_35_ctrl_serveStealReq_valid(_stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_35_ctrl_serveStealReq_ready(_stealNet_io_connSS_35_ctrl_serveStealReq_ready),
		.io_connSS_35_ctrl_stealReq_valid(_stealServers_17_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_35_ctrl_stealReq_ready(_stealNet_io_connSS_35_ctrl_stealReq_ready),
		.io_connSS_35_data_availableTask_ready(_stealServers_17_io_connNetwork_data_availableTask_ready),
		.io_connSS_35_data_availableTask_valid(_stealNet_io_connSS_35_data_availableTask_valid),
		.io_connSS_35_data_availableTask_bits(_stealNet_io_connSS_35_data_availableTask_bits),
		.io_connSS_35_data_qOutTask_ready(_stealNet_io_connSS_35_data_qOutTask_ready),
		.io_connSS_35_data_qOutTask_valid(_stealServers_17_io_connNetwork_data_qOutTask_valid),
		.io_connSS_35_data_qOutTask_bits(_stealServers_17_io_connNetwork_data_qOutTask_bits),
		.io_connSS_36_ctrl_serveStealReq_valid(_stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_36_ctrl_serveStealReq_ready(_stealNet_io_connSS_36_ctrl_serveStealReq_ready),
		.io_connSS_36_ctrl_stealReq_valid(_stealServers_18_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_36_ctrl_stealReq_ready(_stealNet_io_connSS_36_ctrl_stealReq_ready),
		.io_connSS_36_data_availableTask_ready(_stealServers_18_io_connNetwork_data_availableTask_ready),
		.io_connSS_36_data_availableTask_valid(_stealNet_io_connSS_36_data_availableTask_valid),
		.io_connSS_36_data_availableTask_bits(_stealNet_io_connSS_36_data_availableTask_bits),
		.io_connSS_36_data_qOutTask_ready(_stealNet_io_connSS_36_data_qOutTask_ready),
		.io_connSS_36_data_qOutTask_valid(_stealServers_18_io_connNetwork_data_qOutTask_valid),
		.io_connSS_36_data_qOutTask_bits(_stealServers_18_io_connNetwork_data_qOutTask_bits),
		.io_connSS_37_ctrl_serveStealReq_valid(_stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_37_ctrl_serveStealReq_ready(_stealNet_io_connSS_37_ctrl_serveStealReq_ready),
		.io_connSS_37_ctrl_stealReq_valid(_stealServers_19_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_37_ctrl_stealReq_ready(_stealNet_io_connSS_37_ctrl_stealReq_ready),
		.io_connSS_37_data_availableTask_ready(_stealServers_19_io_connNetwork_data_availableTask_ready),
		.io_connSS_37_data_availableTask_valid(_stealNet_io_connSS_37_data_availableTask_valid),
		.io_connSS_37_data_availableTask_bits(_stealNet_io_connSS_37_data_availableTask_bits),
		.io_connSS_37_data_qOutTask_ready(_stealNet_io_connSS_37_data_qOutTask_ready),
		.io_connSS_37_data_qOutTask_valid(_stealServers_19_io_connNetwork_data_qOutTask_valid),
		.io_connSS_37_data_qOutTask_bits(_stealServers_19_io_connNetwork_data_qOutTask_bits),
		.io_connSS_38_ctrl_serveStealReq_valid(_stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_38_ctrl_serveStealReq_ready(_stealNet_io_connSS_38_ctrl_serveStealReq_ready),
		.io_connSS_38_ctrl_stealReq_valid(_stealServers_20_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_38_ctrl_stealReq_ready(_stealNet_io_connSS_38_ctrl_stealReq_ready),
		.io_connSS_38_data_availableTask_ready(_stealServers_20_io_connNetwork_data_availableTask_ready),
		.io_connSS_38_data_availableTask_valid(_stealNet_io_connSS_38_data_availableTask_valid),
		.io_connSS_38_data_availableTask_bits(_stealNet_io_connSS_38_data_availableTask_bits),
		.io_connSS_38_data_qOutTask_ready(_stealNet_io_connSS_38_data_qOutTask_ready),
		.io_connSS_38_data_qOutTask_valid(_stealServers_20_io_connNetwork_data_qOutTask_valid),
		.io_connSS_38_data_qOutTask_bits(_stealServers_20_io_connNetwork_data_qOutTask_bits),
		.io_connSS_39_ctrl_serveStealReq_valid(_stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_39_ctrl_serveStealReq_ready(_stealNet_io_connSS_39_ctrl_serveStealReq_ready),
		.io_connSS_39_ctrl_stealReq_valid(_stealServers_21_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_39_ctrl_stealReq_ready(_stealNet_io_connSS_39_ctrl_stealReq_ready),
		.io_connSS_39_data_availableTask_ready(_stealServers_21_io_connNetwork_data_availableTask_ready),
		.io_connSS_39_data_availableTask_valid(_stealNet_io_connSS_39_data_availableTask_valid),
		.io_connSS_39_data_availableTask_bits(_stealNet_io_connSS_39_data_availableTask_bits),
		.io_connSS_39_data_qOutTask_ready(_stealNet_io_connSS_39_data_qOutTask_ready),
		.io_connSS_39_data_qOutTask_valid(_stealServers_21_io_connNetwork_data_qOutTask_valid),
		.io_connSS_39_data_qOutTask_bits(_stealServers_21_io_connNetwork_data_qOutTask_bits),
		.io_connSS_40_ctrl_serveStealReq_valid(_stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_40_ctrl_serveStealReq_ready(_stealNet_io_connSS_40_ctrl_serveStealReq_ready),
		.io_connSS_40_ctrl_stealReq_valid(_stealServers_22_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_40_ctrl_stealReq_ready(_stealNet_io_connSS_40_ctrl_stealReq_ready),
		.io_connSS_40_data_availableTask_ready(_stealServers_22_io_connNetwork_data_availableTask_ready),
		.io_connSS_40_data_availableTask_valid(_stealNet_io_connSS_40_data_availableTask_valid),
		.io_connSS_40_data_availableTask_bits(_stealNet_io_connSS_40_data_availableTask_bits),
		.io_connSS_40_data_qOutTask_ready(_stealNet_io_connSS_40_data_qOutTask_ready),
		.io_connSS_40_data_qOutTask_valid(_stealServers_22_io_connNetwork_data_qOutTask_valid),
		.io_connSS_40_data_qOutTask_bits(_stealServers_22_io_connNetwork_data_qOutTask_bits),
		.io_connSS_41_ctrl_serveStealReq_valid(_stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_41_ctrl_serveStealReq_ready(_stealNet_io_connSS_41_ctrl_serveStealReq_ready),
		.io_connSS_41_ctrl_stealReq_valid(_stealServers_23_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_41_ctrl_stealReq_ready(_stealNet_io_connSS_41_ctrl_stealReq_ready),
		.io_connSS_41_data_availableTask_ready(_stealServers_23_io_connNetwork_data_availableTask_ready),
		.io_connSS_41_data_availableTask_valid(_stealNet_io_connSS_41_data_availableTask_valid),
		.io_connSS_41_data_availableTask_bits(_stealNet_io_connSS_41_data_availableTask_bits),
		.io_connSS_41_data_qOutTask_ready(_stealNet_io_connSS_41_data_qOutTask_ready),
		.io_connSS_41_data_qOutTask_valid(_stealServers_23_io_connNetwork_data_qOutTask_valid),
		.io_connSS_41_data_qOutTask_bits(_stealServers_23_io_connNetwork_data_qOutTask_bits),
		.io_connSS_42_ctrl_serveStealReq_valid(_stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_42_ctrl_serveStealReq_ready(_stealNet_io_connSS_42_ctrl_serveStealReq_ready),
		.io_connSS_42_ctrl_stealReq_valid(_stealServers_24_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_42_ctrl_stealReq_ready(_stealNet_io_connSS_42_ctrl_stealReq_ready),
		.io_connSS_42_data_availableTask_ready(_stealServers_24_io_connNetwork_data_availableTask_ready),
		.io_connSS_42_data_availableTask_valid(_stealNet_io_connSS_42_data_availableTask_valid),
		.io_connSS_42_data_availableTask_bits(_stealNet_io_connSS_42_data_availableTask_bits),
		.io_connSS_42_data_qOutTask_ready(_stealNet_io_connSS_42_data_qOutTask_ready),
		.io_connSS_42_data_qOutTask_valid(_stealServers_24_io_connNetwork_data_qOutTask_valid),
		.io_connSS_42_data_qOutTask_bits(_stealServers_24_io_connNetwork_data_qOutTask_bits),
		.io_connSS_43_ctrl_serveStealReq_valid(_stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_43_ctrl_serveStealReq_ready(_stealNet_io_connSS_43_ctrl_serveStealReq_ready),
		.io_connSS_43_ctrl_stealReq_valid(_stealServers_25_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_43_ctrl_stealReq_ready(_stealNet_io_connSS_43_ctrl_stealReq_ready),
		.io_connSS_43_data_availableTask_ready(_stealServers_25_io_connNetwork_data_availableTask_ready),
		.io_connSS_43_data_availableTask_valid(_stealNet_io_connSS_43_data_availableTask_valid),
		.io_connSS_43_data_availableTask_bits(_stealNet_io_connSS_43_data_availableTask_bits),
		.io_connSS_43_data_qOutTask_ready(_stealNet_io_connSS_43_data_qOutTask_ready),
		.io_connSS_43_data_qOutTask_valid(_stealServers_25_io_connNetwork_data_qOutTask_valid),
		.io_connSS_43_data_qOutTask_bits(_stealServers_25_io_connNetwork_data_qOutTask_bits),
		.io_connSS_44_ctrl_serveStealReq_valid(_stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_44_ctrl_serveStealReq_ready(_stealNet_io_connSS_44_ctrl_serveStealReq_ready),
		.io_connSS_44_ctrl_stealReq_valid(_stealServers_26_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_44_ctrl_stealReq_ready(_stealNet_io_connSS_44_ctrl_stealReq_ready),
		.io_connSS_44_data_availableTask_ready(_stealServers_26_io_connNetwork_data_availableTask_ready),
		.io_connSS_44_data_availableTask_valid(_stealNet_io_connSS_44_data_availableTask_valid),
		.io_connSS_44_data_availableTask_bits(_stealNet_io_connSS_44_data_availableTask_bits),
		.io_connSS_44_data_qOutTask_ready(_stealNet_io_connSS_44_data_qOutTask_ready),
		.io_connSS_44_data_qOutTask_valid(_stealServers_26_io_connNetwork_data_qOutTask_valid),
		.io_connSS_44_data_qOutTask_bits(_stealServers_26_io_connNetwork_data_qOutTask_bits),
		.io_connSS_45_ctrl_serveStealReq_valid(_stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_45_ctrl_serveStealReq_ready(_stealNet_io_connSS_45_ctrl_serveStealReq_ready),
		.io_connSS_45_ctrl_stealReq_valid(_stealServers_27_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_45_ctrl_stealReq_ready(_stealNet_io_connSS_45_ctrl_stealReq_ready),
		.io_connSS_45_data_availableTask_ready(_stealServers_27_io_connNetwork_data_availableTask_ready),
		.io_connSS_45_data_availableTask_valid(_stealNet_io_connSS_45_data_availableTask_valid),
		.io_connSS_45_data_availableTask_bits(_stealNet_io_connSS_45_data_availableTask_bits),
		.io_connSS_45_data_qOutTask_ready(_stealNet_io_connSS_45_data_qOutTask_ready),
		.io_connSS_45_data_qOutTask_valid(_stealServers_27_io_connNetwork_data_qOutTask_valid),
		.io_connSS_45_data_qOutTask_bits(_stealServers_27_io_connNetwork_data_qOutTask_bits),
		.io_connSS_46_ctrl_serveStealReq_valid(_stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_46_ctrl_serveStealReq_ready(_stealNet_io_connSS_46_ctrl_serveStealReq_ready),
		.io_connSS_46_ctrl_stealReq_valid(_stealServers_28_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_46_ctrl_stealReq_ready(_stealNet_io_connSS_46_ctrl_stealReq_ready),
		.io_connSS_46_data_availableTask_ready(_stealServers_28_io_connNetwork_data_availableTask_ready),
		.io_connSS_46_data_availableTask_valid(_stealNet_io_connSS_46_data_availableTask_valid),
		.io_connSS_46_data_availableTask_bits(_stealNet_io_connSS_46_data_availableTask_bits),
		.io_connSS_46_data_qOutTask_ready(_stealNet_io_connSS_46_data_qOutTask_ready),
		.io_connSS_46_data_qOutTask_valid(_stealServers_28_io_connNetwork_data_qOutTask_valid),
		.io_connSS_46_data_qOutTask_bits(_stealServers_28_io_connNetwork_data_qOutTask_bits),
		.io_connSS_47_ctrl_serveStealReq_valid(_stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_47_ctrl_serveStealReq_ready(_stealNet_io_connSS_47_ctrl_serveStealReq_ready),
		.io_connSS_47_ctrl_stealReq_valid(_stealServers_29_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_47_ctrl_stealReq_ready(_stealNet_io_connSS_47_ctrl_stealReq_ready),
		.io_connSS_47_data_availableTask_ready(_stealServers_29_io_connNetwork_data_availableTask_ready),
		.io_connSS_47_data_availableTask_valid(_stealNet_io_connSS_47_data_availableTask_valid),
		.io_connSS_47_data_availableTask_bits(_stealNet_io_connSS_47_data_availableTask_bits),
		.io_connSS_47_data_qOutTask_ready(_stealNet_io_connSS_47_data_qOutTask_ready),
		.io_connSS_47_data_qOutTask_valid(_stealServers_29_io_connNetwork_data_qOutTask_valid),
		.io_connSS_47_data_qOutTask_bits(_stealServers_29_io_connNetwork_data_qOutTask_bits),
		.io_connSS_48_ctrl_serveStealReq_valid(_stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_48_ctrl_serveStealReq_ready(_stealNet_io_connSS_48_ctrl_serveStealReq_ready),
		.io_connSS_48_ctrl_stealReq_valid(_stealServers_30_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_48_ctrl_stealReq_ready(_stealNet_io_connSS_48_ctrl_stealReq_ready),
		.io_connSS_48_data_availableTask_ready(_stealServers_30_io_connNetwork_data_availableTask_ready),
		.io_connSS_48_data_availableTask_valid(_stealNet_io_connSS_48_data_availableTask_valid),
		.io_connSS_48_data_availableTask_bits(_stealNet_io_connSS_48_data_availableTask_bits),
		.io_connSS_48_data_qOutTask_ready(_stealNet_io_connSS_48_data_qOutTask_ready),
		.io_connSS_48_data_qOutTask_valid(_stealServers_30_io_connNetwork_data_qOutTask_valid),
		.io_connSS_48_data_qOutTask_bits(_stealServers_30_io_connNetwork_data_qOutTask_bits),
		.io_connSS_49_ctrl_serveStealReq_valid(_stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_49_ctrl_serveStealReq_ready(_stealNet_io_connSS_49_ctrl_serveStealReq_ready),
		.io_connSS_49_ctrl_stealReq_valid(_stealServers_31_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_49_ctrl_stealReq_ready(_stealNet_io_connSS_49_ctrl_stealReq_ready),
		.io_connSS_49_data_availableTask_ready(_stealServers_31_io_connNetwork_data_availableTask_ready),
		.io_connSS_49_data_availableTask_valid(_stealNet_io_connSS_49_data_availableTask_valid),
		.io_connSS_49_data_availableTask_bits(_stealNet_io_connSS_49_data_availableTask_bits),
		.io_connSS_49_data_qOutTask_ready(_stealNet_io_connSS_49_data_qOutTask_ready),
		.io_connSS_49_data_qOutTask_valid(_stealServers_31_io_connNetwork_data_qOutTask_valid),
		.io_connSS_49_data_qOutTask_bits(_stealServers_31_io_connNetwork_data_qOutTask_bits),
		.io_connSS_50_ctrl_serveStealReq_valid(_stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_50_ctrl_serveStealReq_ready(_stealNet_io_connSS_50_ctrl_serveStealReq_ready),
		.io_connSS_50_ctrl_stealReq_valid(_stealServers_32_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_50_ctrl_stealReq_ready(_stealNet_io_connSS_50_ctrl_stealReq_ready),
		.io_connSS_50_data_availableTask_ready(_stealServers_32_io_connNetwork_data_availableTask_ready),
		.io_connSS_50_data_availableTask_valid(_stealNet_io_connSS_50_data_availableTask_valid),
		.io_connSS_50_data_availableTask_bits(_stealNet_io_connSS_50_data_availableTask_bits),
		.io_connSS_50_data_qOutTask_ready(_stealNet_io_connSS_50_data_qOutTask_ready),
		.io_connSS_50_data_qOutTask_valid(_stealServers_32_io_connNetwork_data_qOutTask_valid),
		.io_connSS_50_data_qOutTask_bits(_stealServers_32_io_connNetwork_data_qOutTask_bits),
		.io_connSS_51_ctrl_serveStealReq_valid(_stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_51_ctrl_serveStealReq_ready(_stealNet_io_connSS_51_ctrl_serveStealReq_ready),
		.io_connSS_51_ctrl_stealReq_valid(_stealServers_33_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_51_ctrl_stealReq_ready(_stealNet_io_connSS_51_ctrl_stealReq_ready),
		.io_connSS_51_data_availableTask_ready(_stealServers_33_io_connNetwork_data_availableTask_ready),
		.io_connSS_51_data_availableTask_valid(_stealNet_io_connSS_51_data_availableTask_valid),
		.io_connSS_51_data_availableTask_bits(_stealNet_io_connSS_51_data_availableTask_bits),
		.io_connSS_51_data_qOutTask_ready(_stealNet_io_connSS_51_data_qOutTask_ready),
		.io_connSS_51_data_qOutTask_valid(_stealServers_33_io_connNetwork_data_qOutTask_valid),
		.io_connSS_51_data_qOutTask_bits(_stealServers_33_io_connNetwork_data_qOutTask_bits),
		.io_connSS_52_ctrl_serveStealReq_valid(_stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_52_ctrl_serveStealReq_ready(_stealNet_io_connSS_52_ctrl_serveStealReq_ready),
		.io_connSS_52_ctrl_stealReq_valid(_stealServers_34_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_52_ctrl_stealReq_ready(_stealNet_io_connSS_52_ctrl_stealReq_ready),
		.io_connSS_52_data_availableTask_ready(_stealServers_34_io_connNetwork_data_availableTask_ready),
		.io_connSS_52_data_availableTask_valid(_stealNet_io_connSS_52_data_availableTask_valid),
		.io_connSS_52_data_availableTask_bits(_stealNet_io_connSS_52_data_availableTask_bits),
		.io_connSS_52_data_qOutTask_ready(_stealNet_io_connSS_52_data_qOutTask_ready),
		.io_connSS_52_data_qOutTask_valid(_stealServers_34_io_connNetwork_data_qOutTask_valid),
		.io_connSS_52_data_qOutTask_bits(_stealServers_34_io_connNetwork_data_qOutTask_bits),
		.io_connSS_53_ctrl_serveStealReq_valid(_stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_53_ctrl_serveStealReq_ready(_stealNet_io_connSS_53_ctrl_serveStealReq_ready),
		.io_connSS_53_ctrl_stealReq_valid(_stealServers_35_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_53_ctrl_stealReq_ready(_stealNet_io_connSS_53_ctrl_stealReq_ready),
		.io_connSS_53_data_availableTask_ready(_stealServers_35_io_connNetwork_data_availableTask_ready),
		.io_connSS_53_data_availableTask_valid(_stealNet_io_connSS_53_data_availableTask_valid),
		.io_connSS_53_data_availableTask_bits(_stealNet_io_connSS_53_data_availableTask_bits),
		.io_connSS_53_data_qOutTask_ready(_stealNet_io_connSS_53_data_qOutTask_ready),
		.io_connSS_53_data_qOutTask_valid(_stealServers_35_io_connNetwork_data_qOutTask_valid),
		.io_connSS_53_data_qOutTask_bits(_stealServers_35_io_connNetwork_data_qOutTask_bits),
		.io_connSS_54_ctrl_serveStealReq_valid(_stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_54_ctrl_serveStealReq_ready(_stealNet_io_connSS_54_ctrl_serveStealReq_ready),
		.io_connSS_54_ctrl_stealReq_valid(_stealServers_36_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_54_ctrl_stealReq_ready(_stealNet_io_connSS_54_ctrl_stealReq_ready),
		.io_connSS_54_data_availableTask_ready(_stealServers_36_io_connNetwork_data_availableTask_ready),
		.io_connSS_54_data_availableTask_valid(_stealNet_io_connSS_54_data_availableTask_valid),
		.io_connSS_54_data_availableTask_bits(_stealNet_io_connSS_54_data_availableTask_bits),
		.io_connSS_54_data_qOutTask_ready(_stealNet_io_connSS_54_data_qOutTask_ready),
		.io_connSS_54_data_qOutTask_valid(_stealServers_36_io_connNetwork_data_qOutTask_valid),
		.io_connSS_54_data_qOutTask_bits(_stealServers_36_io_connNetwork_data_qOutTask_bits),
		.io_connSS_55_ctrl_serveStealReq_valid(_stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_55_ctrl_serveStealReq_ready(_stealNet_io_connSS_55_ctrl_serveStealReq_ready),
		.io_connSS_55_ctrl_stealReq_valid(_stealServers_37_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_55_ctrl_stealReq_ready(_stealNet_io_connSS_55_ctrl_stealReq_ready),
		.io_connSS_55_data_availableTask_ready(_stealServers_37_io_connNetwork_data_availableTask_ready),
		.io_connSS_55_data_availableTask_valid(_stealNet_io_connSS_55_data_availableTask_valid),
		.io_connSS_55_data_availableTask_bits(_stealNet_io_connSS_55_data_availableTask_bits),
		.io_connSS_55_data_qOutTask_ready(_stealNet_io_connSS_55_data_qOutTask_ready),
		.io_connSS_55_data_qOutTask_valid(_stealServers_37_io_connNetwork_data_qOutTask_valid),
		.io_connSS_55_data_qOutTask_bits(_stealServers_37_io_connNetwork_data_qOutTask_bits),
		.io_connSS_56_ctrl_serveStealReq_valid(_stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_56_ctrl_serveStealReq_ready(_stealNet_io_connSS_56_ctrl_serveStealReq_ready),
		.io_connSS_56_ctrl_stealReq_valid(_stealServers_38_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_56_ctrl_stealReq_ready(_stealNet_io_connSS_56_ctrl_stealReq_ready),
		.io_connSS_56_data_availableTask_ready(_stealServers_38_io_connNetwork_data_availableTask_ready),
		.io_connSS_56_data_availableTask_valid(_stealNet_io_connSS_56_data_availableTask_valid),
		.io_connSS_56_data_availableTask_bits(_stealNet_io_connSS_56_data_availableTask_bits),
		.io_connSS_56_data_qOutTask_ready(_stealNet_io_connSS_56_data_qOutTask_ready),
		.io_connSS_56_data_qOutTask_valid(_stealServers_38_io_connNetwork_data_qOutTask_valid),
		.io_connSS_56_data_qOutTask_bits(_stealServers_38_io_connNetwork_data_qOutTask_bits),
		.io_connSS_57_ctrl_serveStealReq_valid(_stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_57_ctrl_serveStealReq_ready(_stealNet_io_connSS_57_ctrl_serveStealReq_ready),
		.io_connSS_57_ctrl_stealReq_valid(_stealServers_39_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_57_ctrl_stealReq_ready(_stealNet_io_connSS_57_ctrl_stealReq_ready),
		.io_connSS_57_data_availableTask_ready(_stealServers_39_io_connNetwork_data_availableTask_ready),
		.io_connSS_57_data_availableTask_valid(_stealNet_io_connSS_57_data_availableTask_valid),
		.io_connSS_57_data_availableTask_bits(_stealNet_io_connSS_57_data_availableTask_bits),
		.io_connSS_57_data_qOutTask_ready(_stealNet_io_connSS_57_data_qOutTask_ready),
		.io_connSS_57_data_qOutTask_valid(_stealServers_39_io_connNetwork_data_qOutTask_valid),
		.io_connSS_57_data_qOutTask_bits(_stealServers_39_io_connNetwork_data_qOutTask_bits),
		.io_connSS_58_ctrl_serveStealReq_valid(_stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_58_ctrl_serveStealReq_ready(_stealNet_io_connSS_58_ctrl_serveStealReq_ready),
		.io_connSS_58_ctrl_stealReq_valid(_stealServers_40_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_58_ctrl_stealReq_ready(_stealNet_io_connSS_58_ctrl_stealReq_ready),
		.io_connSS_58_data_availableTask_ready(_stealServers_40_io_connNetwork_data_availableTask_ready),
		.io_connSS_58_data_availableTask_valid(_stealNet_io_connSS_58_data_availableTask_valid),
		.io_connSS_58_data_availableTask_bits(_stealNet_io_connSS_58_data_availableTask_bits),
		.io_connSS_58_data_qOutTask_ready(_stealNet_io_connSS_58_data_qOutTask_ready),
		.io_connSS_58_data_qOutTask_valid(_stealServers_40_io_connNetwork_data_qOutTask_valid),
		.io_connSS_58_data_qOutTask_bits(_stealServers_40_io_connNetwork_data_qOutTask_bits),
		.io_connSS_59_ctrl_serveStealReq_valid(_stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_59_ctrl_serveStealReq_ready(_stealNet_io_connSS_59_ctrl_serveStealReq_ready),
		.io_connSS_59_ctrl_stealReq_valid(_stealServers_41_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_59_ctrl_stealReq_ready(_stealNet_io_connSS_59_ctrl_stealReq_ready),
		.io_connSS_59_data_availableTask_ready(_stealServers_41_io_connNetwork_data_availableTask_ready),
		.io_connSS_59_data_availableTask_valid(_stealNet_io_connSS_59_data_availableTask_valid),
		.io_connSS_59_data_availableTask_bits(_stealNet_io_connSS_59_data_availableTask_bits),
		.io_connSS_59_data_qOutTask_ready(_stealNet_io_connSS_59_data_qOutTask_ready),
		.io_connSS_59_data_qOutTask_valid(_stealServers_41_io_connNetwork_data_qOutTask_valid),
		.io_connSS_59_data_qOutTask_bits(_stealServers_41_io_connNetwork_data_qOutTask_bits),
		.io_connSS_60_ctrl_serveStealReq_valid(_stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_60_ctrl_serveStealReq_ready(_stealNet_io_connSS_60_ctrl_serveStealReq_ready),
		.io_connSS_60_ctrl_stealReq_valid(_stealServers_42_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_60_ctrl_stealReq_ready(_stealNet_io_connSS_60_ctrl_stealReq_ready),
		.io_connSS_60_data_availableTask_ready(_stealServers_42_io_connNetwork_data_availableTask_ready),
		.io_connSS_60_data_availableTask_valid(_stealNet_io_connSS_60_data_availableTask_valid),
		.io_connSS_60_data_availableTask_bits(_stealNet_io_connSS_60_data_availableTask_bits),
		.io_connSS_60_data_qOutTask_ready(_stealNet_io_connSS_60_data_qOutTask_ready),
		.io_connSS_60_data_qOutTask_valid(_stealServers_42_io_connNetwork_data_qOutTask_valid),
		.io_connSS_60_data_qOutTask_bits(_stealServers_42_io_connNetwork_data_qOutTask_bits),
		.io_connSS_61_ctrl_serveStealReq_valid(_stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_61_ctrl_serveStealReq_ready(_stealNet_io_connSS_61_ctrl_serveStealReq_ready),
		.io_connSS_61_ctrl_stealReq_valid(_stealServers_43_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_61_ctrl_stealReq_ready(_stealNet_io_connSS_61_ctrl_stealReq_ready),
		.io_connSS_61_data_availableTask_ready(_stealServers_43_io_connNetwork_data_availableTask_ready),
		.io_connSS_61_data_availableTask_valid(_stealNet_io_connSS_61_data_availableTask_valid),
		.io_connSS_61_data_availableTask_bits(_stealNet_io_connSS_61_data_availableTask_bits),
		.io_connSS_61_data_qOutTask_ready(_stealNet_io_connSS_61_data_qOutTask_ready),
		.io_connSS_61_data_qOutTask_valid(_stealServers_43_io_connNetwork_data_qOutTask_valid),
		.io_connSS_61_data_qOutTask_bits(_stealServers_43_io_connNetwork_data_qOutTask_bits),
		.io_connSS_62_ctrl_serveStealReq_valid(_stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_62_ctrl_serveStealReq_ready(_stealNet_io_connSS_62_ctrl_serveStealReq_ready),
		.io_connSS_62_ctrl_stealReq_valid(_stealServers_44_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_62_ctrl_stealReq_ready(_stealNet_io_connSS_62_ctrl_stealReq_ready),
		.io_connSS_62_data_availableTask_ready(_stealServers_44_io_connNetwork_data_availableTask_ready),
		.io_connSS_62_data_availableTask_valid(_stealNet_io_connSS_62_data_availableTask_valid),
		.io_connSS_62_data_availableTask_bits(_stealNet_io_connSS_62_data_availableTask_bits),
		.io_connSS_62_data_qOutTask_ready(_stealNet_io_connSS_62_data_qOutTask_ready),
		.io_connSS_62_data_qOutTask_valid(_stealServers_44_io_connNetwork_data_qOutTask_valid),
		.io_connSS_62_data_qOutTask_bits(_stealServers_44_io_connNetwork_data_qOutTask_bits),
		.io_connSS_63_ctrl_serveStealReq_valid(_stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_63_ctrl_serveStealReq_ready(_stealNet_io_connSS_63_ctrl_serveStealReq_ready),
		.io_connSS_63_ctrl_stealReq_valid(_stealServers_45_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_63_ctrl_stealReq_ready(_stealNet_io_connSS_63_ctrl_stealReq_ready),
		.io_connSS_63_data_availableTask_ready(_stealServers_45_io_connNetwork_data_availableTask_ready),
		.io_connSS_63_data_availableTask_valid(_stealNet_io_connSS_63_data_availableTask_valid),
		.io_connSS_63_data_availableTask_bits(_stealNet_io_connSS_63_data_availableTask_bits),
		.io_connSS_63_data_qOutTask_ready(_stealNet_io_connSS_63_data_qOutTask_ready),
		.io_connSS_63_data_qOutTask_valid(_stealServers_45_io_connNetwork_data_qOutTask_valid),
		.io_connSS_63_data_qOutTask_bits(_stealServers_45_io_connNetwork_data_qOutTask_bits),
		.io_connSS_64_ctrl_serveStealReq_valid(_stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_64_ctrl_serveStealReq_ready(_stealNet_io_connSS_64_ctrl_serveStealReq_ready),
		.io_connSS_64_ctrl_stealReq_valid(_stealServers_46_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_64_ctrl_stealReq_ready(_stealNet_io_connSS_64_ctrl_stealReq_ready),
		.io_connSS_64_data_availableTask_ready(_stealServers_46_io_connNetwork_data_availableTask_ready),
		.io_connSS_64_data_availableTask_valid(_stealNet_io_connSS_64_data_availableTask_valid),
		.io_connSS_64_data_availableTask_bits(_stealNet_io_connSS_64_data_availableTask_bits),
		.io_connSS_64_data_qOutTask_ready(_stealNet_io_connSS_64_data_qOutTask_ready),
		.io_connSS_64_data_qOutTask_valid(_stealServers_46_io_connNetwork_data_qOutTask_valid),
		.io_connSS_64_data_qOutTask_bits(_stealServers_46_io_connNetwork_data_qOutTask_bits),
		.io_connSS_65_ctrl_serveStealReq_valid(_stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_65_ctrl_serveStealReq_ready(_stealNet_io_connSS_65_ctrl_serveStealReq_ready),
		.io_connSS_65_ctrl_stealReq_valid(_stealServers_47_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_65_ctrl_stealReq_ready(_stealNet_io_connSS_65_ctrl_stealReq_ready),
		.io_connSS_65_data_availableTask_ready(_stealServers_47_io_connNetwork_data_availableTask_ready),
		.io_connSS_65_data_availableTask_valid(_stealNet_io_connSS_65_data_availableTask_valid),
		.io_connSS_65_data_availableTask_bits(_stealNet_io_connSS_65_data_availableTask_bits),
		.io_connSS_65_data_qOutTask_ready(_stealNet_io_connSS_65_data_qOutTask_ready),
		.io_connSS_65_data_qOutTask_valid(_stealServers_47_io_connNetwork_data_qOutTask_valid),
		.io_connSS_65_data_qOutTask_bits(_stealServers_47_io_connNetwork_data_qOutTask_bits),
		.io_connSS_66_ctrl_serveStealReq_valid(_stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_66_ctrl_serveStealReq_ready(_stealNet_io_connSS_66_ctrl_serveStealReq_ready),
		.io_connSS_66_ctrl_stealReq_valid(_stealServers_48_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_66_ctrl_stealReq_ready(_stealNet_io_connSS_66_ctrl_stealReq_ready),
		.io_connSS_66_data_availableTask_ready(_stealServers_48_io_connNetwork_data_availableTask_ready),
		.io_connSS_66_data_availableTask_valid(_stealNet_io_connSS_66_data_availableTask_valid),
		.io_connSS_66_data_availableTask_bits(_stealNet_io_connSS_66_data_availableTask_bits),
		.io_connSS_66_data_qOutTask_ready(_stealNet_io_connSS_66_data_qOutTask_ready),
		.io_connSS_66_data_qOutTask_valid(_stealServers_48_io_connNetwork_data_qOutTask_valid),
		.io_connSS_66_data_qOutTask_bits(_stealServers_48_io_connNetwork_data_qOutTask_bits),
		.io_connSS_67_ctrl_serveStealReq_valid(_stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_67_ctrl_serveStealReq_ready(_stealNet_io_connSS_67_ctrl_serveStealReq_ready),
		.io_connSS_67_ctrl_stealReq_valid(_stealServers_49_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_67_ctrl_stealReq_ready(_stealNet_io_connSS_67_ctrl_stealReq_ready),
		.io_connSS_67_data_availableTask_ready(_stealServers_49_io_connNetwork_data_availableTask_ready),
		.io_connSS_67_data_availableTask_valid(_stealNet_io_connSS_67_data_availableTask_valid),
		.io_connSS_67_data_availableTask_bits(_stealNet_io_connSS_67_data_availableTask_bits),
		.io_connSS_67_data_qOutTask_ready(_stealNet_io_connSS_67_data_qOutTask_ready),
		.io_connSS_67_data_qOutTask_valid(_stealServers_49_io_connNetwork_data_qOutTask_valid),
		.io_connSS_67_data_qOutTask_bits(_stealServers_49_io_connNetwork_data_qOutTask_bits),
		.io_connSS_68_ctrl_serveStealReq_valid(_stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_68_ctrl_serveStealReq_ready(_stealNet_io_connSS_68_ctrl_serveStealReq_ready),
		.io_connSS_68_ctrl_stealReq_valid(_stealServers_50_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_68_ctrl_stealReq_ready(_stealNet_io_connSS_68_ctrl_stealReq_ready),
		.io_connSS_68_data_availableTask_ready(_stealServers_50_io_connNetwork_data_availableTask_ready),
		.io_connSS_68_data_availableTask_valid(_stealNet_io_connSS_68_data_availableTask_valid),
		.io_connSS_68_data_availableTask_bits(_stealNet_io_connSS_68_data_availableTask_bits),
		.io_connSS_68_data_qOutTask_ready(_stealNet_io_connSS_68_data_qOutTask_ready),
		.io_connSS_68_data_qOutTask_valid(_stealServers_50_io_connNetwork_data_qOutTask_valid),
		.io_connSS_68_data_qOutTask_bits(_stealServers_50_io_connNetwork_data_qOutTask_bits),
		.io_connSS_69_ctrl_serveStealReq_valid(_stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_69_ctrl_serveStealReq_ready(_stealNet_io_connSS_69_ctrl_serveStealReq_ready),
		.io_connSS_69_ctrl_stealReq_valid(_stealServers_51_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_69_ctrl_stealReq_ready(_stealNet_io_connSS_69_ctrl_stealReq_ready),
		.io_connSS_69_data_availableTask_ready(_stealServers_51_io_connNetwork_data_availableTask_ready),
		.io_connSS_69_data_availableTask_valid(_stealNet_io_connSS_69_data_availableTask_valid),
		.io_connSS_69_data_availableTask_bits(_stealNet_io_connSS_69_data_availableTask_bits),
		.io_connSS_69_data_qOutTask_ready(_stealNet_io_connSS_69_data_qOutTask_ready),
		.io_connSS_69_data_qOutTask_valid(_stealServers_51_io_connNetwork_data_qOutTask_valid),
		.io_connSS_69_data_qOutTask_bits(_stealServers_51_io_connNetwork_data_qOutTask_bits),
		.io_connSS_70_ctrl_serveStealReq_valid(_stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_70_ctrl_serveStealReq_ready(_stealNet_io_connSS_70_ctrl_serveStealReq_ready),
		.io_connSS_70_ctrl_stealReq_valid(_stealServers_52_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_70_ctrl_stealReq_ready(_stealNet_io_connSS_70_ctrl_stealReq_ready),
		.io_connSS_70_data_availableTask_ready(_stealServers_52_io_connNetwork_data_availableTask_ready),
		.io_connSS_70_data_availableTask_valid(_stealNet_io_connSS_70_data_availableTask_valid),
		.io_connSS_70_data_availableTask_bits(_stealNet_io_connSS_70_data_availableTask_bits),
		.io_connSS_70_data_qOutTask_ready(_stealNet_io_connSS_70_data_qOutTask_ready),
		.io_connSS_70_data_qOutTask_valid(_stealServers_52_io_connNetwork_data_qOutTask_valid),
		.io_connSS_70_data_qOutTask_bits(_stealServers_52_io_connNetwork_data_qOutTask_bits),
		.io_connSS_71_ctrl_serveStealReq_valid(_stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_71_ctrl_serveStealReq_ready(_stealNet_io_connSS_71_ctrl_serveStealReq_ready),
		.io_connSS_71_ctrl_stealReq_valid(_stealServers_53_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_71_ctrl_stealReq_ready(_stealNet_io_connSS_71_ctrl_stealReq_ready),
		.io_connSS_71_data_availableTask_ready(_stealServers_53_io_connNetwork_data_availableTask_ready),
		.io_connSS_71_data_availableTask_valid(_stealNet_io_connSS_71_data_availableTask_valid),
		.io_connSS_71_data_availableTask_bits(_stealNet_io_connSS_71_data_availableTask_bits),
		.io_connSS_71_data_qOutTask_ready(_stealNet_io_connSS_71_data_qOutTask_ready),
		.io_connSS_71_data_qOutTask_valid(_stealServers_53_io_connNetwork_data_qOutTask_valid),
		.io_connSS_71_data_qOutTask_bits(_stealServers_53_io_connNetwork_data_qOutTask_bits),
		.io_connSS_72_ctrl_serveStealReq_valid(_stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_72_ctrl_serveStealReq_ready(_stealNet_io_connSS_72_ctrl_serveStealReq_ready),
		.io_connSS_72_ctrl_stealReq_valid(_stealServers_54_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_72_ctrl_stealReq_ready(_stealNet_io_connSS_72_ctrl_stealReq_ready),
		.io_connSS_72_data_availableTask_ready(_stealServers_54_io_connNetwork_data_availableTask_ready),
		.io_connSS_72_data_availableTask_valid(_stealNet_io_connSS_72_data_availableTask_valid),
		.io_connSS_72_data_availableTask_bits(_stealNet_io_connSS_72_data_availableTask_bits),
		.io_connSS_72_data_qOutTask_ready(_stealNet_io_connSS_72_data_qOutTask_ready),
		.io_connSS_72_data_qOutTask_valid(_stealServers_54_io_connNetwork_data_qOutTask_valid),
		.io_connSS_72_data_qOutTask_bits(_stealServers_54_io_connNetwork_data_qOutTask_bits),
		.io_connSS_73_ctrl_serveStealReq_valid(_stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_73_ctrl_serveStealReq_ready(_stealNet_io_connSS_73_ctrl_serveStealReq_ready),
		.io_connSS_73_ctrl_stealReq_valid(_stealServers_55_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_73_ctrl_stealReq_ready(_stealNet_io_connSS_73_ctrl_stealReq_ready),
		.io_connSS_73_data_availableTask_ready(_stealServers_55_io_connNetwork_data_availableTask_ready),
		.io_connSS_73_data_availableTask_valid(_stealNet_io_connSS_73_data_availableTask_valid),
		.io_connSS_73_data_availableTask_bits(_stealNet_io_connSS_73_data_availableTask_bits),
		.io_connSS_73_data_qOutTask_ready(_stealNet_io_connSS_73_data_qOutTask_ready),
		.io_connSS_73_data_qOutTask_valid(_stealServers_55_io_connNetwork_data_qOutTask_valid),
		.io_connSS_73_data_qOutTask_bits(_stealServers_55_io_connNetwork_data_qOutTask_bits),
		.io_connSS_74_ctrl_serveStealReq_valid(_stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_74_ctrl_serveStealReq_ready(_stealNet_io_connSS_74_ctrl_serveStealReq_ready),
		.io_connSS_74_ctrl_stealReq_valid(_stealServers_56_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_74_ctrl_stealReq_ready(_stealNet_io_connSS_74_ctrl_stealReq_ready),
		.io_connSS_74_data_availableTask_ready(_stealServers_56_io_connNetwork_data_availableTask_ready),
		.io_connSS_74_data_availableTask_valid(_stealNet_io_connSS_74_data_availableTask_valid),
		.io_connSS_74_data_availableTask_bits(_stealNet_io_connSS_74_data_availableTask_bits),
		.io_connSS_74_data_qOutTask_ready(_stealNet_io_connSS_74_data_qOutTask_ready),
		.io_connSS_74_data_qOutTask_valid(_stealServers_56_io_connNetwork_data_qOutTask_valid),
		.io_connSS_74_data_qOutTask_bits(_stealServers_56_io_connNetwork_data_qOutTask_bits),
		.io_connSS_75_ctrl_serveStealReq_valid(_stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_75_ctrl_serveStealReq_ready(_stealNet_io_connSS_75_ctrl_serveStealReq_ready),
		.io_connSS_75_ctrl_stealReq_valid(_stealServers_57_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_75_ctrl_stealReq_ready(_stealNet_io_connSS_75_ctrl_stealReq_ready),
		.io_connSS_75_data_availableTask_ready(_stealServers_57_io_connNetwork_data_availableTask_ready),
		.io_connSS_75_data_availableTask_valid(_stealNet_io_connSS_75_data_availableTask_valid),
		.io_connSS_75_data_availableTask_bits(_stealNet_io_connSS_75_data_availableTask_bits),
		.io_connSS_75_data_qOutTask_ready(_stealNet_io_connSS_75_data_qOutTask_ready),
		.io_connSS_75_data_qOutTask_valid(_stealServers_57_io_connNetwork_data_qOutTask_valid),
		.io_connSS_75_data_qOutTask_bits(_stealServers_57_io_connNetwork_data_qOutTask_bits),
		.io_connSS_76_ctrl_serveStealReq_valid(_stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_76_ctrl_serveStealReq_ready(_stealNet_io_connSS_76_ctrl_serveStealReq_ready),
		.io_connSS_76_ctrl_stealReq_valid(_stealServers_58_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_76_ctrl_stealReq_ready(_stealNet_io_connSS_76_ctrl_stealReq_ready),
		.io_connSS_76_data_availableTask_ready(_stealServers_58_io_connNetwork_data_availableTask_ready),
		.io_connSS_76_data_availableTask_valid(_stealNet_io_connSS_76_data_availableTask_valid),
		.io_connSS_76_data_availableTask_bits(_stealNet_io_connSS_76_data_availableTask_bits),
		.io_connSS_76_data_qOutTask_ready(_stealNet_io_connSS_76_data_qOutTask_ready),
		.io_connSS_76_data_qOutTask_valid(_stealServers_58_io_connNetwork_data_qOutTask_valid),
		.io_connSS_76_data_qOutTask_bits(_stealServers_58_io_connNetwork_data_qOutTask_bits),
		.io_connSS_77_ctrl_serveStealReq_valid(_stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_77_ctrl_serveStealReq_ready(_stealNet_io_connSS_77_ctrl_serveStealReq_ready),
		.io_connSS_77_ctrl_stealReq_valid(_stealServers_59_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_77_ctrl_stealReq_ready(_stealNet_io_connSS_77_ctrl_stealReq_ready),
		.io_connSS_77_data_availableTask_ready(_stealServers_59_io_connNetwork_data_availableTask_ready),
		.io_connSS_77_data_availableTask_valid(_stealNet_io_connSS_77_data_availableTask_valid),
		.io_connSS_77_data_availableTask_bits(_stealNet_io_connSS_77_data_availableTask_bits),
		.io_connSS_77_data_qOutTask_ready(_stealNet_io_connSS_77_data_qOutTask_ready),
		.io_connSS_77_data_qOutTask_valid(_stealServers_59_io_connNetwork_data_qOutTask_valid),
		.io_connSS_77_data_qOutTask_bits(_stealServers_59_io_connNetwork_data_qOutTask_bits),
		.io_connSS_78_ctrl_serveStealReq_valid(_stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_78_ctrl_serveStealReq_ready(_stealNet_io_connSS_78_ctrl_serveStealReq_ready),
		.io_connSS_78_ctrl_stealReq_valid(_stealServers_60_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_78_ctrl_stealReq_ready(_stealNet_io_connSS_78_ctrl_stealReq_ready),
		.io_connSS_78_data_availableTask_ready(_stealServers_60_io_connNetwork_data_availableTask_ready),
		.io_connSS_78_data_availableTask_valid(_stealNet_io_connSS_78_data_availableTask_valid),
		.io_connSS_78_data_availableTask_bits(_stealNet_io_connSS_78_data_availableTask_bits),
		.io_connSS_78_data_qOutTask_ready(_stealNet_io_connSS_78_data_qOutTask_ready),
		.io_connSS_78_data_qOutTask_valid(_stealServers_60_io_connNetwork_data_qOutTask_valid),
		.io_connSS_78_data_qOutTask_bits(_stealServers_60_io_connNetwork_data_qOutTask_bits),
		.io_connSS_79_ctrl_serveStealReq_valid(_stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_79_ctrl_serveStealReq_ready(_stealNet_io_connSS_79_ctrl_serveStealReq_ready),
		.io_connSS_79_ctrl_stealReq_valid(_stealServers_61_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_79_ctrl_stealReq_ready(_stealNet_io_connSS_79_ctrl_stealReq_ready),
		.io_connSS_79_data_availableTask_ready(_stealServers_61_io_connNetwork_data_availableTask_ready),
		.io_connSS_79_data_availableTask_valid(_stealNet_io_connSS_79_data_availableTask_valid),
		.io_connSS_79_data_availableTask_bits(_stealNet_io_connSS_79_data_availableTask_bits),
		.io_connSS_79_data_qOutTask_ready(_stealNet_io_connSS_79_data_qOutTask_ready),
		.io_connSS_79_data_qOutTask_valid(_stealServers_61_io_connNetwork_data_qOutTask_valid),
		.io_connSS_79_data_qOutTask_bits(_stealServers_61_io_connNetwork_data_qOutTask_bits),
		.io_connSS_80_ctrl_serveStealReq_valid(_stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_80_ctrl_serveStealReq_ready(_stealNet_io_connSS_80_ctrl_serveStealReq_ready),
		.io_connSS_80_ctrl_stealReq_valid(_stealServers_62_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_80_ctrl_stealReq_ready(_stealNet_io_connSS_80_ctrl_stealReq_ready),
		.io_connSS_80_data_availableTask_ready(_stealServers_62_io_connNetwork_data_availableTask_ready),
		.io_connSS_80_data_availableTask_valid(_stealNet_io_connSS_80_data_availableTask_valid),
		.io_connSS_80_data_availableTask_bits(_stealNet_io_connSS_80_data_availableTask_bits),
		.io_connSS_80_data_qOutTask_ready(_stealNet_io_connSS_80_data_qOutTask_ready),
		.io_connSS_80_data_qOutTask_valid(_stealServers_62_io_connNetwork_data_qOutTask_valid),
		.io_connSS_80_data_qOutTask_bits(_stealServers_62_io_connNetwork_data_qOutTask_bits),
		.io_connSS_81_ctrl_serveStealReq_valid(_stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_81_ctrl_serveStealReq_ready(_stealNet_io_connSS_81_ctrl_serveStealReq_ready),
		.io_connSS_81_ctrl_stealReq_valid(_stealServers_63_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_81_ctrl_stealReq_ready(_stealNet_io_connSS_81_ctrl_stealReq_ready),
		.io_connSS_81_data_availableTask_ready(_stealServers_63_io_connNetwork_data_availableTask_ready),
		.io_connSS_81_data_availableTask_valid(_stealNet_io_connSS_81_data_availableTask_valid),
		.io_connSS_81_data_availableTask_bits(_stealNet_io_connSS_81_data_availableTask_bits),
		.io_connSS_81_data_qOutTask_ready(_stealNet_io_connSS_81_data_qOutTask_ready),
		.io_connSS_81_data_qOutTask_valid(_stealServers_63_io_connNetwork_data_qOutTask_valid),
		.io_connSS_81_data_qOutTask_bits(_stealServers_63_io_connNetwork_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(io_ntwDataUnitOccupancyVSS_0),
		.io_ntwDataUnitOccupancyVSS_1(io_ntwDataUnitOccupancyVSS_1)
	);
	SchedulerClient_64 stealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_0_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_1_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_2(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_2_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_3(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_3_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_4(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_4_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_5(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_5_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_6(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_6_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_7(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_7_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_8(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_8_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_9(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_9_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_10(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_10_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_11(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_11_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_12(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_12_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_13(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_13_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_14(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_14_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_15(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_33_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_33_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_33_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_33_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_33_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_15_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_16(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_34_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_16_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_34_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_16_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_34_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_34_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_34_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_16_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_16_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_16_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_16_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_16_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_16_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_16_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_16_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_16_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_17(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_35_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_17_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_35_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_17_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_35_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_35_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_35_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_17_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_17_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_17_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_17_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_17_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_17_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_17_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_17_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_17_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_18(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_36_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_18_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_36_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_18_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_36_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_36_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_36_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_18_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_18_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_18_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_18_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_18_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_18_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_18_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_18_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_18_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_19(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_37_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_19_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_37_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_19_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_37_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_37_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_37_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_19_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_19_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_19_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_19_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_19_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_19_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_19_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_19_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_19_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_20(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_38_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_20_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_38_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_20_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_38_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_38_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_38_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_20_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_20_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_20_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_20_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_20_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_20_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_20_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_20_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_20_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_21(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_39_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_21_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_39_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_21_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_39_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_39_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_39_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_21_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_21_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_21_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_21_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_21_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_21_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_21_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_21_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_21_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_22(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_40_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_22_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_40_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_22_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_40_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_40_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_40_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_22_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_22_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_22_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_22_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_22_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_22_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_22_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_22_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_22_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_23(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_41_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_23_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_41_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_23_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_41_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_41_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_41_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_23_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_23_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_23_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_23_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_23_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_23_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_23_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_23_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_23_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_24(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_42_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_24_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_42_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_24_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_42_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_42_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_42_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_24_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_24_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_24_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_24_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_24_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_24_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_24_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_24_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_24_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_25(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_43_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_25_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_43_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_25_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_43_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_43_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_43_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_25_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_25_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_25_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_25_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_25_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_25_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_25_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_25_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_25_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_26(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_44_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_26_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_44_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_26_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_44_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_44_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_44_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_26_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_26_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_26_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_26_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_26_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_26_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_26_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_26_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_26_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_27(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_45_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_27_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_45_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_27_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_45_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_45_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_45_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_27_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_27_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_27_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_27_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_27_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_27_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_27_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_27_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_27_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_28(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_46_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_28_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_46_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_28_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_46_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_46_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_46_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_28_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_28_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_28_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_28_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_28_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_28_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_28_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_28_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_28_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_29(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_47_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_29_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_47_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_29_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_47_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_47_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_47_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_29_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_29_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_29_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_29_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_29_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_29_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_29_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_29_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_29_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_30(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_48_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_30_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_48_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_30_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_48_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_48_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_48_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_30_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_30_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_30_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_30_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_30_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_30_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_30_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_30_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_30_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_31(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_49_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_31_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_49_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_31_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_49_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_49_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_49_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_31_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_31_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_31_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_31_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_31_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_31_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_31_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_31_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_31_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_32(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_50_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_32_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_50_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_32_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_50_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_50_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_50_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_32_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_32_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_32_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_32_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_32_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_32_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_32_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_32_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_32_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_33(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_51_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_33_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_51_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_33_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_51_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_51_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_51_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_33_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_33_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_33_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_33_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_33_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_33_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_33_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_33_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_33_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_34(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_52_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_34_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_52_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_34_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_52_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_52_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_52_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_34_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_34_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_34_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_34_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_34_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_34_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_34_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_34_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_34_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_35(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_53_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_35_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_53_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_35_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_53_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_53_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_53_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_35_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_35_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_35_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_35_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_35_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_35_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_35_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_35_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_35_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_36(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_54_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_36_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_54_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_36_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_54_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_54_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_54_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_36_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_36_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_36_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_36_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_36_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_36_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_36_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_36_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_36_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_37(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_55_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_37_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_55_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_37_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_55_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_55_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_55_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_37_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_37_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_37_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_37_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_37_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_37_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_37_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_37_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_37_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_38(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_56_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_38_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_56_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_38_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_56_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_56_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_56_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_38_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_38_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_38_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_38_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_38_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_38_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_38_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_38_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_38_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_39(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_57_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_39_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_57_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_39_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_57_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_57_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_57_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_39_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_39_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_39_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_39_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_39_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_39_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_39_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_39_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_39_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_40(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_58_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_40_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_58_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_40_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_58_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_58_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_58_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_40_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_40_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_40_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_40_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_40_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_40_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_40_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_40_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_40_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_41(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_59_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_41_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_59_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_41_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_59_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_59_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_59_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_41_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_41_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_41_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_41_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_41_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_41_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_41_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_41_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_41_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_42(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_60_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_42_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_60_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_42_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_60_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_60_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_60_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_42_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_42_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_42_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_42_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_42_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_42_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_42_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_42_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_42_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_43(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_61_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_43_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_61_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_43_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_61_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_61_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_61_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_43_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_43_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_43_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_43_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_43_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_43_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_43_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_43_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_43_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_44(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_62_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_44_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_62_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_44_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_62_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_62_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_62_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_44_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_44_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_44_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_44_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_44_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_44_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_44_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_44_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_44_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_45(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_63_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_45_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_63_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_45_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_63_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_63_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_63_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_45_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_45_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_45_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_45_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_45_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_45_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_45_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_45_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_45_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_46(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_64_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_46_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_64_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_46_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_64_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_64_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_64_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_46_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_46_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_46_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_46_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_46_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_46_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_46_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_46_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_46_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_47(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_65_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_47_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_65_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_47_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_65_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_65_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_65_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_47_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_47_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_47_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_47_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_47_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_47_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_47_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_47_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_47_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_48(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_66_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_48_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_66_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_48_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_66_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_66_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_66_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_48_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_48_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_48_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_48_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_48_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_48_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_48_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_48_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_48_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_49(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_67_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_49_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_67_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_49_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_67_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_67_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_67_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_49_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_49_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_49_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_49_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_49_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_49_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_49_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_49_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_49_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_50(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_68_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_50_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_68_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_50_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_68_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_68_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_68_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_50_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_50_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_50_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_50_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_50_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_50_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_50_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_50_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_50_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_51(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_69_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_51_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_69_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_51_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_69_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_69_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_69_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_51_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_51_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_51_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_51_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_51_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_51_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_51_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_51_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_51_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_52(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_70_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_52_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_70_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_52_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_70_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_70_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_70_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_52_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_52_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_52_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_52_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_52_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_52_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_52_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_52_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_52_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_53(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_71_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_53_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_71_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_53_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_71_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_71_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_71_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_53_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_53_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_53_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_53_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_53_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_53_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_53_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_53_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_53_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_54(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_72_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_54_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_72_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_54_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_72_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_72_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_72_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_54_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_54_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_54_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_54_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_54_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_54_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_54_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_54_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_54_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_55(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_73_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_55_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_73_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_55_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_73_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_73_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_73_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_55_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_55_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_55_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_55_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_55_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_55_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_55_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_55_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_55_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_56(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_74_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_56_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_74_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_56_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_74_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_74_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_74_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_56_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_56_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_56_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_56_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_56_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_56_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_56_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_56_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_56_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_57(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_75_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_57_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_75_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_57_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_75_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_75_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_75_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_57_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_57_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_57_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_57_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_57_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_57_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_57_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_57_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_57_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_58(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_76_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_58_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_76_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_58_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_76_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_76_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_76_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_58_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_58_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_58_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_58_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_58_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_58_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_58_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_58_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_58_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_59(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_77_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_59_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_77_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_59_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_77_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_77_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_77_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_59_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_59_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_59_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_59_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_59_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_59_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_59_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_59_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_59_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_60(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_78_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_60_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_78_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_60_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_78_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_78_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_78_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_60_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_60_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_60_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_60_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_60_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_60_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_60_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_60_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_60_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_61(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_79_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_61_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_79_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_61_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_79_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_79_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_79_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_61_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_61_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_61_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_61_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_61_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_61_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_61_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_61_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_61_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_62(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_80_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_62_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_80_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_62_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_80_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_80_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_80_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_62_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_62_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_62_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_62_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_62_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_62_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_62_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_62_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_62_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_63(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_81_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_63_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_81_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_63_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_81_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_81_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_81_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_63_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_63_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_63_io_connVec_1_currLength[3:0]),
		.io_connQ_push_ready(_taskQueues_63_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_63_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_63_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_63_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_63_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_63_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_0(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_0_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_0_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_0_pop_bits),
		.io_connVec_1_currLength(_taskQueues_0_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_1(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_1_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_1_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_1_pop_bits),
		.io_connVec_1_currLength(_taskQueues_1_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_2(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_2_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_2_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_2_pop_bits),
		.io_connVec_1_currLength(_taskQueues_2_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_3(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_3_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_3_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_3_pop_bits),
		.io_connVec_1_currLength(_taskQueues_3_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_4(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_4_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_4_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_4_pop_bits),
		.io_connVec_1_currLength(_taskQueues_4_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_5(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_5_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_5_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_5_pop_bits),
		.io_connVec_1_currLength(_taskQueues_5_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_6(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_6_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_6_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_6_pop_bits),
		.io_connVec_1_currLength(_taskQueues_6_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_7(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_7_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_7_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_7_pop_bits),
		.io_connVec_1_currLength(_taskQueues_7_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_8(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_8_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_8_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_8_pop_bits),
		.io_connVec_1_currLength(_taskQueues_8_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_9(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_9_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_9_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_9_pop_bits),
		.io_connVec_1_currLength(_taskQueues_9_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_10(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_10_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_10_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_10_pop_bits),
		.io_connVec_1_currLength(_taskQueues_10_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_11(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_11_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_11_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_11_pop_bits),
		.io_connVec_1_currLength(_taskQueues_11_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_12(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_12_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_12_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_12_pop_bits),
		.io_connVec_1_currLength(_taskQueues_12_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_13(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_13_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_13_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_13_pop_bits),
		.io_connVec_1_currLength(_taskQueues_13_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_14(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_14_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_14_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_14_pop_bits),
		.io_connVec_1_currLength(_taskQueues_14_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_15(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_15_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_15_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_15_pop_bits),
		.io_connVec_1_currLength(_taskQueues_15_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_16(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_16_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_16_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_16_pop_bits),
		.io_connVec_1_currLength(_taskQueues_16_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_16_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_16_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_16_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_16_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_16_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_16_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_17(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_17_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_17_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_17_pop_bits),
		.io_connVec_1_currLength(_taskQueues_17_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_17_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_17_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_17_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_17_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_17_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_17_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_18(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_18_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_18_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_18_pop_bits),
		.io_connVec_1_currLength(_taskQueues_18_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_18_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_18_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_18_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_18_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_18_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_18_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_19(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_19_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_19_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_19_pop_bits),
		.io_connVec_1_currLength(_taskQueues_19_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_19_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_19_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_19_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_19_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_19_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_19_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_20(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_20_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_20_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_20_pop_bits),
		.io_connVec_1_currLength(_taskQueues_20_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_20_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_20_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_20_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_20_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_20_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_20_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_21(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_21_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_21_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_21_pop_bits),
		.io_connVec_1_currLength(_taskQueues_21_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_21_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_21_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_21_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_21_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_21_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_21_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_22(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_22_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_22_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_22_pop_bits),
		.io_connVec_1_currLength(_taskQueues_22_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_22_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_22_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_22_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_22_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_22_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_22_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_23(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_23_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_23_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_23_pop_bits),
		.io_connVec_1_currLength(_taskQueues_23_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_23_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_23_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_23_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_23_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_23_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_23_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_24(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_24_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_24_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_24_pop_bits),
		.io_connVec_1_currLength(_taskQueues_24_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_24_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_24_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_24_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_24_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_24_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_24_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_25(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_25_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_25_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_25_pop_bits),
		.io_connVec_1_currLength(_taskQueues_25_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_25_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_25_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_25_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_25_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_25_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_25_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_26(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_26_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_26_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_26_pop_bits),
		.io_connVec_1_currLength(_taskQueues_26_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_26_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_26_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_26_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_26_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_26_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_26_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_27(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_27_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_27_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_27_pop_bits),
		.io_connVec_1_currLength(_taskQueues_27_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_27_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_27_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_27_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_27_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_27_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_27_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_28(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_28_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_28_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_28_pop_bits),
		.io_connVec_1_currLength(_taskQueues_28_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_28_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_28_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_28_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_28_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_28_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_28_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_29(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_29_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_29_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_29_pop_bits),
		.io_connVec_1_currLength(_taskQueues_29_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_29_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_29_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_29_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_29_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_29_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_29_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_30(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_30_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_30_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_30_pop_bits),
		.io_connVec_1_currLength(_taskQueues_30_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_30_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_30_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_30_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_30_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_30_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_30_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_31(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_31_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_31_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_31_pop_bits),
		.io_connVec_1_currLength(_taskQueues_31_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_31_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_31_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_31_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_31_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_31_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_31_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_32(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_32_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_32_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_32_pop_bits),
		.io_connVec_1_currLength(_taskQueues_32_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_32_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_32_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_32_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_32_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_32_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_32_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_33(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_33_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_33_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_33_pop_bits),
		.io_connVec_1_currLength(_taskQueues_33_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_33_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_33_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_33_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_33_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_33_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_33_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_34(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_34_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_34_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_34_pop_bits),
		.io_connVec_1_currLength(_taskQueues_34_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_34_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_34_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_34_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_34_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_34_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_34_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_35(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_35_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_35_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_35_pop_bits),
		.io_connVec_1_currLength(_taskQueues_35_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_35_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_35_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_35_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_35_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_35_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_35_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_36(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_36_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_36_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_36_pop_bits),
		.io_connVec_1_currLength(_taskQueues_36_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_36_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_36_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_36_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_36_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_36_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_36_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_37(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_37_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_37_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_37_pop_bits),
		.io_connVec_1_currLength(_taskQueues_37_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_37_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_37_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_37_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_37_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_37_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_37_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_38(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_38_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_38_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_38_pop_bits),
		.io_connVec_1_currLength(_taskQueues_38_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_38_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_38_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_38_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_38_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_38_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_38_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_39(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_39_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_39_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_39_pop_bits),
		.io_connVec_1_currLength(_taskQueues_39_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_39_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_39_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_39_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_39_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_39_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_39_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_40(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_40_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_40_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_40_pop_bits),
		.io_connVec_1_currLength(_taskQueues_40_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_40_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_40_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_40_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_40_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_40_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_40_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_41(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_41_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_41_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_41_pop_bits),
		.io_connVec_1_currLength(_taskQueues_41_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_41_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_41_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_41_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_41_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_41_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_41_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_42(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_42_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_42_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_42_pop_bits),
		.io_connVec_1_currLength(_taskQueues_42_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_42_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_42_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_42_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_42_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_42_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_42_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_43(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_43_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_43_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_43_pop_bits),
		.io_connVec_1_currLength(_taskQueues_43_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_43_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_43_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_43_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_43_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_43_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_43_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_44(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_44_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_44_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_44_pop_bits),
		.io_connVec_1_currLength(_taskQueues_44_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_44_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_44_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_44_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_44_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_44_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_44_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_45(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_45_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_45_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_45_pop_bits),
		.io_connVec_1_currLength(_taskQueues_45_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_45_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_45_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_45_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_45_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_45_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_45_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_46(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_46_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_46_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_46_pop_bits),
		.io_connVec_1_currLength(_taskQueues_46_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_46_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_46_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_46_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_46_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_46_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_46_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_47(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_47_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_47_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_47_pop_bits),
		.io_connVec_1_currLength(_taskQueues_47_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_47_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_47_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_47_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_47_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_47_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_47_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_48(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_48_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_48_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_48_pop_bits),
		.io_connVec_1_currLength(_taskQueues_48_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_48_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_48_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_48_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_48_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_48_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_48_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_49(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_49_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_49_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_49_pop_bits),
		.io_connVec_1_currLength(_taskQueues_49_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_49_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_49_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_49_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_49_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_49_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_49_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_50(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_50_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_50_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_50_pop_bits),
		.io_connVec_1_currLength(_taskQueues_50_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_50_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_50_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_50_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_50_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_50_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_50_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_51(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_51_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_51_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_51_pop_bits),
		.io_connVec_1_currLength(_taskQueues_51_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_51_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_51_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_51_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_51_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_51_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_51_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_52(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_52_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_52_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_52_pop_bits),
		.io_connVec_1_currLength(_taskQueues_52_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_52_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_52_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_52_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_52_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_52_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_52_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_53(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_53_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_53_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_53_pop_bits),
		.io_connVec_1_currLength(_taskQueues_53_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_53_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_53_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_53_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_53_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_53_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_53_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_54(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_54_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_54_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_54_pop_bits),
		.io_connVec_1_currLength(_taskQueues_54_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_54_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_54_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_54_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_54_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_54_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_54_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_55(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_55_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_55_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_55_pop_bits),
		.io_connVec_1_currLength(_taskQueues_55_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_55_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_55_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_55_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_55_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_55_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_55_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_56(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_56_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_56_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_56_pop_bits),
		.io_connVec_1_currLength(_taskQueues_56_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_56_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_56_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_56_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_56_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_56_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_56_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_57(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_57_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_57_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_57_pop_bits),
		.io_connVec_1_currLength(_taskQueues_57_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_57_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_57_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_57_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_57_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_57_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_57_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_58(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_58_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_58_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_58_pop_bits),
		.io_connVec_1_currLength(_taskQueues_58_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_58_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_58_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_58_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_58_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_58_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_58_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_59(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_59_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_59_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_59_pop_bits),
		.io_connVec_1_currLength(_taskQueues_59_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_59_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_59_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_59_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_59_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_59_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_59_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_60(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_60_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_60_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_60_pop_bits),
		.io_connVec_1_currLength(_taskQueues_60_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_60_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_60_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_60_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_60_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_60_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_60_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_61(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_61_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_61_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_61_pop_bits),
		.io_connVec_1_currLength(_taskQueues_61_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_61_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_61_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_61_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_61_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_61_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_61_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_62(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_62_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_62_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_62_pop_bits),
		.io_connVec_1_currLength(_taskQueues_62_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_62_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_62_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_62_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_62_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_62_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_62_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_63(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_63_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_63_pop_valid),
		.io_connVec_0_pop_bits(io_connPE_63_pop_bits),
		.io_connVec_1_currLength(_taskQueues_63_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_63_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_63_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_63_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_63_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_63_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_63_io_connVec_1_pop_bits)
	);
endmodule
module ram_16x256 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [3:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [255:0] R0_data;
	input [3:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [255:0] W0_data;
	reg [255:0] Memory [0:15];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 256'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue16_UInt_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits,
	io_count
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [255:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [255:0] io_deq_bits;
	output wire [4:0] io_count;
	reg [3:0] enq_ptr_value;
	reg [3:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 4'h0;
			deq_ptr_value <= 4'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 4'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 4'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_16x256 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_count = {maybe_full & ptr_match, enq_ptr_value - deq_ptr_value};
endmodule
module SchedulerServer_2 (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_axi_mgmt_ar_ready,
	io_axi_mgmt_ar_valid,
	io_axi_mgmt_ar_bits_addr,
	io_axi_mgmt_ar_bits_prot,
	io_axi_mgmt_r_ready,
	io_axi_mgmt_r_valid,
	io_axi_mgmt_r_bits_data,
	io_axi_mgmt_r_bits_resp,
	io_axi_mgmt_aw_ready,
	io_axi_mgmt_aw_valid,
	io_axi_mgmt_aw_bits_addr,
	io_axi_mgmt_aw_bits_prot,
	io_axi_mgmt_w_ready,
	io_axi_mgmt_w_valid,
	io_axi_mgmt_w_bits_data,
	io_axi_mgmt_w_bits_strb,
	io_axi_mgmt_b_ready,
	io_axi_mgmt_b_valid,
	io_axi_mgmt_b_bits_resp,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_read_burst_len,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_write_burst_len,
	io_write_last,
	io_ntwDataUnitOccupancy
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [255:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [255:0] io_connNetwork_data_qOutTask_bits;
	output wire io_axi_mgmt_ar_ready;
	input io_axi_mgmt_ar_valid;
	input [5:0] io_axi_mgmt_ar_bits_addr;
	input [2:0] io_axi_mgmt_ar_bits_prot;
	input io_axi_mgmt_r_ready;
	output wire io_axi_mgmt_r_valid;
	output wire [63:0] io_axi_mgmt_r_bits_data;
	output wire [1:0] io_axi_mgmt_r_bits_resp;
	output wire io_axi_mgmt_aw_ready;
	input io_axi_mgmt_aw_valid;
	input [5:0] io_axi_mgmt_aw_bits_addr;
	input [2:0] io_axi_mgmt_aw_bits_prot;
	output wire io_axi_mgmt_w_ready;
	input io_axi_mgmt_w_valid;
	input [63:0] io_axi_mgmt_w_bits_data;
	input [7:0] io_axi_mgmt_w_bits_strb;
	input io_axi_mgmt_b_ready;
	output wire io_axi_mgmt_b_valid;
	output wire [1:0] io_axi_mgmt_b_bits_resp;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [255:0] io_read_data_bits;
	output wire [3:0] io_read_burst_len;
	input io_write_address_ready;
	output wire io_write_address_valid;
	output wire [63:0] io_write_address_bits;
	input io_write_data_ready;
	output wire io_write_data_valid;
	output wire [255:0] io_write_data_bits;
	output wire [3:0] io_write_burst_len;
	output wire io_write_last;
	input io_ntwDataUnitOccupancy;
	wire _taskQueueBuffer_io_enq_ready;
	wire [255:0] _taskQueueBuffer_io_deq_bits;
	wire [4:0] _taskQueueBuffer_io_count;
	wire _wrRespQueue__io_enq_ready;
	wire _wrRespQueue__io_deq_valid;
	wire _wrReqData__deq_q_io_enq_ready;
	wire _wrReqData__deq_q_io_deq_valid;
	wire [63:0] _wrReqData__deq_q_io_deq_bits_data;
	wire [7:0] _wrReqData__deq_q_io_deq_bits_strb;
	wire _wrReq__deq_q_io_enq_ready;
	wire _wrReq__deq_q_io_deq_valid;
	wire [5:0] _wrReq__deq_q_io_deq_bits_addr;
	wire _rdRespQueue__io_enq_ready;
	wire _rdRespQueue__io_deq_valid;
	wire [63:0] _rdRespQueue__io_deq_bits_data;
	wire [1:0] _rdRespQueue__io_deq_bits_resp;
	wire _rdReq__deq_q_io_enq_ready;
	wire _rdReq__deq_q_io_deq_valid;
	wire [5:0] _rdReq__deq_q_io_deq_bits_addr;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	wire rdReq = _rdReq__deq_q_io_deq_valid & _rdRespQueue__io_enq_ready;
	wire wrReq = (_wrReq__deq_q_io_deq_valid & _wrReqData__deq_q_io_deq_valid) & _wrRespQueue__io_enq_ready;
	reg [63:0] rAddr;
	reg [63:0] rPause;
	reg [63:0] procInterrupt;
	reg [63:0] maxLength;
	reg [3:0] stateReg;
	reg [63:0] currLen;
	reg [63:0] contentionCounter;
	reg networkCongested;
	reg [63:0] fifoTailReg;
	reg [63:0] fifoHeadReg;
	reg [4:0] memDataCounter;
	wire _GEN = stateReg == 4'h2;
	wire _GEN_0 = stateReg == 4'h4;
	wire _GEN_1 = stateReg == 4'h3;
	wire _GEN_2 = memDataCounter == 5'h01;
	wire _GEN_3 = _GEN | _GEN_0;
	wire _GEN_4 = stateReg == 4'h6;
	wire _GEN_5 = stateReg == 4'h5;
	wire _GEN_6 = (_GEN_0 | _GEN_1) | _GEN_4;
	wire _GEN_7 = _GEN | _GEN_6;
	wire _GEN_8 = stateReg == 4'h7;
	wire _GEN_9 = (_GEN | _GEN_0) | _GEN_1;
	wire _GEN_10 = _GEN_9 | ~_GEN_4;
	wire _GEN_11 = _GEN_4 | _GEN_5;
	wire [511:0] _GEN_12 = {64'hffffffffffffffff, currLen, procInterrupt, fifoHeadReg, fifoTailReg, maxLength, rAddr, rPause};
	always @(posedge clock)
		if (reset) begin
			rAddr <= 64'h0000000000000000;
			rPause <= 64'h0000000000000000;
			procInterrupt <= 64'h0000000000000000;
			maxLength <= 64'h0000000000000000;
			stateReg <= 4'h0;
			currLen <= 64'h0000000000000000;
			contentionCounter <= 64'h0000000000000000;
			networkCongested <= 1'h0;
			fifoTailReg <= 64'h0000000000000000;
			fifoHeadReg <= 64'h0000000000000000;
			memDataCounter <= 5'h00;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_13;
			reg _GEN_14;
			reg _GEN_15;
			reg [63:0] _GEN_16;
			reg _GEN_17;
			reg _GEN_18;
			reg _GEN_19;
			reg [63:0] _GEN_20;
			_GEN_19 = rPause == 64'h0000000000000000;
			_GEN_13 = stateReg == 4'h0;
			_GEN_14 = ((currLen == maxLength) & networkCongested) | (maxLength < (currLen + 64'h0000000000000010));
			_GEN_15 = io_write_data_ready & _GEN_2;
			_GEN_16 = maxLength - 64'h0000000000000001;
			_GEN_17 = _GEN_13 | _GEN_3;
			_GEN_18 = io_read_data_valid & _GEN_2;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h1))
				rAddr <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rAddr[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rAddr[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rAddr[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rAddr[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rAddr[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rAddr[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rAddr[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rAddr[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h0))
				rPause <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rPause[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rPause[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rPause[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rPause[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rPause[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rPause[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rPause[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rPause[7:0])};
			else if (_GEN_13 & (|procInterrupt | _GEN_14))
				rPause <= 64'hffffffffffffffff;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h5))
				procInterrupt <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : procInterrupt[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : procInterrupt[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : procInterrupt[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : procInterrupt[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : procInterrupt[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : procInterrupt[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : procInterrupt[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : procInterrupt[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h2))
				maxLength <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : maxLength[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : maxLength[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : maxLength[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : maxLength[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : maxLength[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : maxLength[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : maxLength[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : maxLength[7:0])};
			_GEN_20 = {stateReg, stateReg, stateReg, stateReg, stateReg, (_GEN_19 ? 4'h0 : 4'ha), (_GEN_19 ? 4'h0 : 4'h9), (io_connNetwork_ctrl_serveStealReq_ready ? 4'h7 : (networkCongested | (|procInterrupt) ? 4'h0 : stateReg)), (io_connNetwork_data_qOutTask_ready | networkCongested ? 4'h0 : 4'h7), (io_read_address_ready ? 4'h5 : stateReg), (_GEN_18 ? 4'h8 : stateReg), (io_write_address_ready ? 4'h3 : stateReg), (_GEN_15 ? 4'h0 : stateReg), ((_taskQueueBuffer_io_count == 5'h0f) & io_connNetwork_data_availableTask_valid ? 4'h4 : (io_connNetwork_data_availableTask_valid & networkCongested ? 4'h2 : (networkCongested ? stateReg : 4'h0))), stateReg, (|procInterrupt ? 4'ha : (_GEN_14 ? 4'h9 : (networkCongested & (_taskQueueBuffer_io_count == 5'h10) ? 4'h4 : (networkCongested ? 4'h2 : ((~networkCongested & |currLen) & ~(|_taskQueueBuffer_io_count) ? 4'h6 : (~networkCongested & |_taskQueueBuffer_io_count ? 4'h7 : stateReg))))))};
			stateReg <= _GEN_20[stateReg * 4+:4];
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h6))
				currLen <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : currLen[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : currLen[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : currLen[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : currLen[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : currLen[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : currLen[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : currLen[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : currLen[7:0])};
			else if (~_GEN_17) begin
				if (_GEN_1) begin
					if (_GEN_15)
						currLen <= currLen + 64'h0000000000000001;
					else if (io_write_data_ready)
						currLen <= currLen + 64'h0000000000000001;
				end
				else if (_GEN_4 | ~_GEN_5)
					;
				else if (_GEN_18)
					currLen <= currLen - 64'h0000000000000001;
				else if (io_read_data_valid)
					currLen <= currLen - 64'h0000000000000001;
			end
			if (io_ntwDataUnitOccupancy & (contentionCounter != 64'h0000000000000050))
				contentionCounter <= contentionCounter + 64'h0000000000000001;
			else if (|contentionCounter & ~io_ntwDataUnitOccupancy)
				contentionCounter <= contentionCounter - 64'h0000000000000001;
			networkCongested <= (contentionCounter > 64'h0000000000000042) | ((contentionCounter > 64'h0000000000000040) & networkCongested);
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h3))
				fifoTailReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoTailReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoTailReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoTailReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoTailReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoTailReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoTailReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoTailReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoTailReg[7:0])};
			else if (_GEN_17 | ~_GEN_1)
				;
			else begin : sv2v_autoblock_2
				reg _GEN_21;
				_GEN_21 = fifoTailReg < _GEN_16;
				if (_GEN_15) begin
					if (_GEN_21)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
				else if (io_write_data_ready) begin
					if (_GEN_21)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
			end
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h4))
				fifoHeadReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoHeadReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoHeadReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoHeadReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoHeadReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoHeadReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoHeadReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoHeadReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoHeadReg[7:0])};
			else if ((_GEN_13 | _GEN_7) | ~_GEN_5)
				;
			else begin : sv2v_autoblock_3
				reg _GEN_22;
				_GEN_22 = fifoHeadReg < _GEN_16;
				if (_GEN_18) begin
					if (_GEN_22)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
				else if (io_read_data_valid) begin
					if (_GEN_22)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
			end
			if (~(_GEN_13 | _GEN)) begin
				if (_GEN_0) begin
					if (io_write_address_ready)
						memDataCounter <= 5'h10;
				end
				else if (_GEN_1) begin
					if (_GEN_15 | ~io_write_data_ready)
						;
					else
						memDataCounter <= memDataCounter - 5'h01;
				end
				else if (_GEN_4) begin
					if (io_read_address_ready)
						memDataCounter <= (currLen < 64'h0000000000000010 ? currLen[4:0] : 5'h10);
				end
				else if ((~_GEN_5 | _GEN_18) | ~io_read_data_valid)
					;
				else
					memDataCounter <= memDataCounter - 5'h01;
			end
		end
	Queue2_AddressChannel_2 s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_ar_ready),
		.io_enq_valid(io_axi_mgmt_ar_valid),
		.io_enq_bits_addr(io_axi_mgmt_ar_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_ar_bits_prot),
		.io_deq_ready(_rdReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_rdRespQueue__io_deq_valid),
		.io_enq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_enq_bits_resp(_rdRespQueue__io_deq_bits_resp),
		.io_deq_ready(io_axi_mgmt_r_ready),
		.io_deq_valid(io_axi_mgmt_r_valid),
		.io_deq_bits_data(io_axi_mgmt_r_bits_data),
		.io_deq_bits_resp(io_axi_mgmt_r_bits_resp)
	);
	Queue2_AddressChannel_2 s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_aw_ready),
		.io_enq_valid(io_axi_mgmt_aw_valid),
		.io_enq_bits_addr(io_axi_mgmt_aw_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_aw_bits_prot),
		.io_deq_ready(_wrReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_w_ready),
		.io_enq_valid(io_axi_mgmt_w_valid),
		.io_enq_bits_data(io_axi_mgmt_w_bits_data),
		.io_enq_bits_strb(io_axi_mgmt_w_bits_strb),
		.io_deq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_wrRespQueue__io_deq_valid),
		.io_enq_bits_resp(2'h0),
		.io_deq_ready(io_axi_mgmt_b_ready),
		.io_deq_valid(io_axi_mgmt_b_valid),
		.io_deq_bits_resp(io_axi_mgmt_b_bits_resp)
	);
	Queue1_AddressChannel rdReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_deq_ready(rdReq),
		.io_deq_valid(_rdReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_rdReq__deq_q_io_deq_bits_addr)
	);
	Queue1_ReadDataChannel rdRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdRespQueue__io_enq_ready),
		.io_enq_valid(rdReq),
		.io_enq_bits_data(_GEN_12[_rdReq__deq_q_io_deq_bits_addr[5:3] * 64+:64]),
		.io_deq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_deq_valid(_rdRespQueue__io_deq_valid),
		.io_deq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_deq_bits_resp(_rdRespQueue__io_deq_bits_resp)
	);
	Queue1_AddressChannel wrReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_wrReq__deq_q_io_deq_bits_addr)
	);
	Queue1_WriteDataChannel wrReqData__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_enq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_enq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReqData__deq_q_io_deq_valid),
		.io_deq_bits_data(_wrReqData__deq_q_io_deq_bits_data),
		.io_deq_bits_strb(_wrReqData__deq_q_io_deq_bits_strb)
	);
	Queue1_WriteResponseChannel wrRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrRespQueue__io_enq_ready),
		.io_enq_valid(wrReq),
		.io_deq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_deq_valid(_wrRespQueue__io_deq_valid)
	);
	Queue16_UInt_2 taskQueueBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_taskQueueBuffer_io_enq_ready),
		.io_enq_valid((_GEN ? io_connNetwork_data_availableTask_valid : (~_GEN_6 & _GEN_5) & io_read_data_valid)),
		.io_enq_bits((_GEN ? io_connNetwork_data_availableTask_bits : (_GEN_6 | ~_GEN_5 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : io_read_data_bits))),
		.io_deq_ready(~_GEN_3 & (_GEN_1 ? io_write_data_ready : (~_GEN_11 & _GEN_8) & io_connNetwork_data_qOutTask_ready)),
		.io_deq_valid(),
		.io_deq_bits(_taskQueueBuffer_io_deq_bits),
		.io_count(_taskQueueBuffer_io_count)
	);
	assign io_connNetwork_ctrl_serveStealReq_valid = ~(((((_GEN | _GEN_0) | _GEN_1) | _GEN_4) | _GEN_5) | _GEN_8) & (stateReg == 4'h8);
	assign io_connNetwork_data_availableTask_ready = _GEN & _taskQueueBuffer_io_enq_ready;
	assign io_connNetwork_data_qOutTask_valid = ~(((_GEN | _GEN_0) | _GEN_1) | _GEN_11) & _GEN_8;
	assign io_connNetwork_data_qOutTask_bits = _taskQueueBuffer_io_deq_bits;
	assign io_read_address_valid = ~_GEN_9 & _GEN_4;
	assign io_read_address_bits = (_GEN_10 ? 64'h0000000000000000 : {fifoHeadReg[58:0], 5'h00} + rAddr);
	assign io_read_data_ready = ~_GEN_7 & _GEN_5;
	assign io_read_burst_len = (_GEN_10 ? 4'h0 : (currLen < 64'h0000000000000010 ? currLen[3:0] - 4'h1 : 4'hf));
	assign io_write_address_valid = ~_GEN & _GEN_0;
	assign io_write_address_bits = (_GEN | ~_GEN_0 ? 64'h0000000000000000 : {fifoTailReg[58:0], 5'h00} + rAddr);
	assign io_write_data_valid = ~_GEN_3 & _GEN_1;
	assign io_write_data_bits = _taskQueueBuffer_io_deq_bits;
	assign io_write_burst_len = (_GEN ? 4'h0 : {4 {_GEN_0}});
	assign io_write_last = (~_GEN_3 & _GEN_1) & _GEN_2;
endmodule
module RVtoAXIBridge_2 (
	clock,
	reset,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_writeBurst_len,
	io_writeBurst_last,
	io_readBurst_len,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_ar_bits_len,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data,
	axi_aw_ready,
	axi_aw_valid,
	axi_aw_bits_addr,
	axi_aw_bits_len,
	axi_w_ready,
	axi_w_valid,
	axi_w_bits_data,
	axi_w_bits_last,
	axi_b_valid
);
	input clock;
	input reset;
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [255:0] io_read_data_bits;
	output wire io_write_address_ready;
	input io_write_address_valid;
	input [63:0] io_write_address_bits;
	output wire io_write_data_ready;
	input io_write_data_valid;
	input [255:0] io_write_data_bits;
	input [3:0] io_writeBurst_len;
	input io_writeBurst_last;
	input [3:0] io_readBurst_len;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire [7:0] axi_ar_bits_len;
	output wire axi_r_ready;
	input axi_r_valid;
	input [255:0] axi_r_bits_data;
	input axi_aw_ready;
	output wire axi_aw_valid;
	output wire [63:0] axi_aw_bits_addr;
	output wire [7:0] axi_aw_bits_len;
	input axi_w_ready;
	output wire axi_w_valid;
	output wire [255:0] axi_w_bits_data;
	output wire axi_w_bits_last;
	input axi_b_valid;
	reg writeHandshakeDetector;
	wire axi_w_valid_0 = (io_write_data_valid & axi_w_ready) & ~writeHandshakeDetector;
	always @(posedge clock)
		if (reset)
			writeHandshakeDetector <= 1'h0;
		else if (axi_w_valid_0)
			writeHandshakeDetector <= io_writeBurst_last | writeHandshakeDetector;
		else
			writeHandshakeDetector <= ~axi_b_valid & writeHandshakeDetector;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign io_write_address_ready = axi_aw_ready;
	assign io_write_data_ready = axi_w_ready & ~writeHandshakeDetector;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_ar_bits_len = {4'h0, io_readBurst_len};
	assign axi_r_ready = io_read_data_ready;
	assign axi_aw_valid = io_write_address_valid;
	assign axi_aw_bits_addr = io_write_address_bits;
	assign axi_aw_bits_len = {4'h0, io_writeBurst_len};
	assign axi_w_valid = axi_w_valid_0;
	assign axi_w_bits_data = io_write_data_bits;
	assign axi_w_bits_last = io_writeBurst_last;
endmodule
module Queue1_ReadDataChannel_6 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits_id;
	input [255:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [255:0] io_deq_bits_data;
	reg [259:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_last, io_enq_bits_resp, io_enq_bits_data, io_enq_bits_id};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[256:1];
endmodule
module Queue1_WriteDataChannel_6 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [255:0] io_enq_bits_data;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [255:0] io_deq_bits_data;
	output wire [31:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	reg [288:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_last, 32'hffffffff, io_enq_bits_data};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[255:0];
	assign io_deq_bits_strb = ram[287:256];
	assign io_deq_bits_last = ram[288];
endmodule
module ram_2x261 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [260:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [260:0] W0_data;
	reg [260:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 261'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel_6 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_data,
	io_deq_bits_resp,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_id;
	input [255:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_id;
	output wire [255:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	output wire io_deq_bits_last;
	wire [260:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x261 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_resp, io_enq_bits_data, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[1:0];
	assign io_deq_bits_data = _ram_ext_R0_data[257:2];
	assign io_deq_bits_resp = _ram_ext_R0_data[259:258];
	assign io_deq_bits_last = _ram_ext_R0_data[260];
endmodule
module ram_2x289 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [288:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [288:0] W0_data;
	reg [288:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteDataChannel_6 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [255:0] io_enq_bits_data;
	input [31:0] io_enq_bits_strb;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [255:0] io_deq_bits_data;
	output wire [31:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	wire [288:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x289 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_strb, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[255:0];
	assign io_deq_bits_strb = _ram_ext_R0_data[287:256];
	assign io_deq_bits_last = _ram_ext_R0_data[288];
endmodule
module elasticDemux_5 (
	io_source_ready,
	io_source_valid,
	io_source_bits_id,
	io_source_bits_data,
	io_source_bits_resp,
	io_source_bits_last,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_id,
	io_sinks_0_bits_data,
	io_sinks_0_bits_resp,
	io_sinks_0_bits_last,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_id,
	io_sinks_1_bits_data,
	io_sinks_1_bits_resp,
	io_sinks_1_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [1:0] io_source_bits_id;
	input [255:0] io_source_bits_data;
	input [1:0] io_source_bits_resp;
	input io_source_bits_last;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [1:0] io_sinks_0_bits_id;
	output wire [255:0] io_sinks_0_bits_data;
	output wire [1:0] io_sinks_0_bits_resp;
	output wire io_sinks_0_bits_last;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [1:0] io_sinks_1_bits_id;
	output wire [255:0] io_sinks_1_bits_data;
	output wire [1:0] io_sinks_1_bits_resp;
	output wire io_sinks_1_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire fire = valid & (io_select_bits ? io_sinks_1_ready : io_sinks_0_ready);
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & ~io_select_bits;
	assign io_sinks_0_bits_id = io_source_bits_id;
	assign io_sinks_0_bits_data = io_source_bits_data;
	assign io_sinks_0_bits_resp = io_source_bits_resp;
	assign io_sinks_0_bits_last = io_source_bits_last;
	assign io_sinks_1_valid = valid & io_select_bits;
	assign io_sinks_1_bits_id = io_source_bits_id;
	assign io_sinks_1_bits_data = io_source_bits_data;
	assign io_sinks_1_bits_resp = io_source_bits_resp;
	assign io_sinks_1_bits_last = io_source_bits_last;
	assign io_select_ready = fire;
endmodule
module elasticMux_3 (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_data,
	io_sources_0_bits_strb,
	io_sources_0_bits_last,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_data,
	io_sources_1_bits_strb,
	io_sources_1_bits_last,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_data,
	io_sink_bits_strb,
	io_sink_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [255:0] io_sources_0_bits_data;
	input [31:0] io_sources_0_bits_strb;
	input io_sources_0_bits_last;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [255:0] io_sources_1_bits_data;
	input [31:0] io_sources_1_bits_strb;
	input io_sources_1_bits_last;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [255:0] io_sink_bits_data;
	output wire [31:0] io_sink_bits_strb;
	output wire io_sink_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input io_select_bits;
	wire io_sink_bits_last_0 = (io_select_bits ? io_sources_1_bits_last : io_sources_0_bits_last);
	wire valid = io_select_valid & (io_select_bits ? io_sources_1_valid : io_sources_0_valid);
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & ~io_select_bits;
	assign io_sources_1_ready = fire & io_select_bits;
	assign io_sink_valid = valid;
	assign io_sink_bits_data = (io_select_bits ? io_sources_1_bits_data : io_sources_0_bits_data);
	assign io_sink_bits_strb = (io_select_bits ? io_sources_1_bits_strb : io_sources_0_bits_strb);
	assign io_sink_bits_last = io_sink_bits_last_0;
	assign io_select_ready = fire & io_sink_bits_last_0;
endmodule
module axi4FullMux_1 (
	clock,
	reset,
	s_axi_0_ar_ready,
	s_axi_0_ar_valid,
	s_axi_0_ar_bits_addr,
	s_axi_0_ar_bits_len,
	s_axi_0_ar_bits_size,
	s_axi_0_ar_bits_burst,
	s_axi_0_ar_bits_lock,
	s_axi_0_ar_bits_cache,
	s_axi_0_ar_bits_prot,
	s_axi_0_ar_bits_qos,
	s_axi_0_ar_bits_region,
	s_axi_0_r_ready,
	s_axi_0_r_valid,
	s_axi_0_r_bits_data,
	s_axi_0_aw_ready,
	s_axi_0_aw_valid,
	s_axi_0_aw_bits_addr,
	s_axi_0_aw_bits_len,
	s_axi_0_aw_bits_size,
	s_axi_0_aw_bits_burst,
	s_axi_0_aw_bits_lock,
	s_axi_0_aw_bits_cache,
	s_axi_0_aw_bits_prot,
	s_axi_0_aw_bits_qos,
	s_axi_0_aw_bits_region,
	s_axi_0_w_ready,
	s_axi_0_w_valid,
	s_axi_0_w_bits_data,
	s_axi_0_w_bits_last,
	s_axi_0_b_valid,
	s_axi_1_ar_ready,
	s_axi_1_ar_valid,
	s_axi_1_ar_bits_addr,
	s_axi_1_ar_bits_len,
	s_axi_1_ar_bits_size,
	s_axi_1_ar_bits_burst,
	s_axi_1_ar_bits_lock,
	s_axi_1_ar_bits_cache,
	s_axi_1_ar_bits_prot,
	s_axi_1_ar_bits_qos,
	s_axi_1_ar_bits_region,
	s_axi_1_r_ready,
	s_axi_1_r_valid,
	s_axi_1_r_bits_data,
	s_axi_1_aw_ready,
	s_axi_1_aw_valid,
	s_axi_1_aw_bits_addr,
	s_axi_1_aw_bits_len,
	s_axi_1_aw_bits_size,
	s_axi_1_aw_bits_burst,
	s_axi_1_aw_bits_lock,
	s_axi_1_aw_bits_cache,
	s_axi_1_aw_bits_prot,
	s_axi_1_aw_bits_qos,
	s_axi_1_aw_bits_region,
	s_axi_1_w_ready,
	s_axi_1_w_valid,
	s_axi_1_w_bits_data,
	s_axi_1_w_bits_last,
	s_axi_1_b_valid,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_id,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_id,
	m_axi_r_bits_data,
	m_axi_r_bits_resp,
	m_axi_r_bits_last,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_id,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_strb,
	m_axi_w_bits_last,
	m_axi_b_ready,
	m_axi_b_valid,
	m_axi_b_bits_id,
	m_axi_b_bits_resp
);
	input clock;
	input reset;
	output wire s_axi_0_ar_ready;
	input s_axi_0_ar_valid;
	input [63:0] s_axi_0_ar_bits_addr;
	input [7:0] s_axi_0_ar_bits_len;
	input [2:0] s_axi_0_ar_bits_size;
	input [1:0] s_axi_0_ar_bits_burst;
	input s_axi_0_ar_bits_lock;
	input [3:0] s_axi_0_ar_bits_cache;
	input [2:0] s_axi_0_ar_bits_prot;
	input [3:0] s_axi_0_ar_bits_qos;
	input [3:0] s_axi_0_ar_bits_region;
	input s_axi_0_r_ready;
	output wire s_axi_0_r_valid;
	output wire [255:0] s_axi_0_r_bits_data;
	output wire s_axi_0_aw_ready;
	input s_axi_0_aw_valid;
	input [63:0] s_axi_0_aw_bits_addr;
	input [7:0] s_axi_0_aw_bits_len;
	input [2:0] s_axi_0_aw_bits_size;
	input [1:0] s_axi_0_aw_bits_burst;
	input s_axi_0_aw_bits_lock;
	input [3:0] s_axi_0_aw_bits_cache;
	input [2:0] s_axi_0_aw_bits_prot;
	input [3:0] s_axi_0_aw_bits_qos;
	input [3:0] s_axi_0_aw_bits_region;
	output wire s_axi_0_w_ready;
	input s_axi_0_w_valid;
	input [255:0] s_axi_0_w_bits_data;
	input s_axi_0_w_bits_last;
	output wire s_axi_0_b_valid;
	output wire s_axi_1_ar_ready;
	input s_axi_1_ar_valid;
	input [63:0] s_axi_1_ar_bits_addr;
	input [7:0] s_axi_1_ar_bits_len;
	input [2:0] s_axi_1_ar_bits_size;
	input [1:0] s_axi_1_ar_bits_burst;
	input s_axi_1_ar_bits_lock;
	input [3:0] s_axi_1_ar_bits_cache;
	input [2:0] s_axi_1_ar_bits_prot;
	input [3:0] s_axi_1_ar_bits_qos;
	input [3:0] s_axi_1_ar_bits_region;
	input s_axi_1_r_ready;
	output wire s_axi_1_r_valid;
	output wire [255:0] s_axi_1_r_bits_data;
	output wire s_axi_1_aw_ready;
	input s_axi_1_aw_valid;
	input [63:0] s_axi_1_aw_bits_addr;
	input [7:0] s_axi_1_aw_bits_len;
	input [2:0] s_axi_1_aw_bits_size;
	input [1:0] s_axi_1_aw_bits_burst;
	input s_axi_1_aw_bits_lock;
	input [3:0] s_axi_1_aw_bits_cache;
	input [2:0] s_axi_1_aw_bits_prot;
	input [3:0] s_axi_1_aw_bits_qos;
	input [3:0] s_axi_1_aw_bits_region;
	output wire s_axi_1_w_ready;
	input s_axi_1_w_valid;
	input [255:0] s_axi_1_w_bits_data;
	input s_axi_1_w_bits_last;
	output wire s_axi_1_b_valid;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [1:0] m_axi_ar_bits_id;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [1:0] m_axi_r_bits_id;
	input [255:0] m_axi_r_bits_data;
	input [1:0] m_axi_r_bits_resp;
	input m_axi_r_bits_last;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [1:0] m_axi_aw_bits_id;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [255:0] m_axi_w_bits_data;
	output wire [31:0] m_axi_w_bits_strb;
	output wire m_axi_w_bits_last;
	output wire m_axi_b_ready;
	input m_axi_b_valid;
	input [1:0] m_axi_b_bits_id;
	input [1:0] m_axi_b_bits_resp;
	wire _write_demux_io_source_ready;
	wire _write_demux_io_sinks_0_valid;
	wire _write_demux_io_sinks_1_valid;
	wire _write_demux_io_select_ready;
	wire _write_mux_io_sources_0_ready;
	wire _write_mux_io_sources_1_ready;
	wire _write_mux_io_sink_valid;
	wire [255:0] _write_mux_io_sink_bits_data;
	wire [31:0] _write_mux_io_sink_bits_strb;
	wire _write_mux_io_sink_bits_last;
	wire _write_mux_io_select_ready;
	wire _write_arbiter_io_sources_0_ready;
	wire _write_arbiter_io_sources_1_ready;
	wire _write_arbiter_io_sink_valid;
	wire [1:0] _write_arbiter_io_sink_bits_id;
	wire [63:0] _write_arbiter_io_sink_bits_addr;
	wire [7:0] _write_arbiter_io_sink_bits_len;
	wire [2:0] _write_arbiter_io_sink_bits_size;
	wire [1:0] _write_arbiter_io_sink_bits_burst;
	wire _write_arbiter_io_sink_bits_lock;
	wire [3:0] _write_arbiter_io_sink_bits_cache;
	wire [2:0] _write_arbiter_io_sink_bits_prot;
	wire [3:0] _write_arbiter_io_sink_bits_qos;
	wire [3:0] _write_arbiter_io_sink_bits_region;
	wire _write_arbiter_io_select_valid;
	wire _write_arbiter_io_select_bits;
	wire _write_portQueue_io_enq_ready;
	wire _write_portQueue_io_deq_valid;
	wire _write_portQueue_io_deq_bits;
	wire _read_demux_io_source_ready;
	wire _read_demux_io_sinks_0_valid;
	wire [1:0] _read_demux_io_sinks_0_bits_id;
	wire [255:0] _read_demux_io_sinks_0_bits_data;
	wire [1:0] _read_demux_io_sinks_0_bits_resp;
	wire _read_demux_io_sinks_0_bits_last;
	wire _read_demux_io_sinks_1_valid;
	wire [1:0] _read_demux_io_sinks_1_bits_id;
	wire [255:0] _read_demux_io_sinks_1_bits_data;
	wire [1:0] _read_demux_io_sinks_1_bits_resp;
	wire _read_demux_io_sinks_1_bits_last;
	wire _read_demux_io_select_ready;
	wire _read_arbiter_io_sources_0_ready;
	wire _read_arbiter_io_sources_1_ready;
	wire _read_arbiter_io_sink_valid;
	wire [1:0] _read_arbiter_io_sink_bits_id;
	wire [63:0] _read_arbiter_io_sink_bits_addr;
	wire [7:0] _read_arbiter_io_sink_bits_len;
	wire [2:0] _read_arbiter_io_sink_bits_size;
	wire [1:0] _read_arbiter_io_sink_bits_burst;
	wire _read_arbiter_io_sink_bits_lock;
	wire [3:0] _read_arbiter_io_sink_bits_cache;
	wire [2:0] _read_arbiter_io_sink_bits_prot;
	wire [3:0] _read_arbiter_io_sink_bits_qos;
	wire [3:0] _read_arbiter_io_sink_bits_region;
	wire _m_axi__sinkBuffer_1_io_deq_valid;
	wire [1:0] _m_axi__sinkBuffer_1_io_deq_bits_id;
	wire _m_axi__sourceBuffer_2_io_enq_ready;
	wire _m_axi__sourceBuffer_1_io_enq_ready;
	wire _m_axi__sinkBuffer_io_deq_valid;
	wire [1:0] _m_axi__sinkBuffer_io_deq_bits_id;
	wire [255:0] _m_axi__sinkBuffer_io_deq_bits_data;
	wire [1:0] _m_axi__sinkBuffer_io_deq_bits_resp;
	wire _m_axi__sinkBuffer_io_deq_bits_last;
	wire _m_axi__sourceBuffer_io_enq_ready;
	wire _s_axi__buffered_sinkBuffer_3_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_valid;
	wire [255:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_data;
	wire [31:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_2_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_1_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_valid;
	wire [255:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_data;
	wire [31:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_region;
	reg read_eagerFork_regs_0;
	reg read_eagerFork_regs_1;
	wire read_eagerFork_m_axi__r_ready_qual1_0 = _read_demux_io_source_ready | read_eagerFork_regs_0;
	wire read_eagerFork_m_axi__r_ready_qual1_1 = _read_demux_io_select_ready | read_eagerFork_regs_1;
	wire m_axi__r_ready = read_eagerFork_m_axi__r_ready_qual1_0 & read_eagerFork_m_axi__r_ready_qual1_1;
	reg write_eagerFork_regs_0;
	reg write_eagerFork_regs_1;
	wire write_eagerFork_m_axi__b_ready_qual1_0 = _write_demux_io_source_ready | write_eagerFork_regs_0;
	wire write_eagerFork_m_axi__b_ready_qual1_1 = _write_demux_io_select_ready | write_eagerFork_regs_1;
	wire m_axi__b_ready = write_eagerFork_m_axi__b_ready_qual1_0 & write_eagerFork_m_axi__b_ready_qual1_1;
	always @(posedge clock)
		if (reset) begin
			read_eagerFork_regs_0 <= 1'h0;
			read_eagerFork_regs_1 <= 1'h0;
			write_eagerFork_regs_0 <= 1'h0;
			write_eagerFork_regs_1 <= 1'h0;
		end
		else begin
			read_eagerFork_regs_0 <= (read_eagerFork_m_axi__r_ready_qual1_0 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			read_eagerFork_regs_1 <= (read_eagerFork_m_axi__r_ready_qual1_1 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			write_eagerFork_regs_0 <= (write_eagerFork_m_axi__b_ready_qual1_0 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
			write_eagerFork_regs_1 <= (write_eagerFork_m_axi__b_ready_qual1_1 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
		end
	Queue1_ReadAddressChannel s_axi__buffered_sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_ar_ready),
		.io_enq_valid(s_axi_0_ar_valid),
		.io_enq_bits_addr(s_axi_0_ar_bits_addr),
		.io_enq_bits_len(s_axi_0_ar_bits_len),
		.io_enq_bits_size(s_axi_0_ar_bits_size),
		.io_enq_bits_burst(s_axi_0_ar_bits_burst),
		.io_enq_bits_lock(s_axi_0_ar_bits_lock),
		.io_enq_bits_cache(s_axi_0_ar_bits_cache),
		.io_enq_bits_prot(s_axi_0_ar_bits_prot),
		.io_enq_bits_qos(s_axi_0_ar_bits_qos),
		.io_enq_bits_region(s_axi_0_ar_bits_region),
		.io_deq_ready(_read_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region)
	);
	Queue1_ReadDataChannel_6 s_axi__buffered_sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_0_valid),
		.io_enq_bits_id(_read_demux_io_sinks_0_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_deq_ready(s_axi_0_r_ready),
		.io_deq_valid(s_axi_0_r_valid),
		.io_deq_bits_data(s_axi_0_r_bits_data)
	);
	Queue1_WriteAddressChannel s_axi__buffered_sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_aw_ready),
		.io_enq_valid(s_axi_0_aw_valid),
		.io_enq_bits_addr(s_axi_0_aw_bits_addr),
		.io_enq_bits_len(s_axi_0_aw_bits_len),
		.io_enq_bits_size(s_axi_0_aw_bits_size),
		.io_enq_bits_burst(s_axi_0_aw_bits_burst),
		.io_enq_bits_lock(s_axi_0_aw_bits_lock),
		.io_enq_bits_cache(s_axi_0_aw_bits_cache),
		.io_enq_bits_prot(s_axi_0_aw_bits_prot),
		.io_enq_bits_qos(s_axi_0_aw_bits_qos),
		.io_enq_bits_region(s_axi_0_aw_bits_region),
		.io_deq_ready(_write_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_1_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region)
	);
	Queue1_WriteDataChannel_6 s_axi__buffered_sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_w_ready),
		.io_enq_valid(s_axi_0_w_valid),
		.io_enq_bits_data(s_axi_0_w_bits_data),
		.io_enq_bits_last(s_axi_0_w_bits_last),
		.io_deq_ready(_write_mux_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last)
	);
	Queue1_WriteResponseChannel_2 s_axi__buffered_sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_0_valid),
		.io_deq_valid(s_axi_0_b_valid)
	);
	Queue1_ReadAddressChannel s_axi__buffered_sourceBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_ar_ready),
		.io_enq_valid(s_axi_1_ar_valid),
		.io_enq_bits_addr(s_axi_1_ar_bits_addr),
		.io_enq_bits_len(s_axi_1_ar_bits_len),
		.io_enq_bits_size(s_axi_1_ar_bits_size),
		.io_enq_bits_burst(s_axi_1_ar_bits_burst),
		.io_enq_bits_lock(s_axi_1_ar_bits_lock),
		.io_enq_bits_cache(s_axi_1_ar_bits_cache),
		.io_enq_bits_prot(s_axi_1_ar_bits_prot),
		.io_enq_bits_qos(s_axi_1_ar_bits_qos),
		.io_enq_bits_region(s_axi_1_ar_bits_region),
		.io_deq_ready(_read_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_3_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region)
	);
	Queue1_ReadDataChannel_6 s_axi__buffered_sinkBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_1_valid),
		.io_enq_bits_id(_read_demux_io_sinks_1_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_deq_ready(s_axi_1_r_ready),
		.io_deq_valid(s_axi_1_r_valid),
		.io_deq_bits_data(s_axi_1_r_bits_data)
	);
	Queue1_WriteAddressChannel s_axi__buffered_sourceBuffer_4(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_aw_ready),
		.io_enq_valid(s_axi_1_aw_valid),
		.io_enq_bits_addr(s_axi_1_aw_bits_addr),
		.io_enq_bits_len(s_axi_1_aw_bits_len),
		.io_enq_bits_size(s_axi_1_aw_bits_size),
		.io_enq_bits_burst(s_axi_1_aw_bits_burst),
		.io_enq_bits_lock(s_axi_1_aw_bits_lock),
		.io_enq_bits_cache(s_axi_1_aw_bits_cache),
		.io_enq_bits_prot(s_axi_1_aw_bits_prot),
		.io_enq_bits_qos(s_axi_1_aw_bits_qos),
		.io_enq_bits_region(s_axi_1_aw_bits_region),
		.io_deq_ready(_write_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_4_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region)
	);
	Queue1_WriteDataChannel_6 s_axi__buffered_sourceBuffer_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_w_ready),
		.io_enq_valid(s_axi_1_w_valid),
		.io_enq_bits_data(s_axi_1_w_bits_data),
		.io_enq_bits_last(s_axi_1_w_bits_last),
		.io_deq_ready(_write_mux_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last)
	);
	Queue1_WriteResponseChannel_2 s_axi__buffered_sinkBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_1_valid),
		.io_deq_valid(s_axi_1_b_valid)
	);
	Queue2_ReadAddressChannel m_axi__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_enq_valid(_read_arbiter_io_sink_valid),
		.io_enq_bits_id(_read_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_read_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_read_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_read_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_id(m_axi_ar_bits_id),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	Queue2_ReadDataChannel_6 m_axi__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_r_ready),
		.io_enq_valid(m_axi_r_valid),
		.io_enq_bits_id(m_axi_r_bits_id),
		.io_enq_bits_data(m_axi_r_bits_data),
		.io_enq_bits_resp(m_axi_r_bits_resp),
		.io_enq_bits_last(m_axi_r_bits_last),
		.io_deq_ready(m_axi__r_ready),
		.io_deq_valid(_m_axi__sinkBuffer_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_deq_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_deq_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_deq_bits_last(_m_axi__sinkBuffer_io_deq_bits_last)
	);
	Queue2_WriteAddressChannel m_axi__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_sink_valid),
		.io_enq_bits_id(_write_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_write_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_write_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_write_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_id(m_axi_aw_bits_id),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_WriteDataChannel_6 m_axi__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_enq_valid(_write_mux_io_sink_valid),
		.io_enq_bits_data(_write_mux_io_sink_bits_data),
		.io_enq_bits_strb(_write_mux_io_sink_bits_strb),
		.io_enq_bits_last(_write_mux_io_sink_bits_last),
		.io_deq_ready(m_axi_w_ready),
		.io_deq_valid(m_axi_w_valid),
		.io_deq_bits_data(m_axi_w_bits_data),
		.io_deq_bits_strb(m_axi_w_bits_strb),
		.io_deq_bits_last(m_axi_w_bits_last)
	);
	Queue2_WriteResponseChannel_3 m_axi__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_b_ready),
		.io_enq_valid(m_axi_b_valid),
		.io_enq_bits_id(m_axi_b_bits_id),
		.io_enq_bits_resp(m_axi_b_bits_resp),
		.io_deq_ready(m_axi__b_ready),
		.io_deq_valid(_m_axi__sinkBuffer_1_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_1_io_deq_bits_id)
	);
	elasticArbiter read_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_read_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_sources_0_bits_id({1'h0, _s_axi__buffered_sourceBuffer_io_deq_bits_id}),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region),
		.io_sources_1_ready(_read_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_sources_1_bits_id({1'h1, _s_axi__buffered_sourceBuffer_3_io_deq_bits_id}),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_sink_valid(_read_arbiter_io_sink_valid),
		.io_sink_bits_id(_read_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_read_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_read_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_read_arbiter_io_sink_bits_region),
		.io_select_ready(1'h1),
		.io_select_valid(),
		.io_select_bits()
	);
	elasticDemux_5 read_demux(
		.io_source_ready(_read_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_0),
		.io_source_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_source_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_source_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_source_bits_last(_m_axi__sinkBuffer_io_deq_bits_last),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_sinks_0_valid(_read_demux_io_sinks_0_valid),
		.io_sinks_0_bits_id(_read_demux_io_sinks_0_bits_id),
		.io_sinks_0_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_sinks_0_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_sinks_0_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_sinks_1_valid(_read_demux_io_sinks_1_valid),
		.io_sinks_1_bits_id(_read_demux_io_sinks_1_bits_id),
		.io_sinks_1_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_sinks_1_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_sinks_1_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_select_ready(_read_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_io_deq_bits_id[1])
	);
	Queue32_UInt1 write_portQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueue_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_select_valid),
		.io_enq_bits(_write_arbiter_io_select_bits),
		.io_deq_ready(_write_mux_io_select_ready),
		.io_deq_valid(_write_portQueue_io_deq_valid),
		.io_deq_bits(_write_portQueue_io_deq_bits)
	);
	elasticArbiter write_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_write_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_sources_0_bits_id({1'h0, _s_axi__buffered_sourceBuffer_1_io_deq_bits_id}),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region),
		.io_sources_1_ready(_write_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_sources_1_bits_id({1'h1, _s_axi__buffered_sourceBuffer_4_io_deq_bits_id}),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_sink_valid(_write_arbiter_io_sink_valid),
		.io_sink_bits_id(_write_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_write_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_write_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_write_arbiter_io_sink_bits_region),
		.io_select_ready(_write_portQueue_io_enq_ready),
		.io_select_valid(_write_arbiter_io_select_valid),
		.io_select_bits(_write_arbiter_io_select_bits)
	);
	elasticMux_3 write_mux(
		.io_sources_0_ready(_write_mux_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_sources_0_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_sources_0_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_sources_0_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last),
		.io_sources_1_ready(_write_mux_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_sources_1_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_sources_1_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_sources_1_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last),
		.io_sink_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_sink_valid(_write_mux_io_sink_valid),
		.io_sink_bits_data(_write_mux_io_sink_bits_data),
		.io_sink_bits_strb(_write_mux_io_sink_bits_strb),
		.io_sink_bits_last(_write_mux_io_sink_bits_last),
		.io_select_ready(_write_mux_io_select_ready),
		.io_select_valid(_write_portQueue_io_deq_valid),
		.io_select_bits(_write_portQueue_io_deq_bits)
	);
	elasticDemux_4 write_demux(
		.io_source_ready(_write_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_0),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_sinks_0_valid(_write_demux_io_sinks_0_valid),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_sinks_1_valid(_write_demux_io_sinks_1_valid),
		.io_select_ready(_write_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_1_io_deq_bits_id[1])
	);
endmodule
module AxiWriteBuffer_2 (
	clock,
	reset,
	s_axi_ar_ready,
	s_axi_ar_valid,
	s_axi_ar_bits_addr,
	s_axi_ar_bits_len,
	s_axi_r_ready,
	s_axi_r_valid,
	s_axi_r_bits_data,
	s_axi_aw_ready,
	s_axi_aw_valid,
	s_axi_aw_bits_addr,
	s_axi_aw_bits_len,
	s_axi_w_ready,
	s_axi_w_valid,
	s_axi_w_bits_data,
	s_axi_w_bits_last,
	s_axi_b_valid,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_data,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_last,
	m_axi_b_valid
);
	input clock;
	input reset;
	output wire s_axi_ar_ready;
	input s_axi_ar_valid;
	input [63:0] s_axi_ar_bits_addr;
	input [7:0] s_axi_ar_bits_len;
	input s_axi_r_ready;
	output wire s_axi_r_valid;
	output wire [255:0] s_axi_r_bits_data;
	output wire s_axi_aw_ready;
	input s_axi_aw_valid;
	input [63:0] s_axi_aw_bits_addr;
	input [7:0] s_axi_aw_bits_len;
	output wire s_axi_w_ready;
	input s_axi_w_valid;
	input [255:0] s_axi_w_bits_data;
	input s_axi_w_bits_last;
	output wire s_axi_b_valid;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [255:0] m_axi_r_bits_data;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [255:0] m_axi_w_bits_data;
	output wire m_axi_w_bits_last;
	input m_axi_b_valid;
	wire s_axi_aw_ready_0;
	wire _sinkBuffered__sinkBuffer_1_io_enq_ready;
	wire _sinkBuffered__sinkBuffer_io_enq_ready;
	wire _counter_io_empty;
	wire _counter_io_full;
	wire _counter_io_incEn_T = s_axi_aw_ready_0 & s_axi_aw_valid;
	assign s_axi_aw_ready_0 = (_sinkBuffered__sinkBuffer_io_enq_ready & s_axi_aw_valid) & ~_counter_io_full;
	wire s_axi_ar_ready_0 = ((_sinkBuffered__sinkBuffer_1_io_enq_ready & s_axi_ar_valid) & _counter_io_empty) & ~_counter_io_incEn_T;
	Counter counter(
		.clock(clock),
		.reset(reset),
		.io_incEn(_counter_io_incEn_T),
		.io_decEn(m_axi_b_valid),
		.io_empty(_counter_io_empty),
		.io_full(_counter_io_full)
	);
	Queue2_WriteAddressChannel_1 sinkBuffered__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_io_enq_ready),
		.io_enq_valid(s_axi_aw_ready_0),
		.io_enq_bits_addr(s_axi_aw_bits_addr),
		.io_enq_bits_len(s_axi_aw_bits_len),
		.io_enq_bits_size(3'h5),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_ReadAddressChannel_1 sinkBuffered__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(s_axi_ar_ready_0),
		.io_enq_bits_addr(s_axi_ar_bits_addr),
		.io_enq_bits_len(s_axi_ar_bits_len),
		.io_enq_bits_size(3'h5),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	assign s_axi_ar_ready = s_axi_ar_ready_0;
	assign s_axi_r_valid = m_axi_r_valid;
	assign s_axi_r_bits_data = m_axi_r_bits_data;
	assign s_axi_aw_ready = s_axi_aw_ready_0;
	assign s_axi_w_ready = m_axi_w_ready;
	assign s_axi_b_valid = m_axi_b_valid;
	assign m_axi_r_ready = s_axi_r_ready;
	assign m_axi_w_valid = s_axi_w_valid;
	assign m_axi_w_bits_data = s_axi_w_bits_data;
	assign m_axi_w_bits_last = s_axi_w_bits_last;
endmodule
module AxisDataWidthConverter_128 (
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [255:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [255:0] io_dataOut_TDATA;
	assign io_dataIn_TREADY = io_dataOut_TREADY;
	assign io_dataOut_TVALID = io_dataIn_TVALID;
	assign io_dataOut_TDATA = io_dataIn_TDATA;
endmodule
module Scheduler_1 (
	clock,
	reset,
	io_export_taskOut_0_TREADY,
	io_export_taskOut_0_TVALID,
	io_export_taskOut_0_TDATA,
	io_export_taskOut_1_TREADY,
	io_export_taskOut_1_TVALID,
	io_export_taskOut_1_TDATA,
	io_export_taskOut_2_TREADY,
	io_export_taskOut_2_TVALID,
	io_export_taskOut_2_TDATA,
	io_export_taskOut_3_TREADY,
	io_export_taskOut_3_TVALID,
	io_export_taskOut_3_TDATA,
	io_export_taskOut_4_TREADY,
	io_export_taskOut_4_TVALID,
	io_export_taskOut_4_TDATA,
	io_export_taskOut_5_TREADY,
	io_export_taskOut_5_TVALID,
	io_export_taskOut_5_TDATA,
	io_export_taskOut_6_TREADY,
	io_export_taskOut_6_TVALID,
	io_export_taskOut_6_TDATA,
	io_export_taskOut_7_TREADY,
	io_export_taskOut_7_TVALID,
	io_export_taskOut_7_TDATA,
	io_export_taskOut_8_TREADY,
	io_export_taskOut_8_TVALID,
	io_export_taskOut_8_TDATA,
	io_export_taskOut_9_TREADY,
	io_export_taskOut_9_TVALID,
	io_export_taskOut_9_TDATA,
	io_export_taskOut_10_TREADY,
	io_export_taskOut_10_TVALID,
	io_export_taskOut_10_TDATA,
	io_export_taskOut_11_TREADY,
	io_export_taskOut_11_TVALID,
	io_export_taskOut_11_TDATA,
	io_export_taskOut_12_TREADY,
	io_export_taskOut_12_TVALID,
	io_export_taskOut_12_TDATA,
	io_export_taskOut_13_TREADY,
	io_export_taskOut_13_TVALID,
	io_export_taskOut_13_TDATA,
	io_export_taskOut_14_TREADY,
	io_export_taskOut_14_TVALID,
	io_export_taskOut_14_TDATA,
	io_export_taskOut_15_TREADY,
	io_export_taskOut_15_TVALID,
	io_export_taskOut_15_TDATA,
	io_export_taskOut_16_TREADY,
	io_export_taskOut_16_TVALID,
	io_export_taskOut_16_TDATA,
	io_export_taskOut_17_TREADY,
	io_export_taskOut_17_TVALID,
	io_export_taskOut_17_TDATA,
	io_export_taskOut_18_TREADY,
	io_export_taskOut_18_TVALID,
	io_export_taskOut_18_TDATA,
	io_export_taskOut_19_TREADY,
	io_export_taskOut_19_TVALID,
	io_export_taskOut_19_TDATA,
	io_export_taskOut_20_TREADY,
	io_export_taskOut_20_TVALID,
	io_export_taskOut_20_TDATA,
	io_export_taskOut_21_TREADY,
	io_export_taskOut_21_TVALID,
	io_export_taskOut_21_TDATA,
	io_export_taskOut_22_TREADY,
	io_export_taskOut_22_TVALID,
	io_export_taskOut_22_TDATA,
	io_export_taskOut_23_TREADY,
	io_export_taskOut_23_TVALID,
	io_export_taskOut_23_TDATA,
	io_export_taskOut_24_TREADY,
	io_export_taskOut_24_TVALID,
	io_export_taskOut_24_TDATA,
	io_export_taskOut_25_TREADY,
	io_export_taskOut_25_TVALID,
	io_export_taskOut_25_TDATA,
	io_export_taskOut_26_TREADY,
	io_export_taskOut_26_TVALID,
	io_export_taskOut_26_TDATA,
	io_export_taskOut_27_TREADY,
	io_export_taskOut_27_TVALID,
	io_export_taskOut_27_TDATA,
	io_export_taskOut_28_TREADY,
	io_export_taskOut_28_TVALID,
	io_export_taskOut_28_TDATA,
	io_export_taskOut_29_TREADY,
	io_export_taskOut_29_TVALID,
	io_export_taskOut_29_TDATA,
	io_export_taskOut_30_TREADY,
	io_export_taskOut_30_TVALID,
	io_export_taskOut_30_TDATA,
	io_export_taskOut_31_TREADY,
	io_export_taskOut_31_TVALID,
	io_export_taskOut_31_TDATA,
	io_export_taskOut_32_TREADY,
	io_export_taskOut_32_TVALID,
	io_export_taskOut_32_TDATA,
	io_export_taskOut_33_TREADY,
	io_export_taskOut_33_TVALID,
	io_export_taskOut_33_TDATA,
	io_export_taskOut_34_TREADY,
	io_export_taskOut_34_TVALID,
	io_export_taskOut_34_TDATA,
	io_export_taskOut_35_TREADY,
	io_export_taskOut_35_TVALID,
	io_export_taskOut_35_TDATA,
	io_export_taskOut_36_TREADY,
	io_export_taskOut_36_TVALID,
	io_export_taskOut_36_TDATA,
	io_export_taskOut_37_TREADY,
	io_export_taskOut_37_TVALID,
	io_export_taskOut_37_TDATA,
	io_export_taskOut_38_TREADY,
	io_export_taskOut_38_TVALID,
	io_export_taskOut_38_TDATA,
	io_export_taskOut_39_TREADY,
	io_export_taskOut_39_TVALID,
	io_export_taskOut_39_TDATA,
	io_export_taskOut_40_TREADY,
	io_export_taskOut_40_TVALID,
	io_export_taskOut_40_TDATA,
	io_export_taskOut_41_TREADY,
	io_export_taskOut_41_TVALID,
	io_export_taskOut_41_TDATA,
	io_export_taskOut_42_TREADY,
	io_export_taskOut_42_TVALID,
	io_export_taskOut_42_TDATA,
	io_export_taskOut_43_TREADY,
	io_export_taskOut_43_TVALID,
	io_export_taskOut_43_TDATA,
	io_export_taskOut_44_TREADY,
	io_export_taskOut_44_TVALID,
	io_export_taskOut_44_TDATA,
	io_export_taskOut_45_TREADY,
	io_export_taskOut_45_TVALID,
	io_export_taskOut_45_TDATA,
	io_export_taskOut_46_TREADY,
	io_export_taskOut_46_TVALID,
	io_export_taskOut_46_TDATA,
	io_export_taskOut_47_TREADY,
	io_export_taskOut_47_TVALID,
	io_export_taskOut_47_TDATA,
	io_export_taskOut_48_TREADY,
	io_export_taskOut_48_TVALID,
	io_export_taskOut_48_TDATA,
	io_export_taskOut_49_TREADY,
	io_export_taskOut_49_TVALID,
	io_export_taskOut_49_TDATA,
	io_export_taskOut_50_TREADY,
	io_export_taskOut_50_TVALID,
	io_export_taskOut_50_TDATA,
	io_export_taskOut_51_TREADY,
	io_export_taskOut_51_TVALID,
	io_export_taskOut_51_TDATA,
	io_export_taskOut_52_TREADY,
	io_export_taskOut_52_TVALID,
	io_export_taskOut_52_TDATA,
	io_export_taskOut_53_TREADY,
	io_export_taskOut_53_TVALID,
	io_export_taskOut_53_TDATA,
	io_export_taskOut_54_TREADY,
	io_export_taskOut_54_TVALID,
	io_export_taskOut_54_TDATA,
	io_export_taskOut_55_TREADY,
	io_export_taskOut_55_TVALID,
	io_export_taskOut_55_TDATA,
	io_export_taskOut_56_TREADY,
	io_export_taskOut_56_TVALID,
	io_export_taskOut_56_TDATA,
	io_export_taskOut_57_TREADY,
	io_export_taskOut_57_TVALID,
	io_export_taskOut_57_TDATA,
	io_export_taskOut_58_TREADY,
	io_export_taskOut_58_TVALID,
	io_export_taskOut_58_TDATA,
	io_export_taskOut_59_TREADY,
	io_export_taskOut_59_TVALID,
	io_export_taskOut_59_TDATA,
	io_export_taskOut_60_TREADY,
	io_export_taskOut_60_TVALID,
	io_export_taskOut_60_TDATA,
	io_export_taskOut_61_TREADY,
	io_export_taskOut_61_TVALID,
	io_export_taskOut_61_TDATA,
	io_export_taskOut_62_TREADY,
	io_export_taskOut_62_TVALID,
	io_export_taskOut_62_TDATA,
	io_export_taskOut_63_TREADY,
	io_export_taskOut_63_TVALID,
	io_export_taskOut_63_TDATA,
	io_internal_vss_axi_full_0_ar_ready,
	io_internal_vss_axi_full_0_ar_valid,
	io_internal_vss_axi_full_0_ar_bits_id,
	io_internal_vss_axi_full_0_ar_bits_addr,
	io_internal_vss_axi_full_0_ar_bits_len,
	io_internal_vss_axi_full_0_ar_bits_size,
	io_internal_vss_axi_full_0_ar_bits_burst,
	io_internal_vss_axi_full_0_ar_bits_lock,
	io_internal_vss_axi_full_0_ar_bits_cache,
	io_internal_vss_axi_full_0_ar_bits_prot,
	io_internal_vss_axi_full_0_ar_bits_qos,
	io_internal_vss_axi_full_0_ar_bits_region,
	io_internal_vss_axi_full_0_r_ready,
	io_internal_vss_axi_full_0_r_valid,
	io_internal_vss_axi_full_0_r_bits_id,
	io_internal_vss_axi_full_0_r_bits_data,
	io_internal_vss_axi_full_0_r_bits_resp,
	io_internal_vss_axi_full_0_r_bits_last,
	io_internal_vss_axi_full_0_aw_ready,
	io_internal_vss_axi_full_0_aw_valid,
	io_internal_vss_axi_full_0_aw_bits_id,
	io_internal_vss_axi_full_0_aw_bits_addr,
	io_internal_vss_axi_full_0_aw_bits_len,
	io_internal_vss_axi_full_0_aw_bits_size,
	io_internal_vss_axi_full_0_aw_bits_burst,
	io_internal_vss_axi_full_0_aw_bits_lock,
	io_internal_vss_axi_full_0_aw_bits_cache,
	io_internal_vss_axi_full_0_aw_bits_prot,
	io_internal_vss_axi_full_0_aw_bits_qos,
	io_internal_vss_axi_full_0_aw_bits_region,
	io_internal_vss_axi_full_0_w_ready,
	io_internal_vss_axi_full_0_w_valid,
	io_internal_vss_axi_full_0_w_bits_data,
	io_internal_vss_axi_full_0_w_bits_strb,
	io_internal_vss_axi_full_0_w_bits_last,
	io_internal_vss_axi_full_0_b_ready,
	io_internal_vss_axi_full_0_b_valid,
	io_internal_vss_axi_full_0_b_bits_id,
	io_internal_vss_axi_full_0_b_bits_resp,
	io_internal_axi_mgmt_vss_0_ar_ready,
	io_internal_axi_mgmt_vss_0_ar_valid,
	io_internal_axi_mgmt_vss_0_ar_bits_addr,
	io_internal_axi_mgmt_vss_0_ar_bits_prot,
	io_internal_axi_mgmt_vss_0_r_ready,
	io_internal_axi_mgmt_vss_0_r_valid,
	io_internal_axi_mgmt_vss_0_r_bits_data,
	io_internal_axi_mgmt_vss_0_r_bits_resp,
	io_internal_axi_mgmt_vss_0_aw_ready,
	io_internal_axi_mgmt_vss_0_aw_valid,
	io_internal_axi_mgmt_vss_0_aw_bits_addr,
	io_internal_axi_mgmt_vss_0_aw_bits_prot,
	io_internal_axi_mgmt_vss_0_w_ready,
	io_internal_axi_mgmt_vss_0_w_valid,
	io_internal_axi_mgmt_vss_0_w_bits_data,
	io_internal_axi_mgmt_vss_0_w_bits_strb,
	io_internal_axi_mgmt_vss_0_b_ready,
	io_internal_axi_mgmt_vss_0_b_valid,
	io_internal_axi_mgmt_vss_0_b_bits_resp,
	io_internal_axi_mgmt_vss_1_ar_ready,
	io_internal_axi_mgmt_vss_1_ar_valid,
	io_internal_axi_mgmt_vss_1_ar_bits_addr,
	io_internal_axi_mgmt_vss_1_ar_bits_prot,
	io_internal_axi_mgmt_vss_1_r_ready,
	io_internal_axi_mgmt_vss_1_r_valid,
	io_internal_axi_mgmt_vss_1_r_bits_data,
	io_internal_axi_mgmt_vss_1_r_bits_resp,
	io_internal_axi_mgmt_vss_1_aw_ready,
	io_internal_axi_mgmt_vss_1_aw_valid,
	io_internal_axi_mgmt_vss_1_aw_bits_addr,
	io_internal_axi_mgmt_vss_1_aw_bits_prot,
	io_internal_axi_mgmt_vss_1_w_ready,
	io_internal_axi_mgmt_vss_1_w_valid,
	io_internal_axi_mgmt_vss_1_w_bits_data,
	io_internal_axi_mgmt_vss_1_w_bits_strb,
	io_internal_axi_mgmt_vss_1_b_ready,
	io_internal_axi_mgmt_vss_1_b_valid,
	io_internal_axi_mgmt_vss_1_b_bits_resp,
	connArgumentNotifier_0_ctrl_serveStealReq_valid,
	connArgumentNotifier_0_ctrl_serveStealReq_ready,
	connArgumentNotifier_0_data_qOutTask_ready,
	connArgumentNotifier_0_data_qOutTask_valid,
	connArgumentNotifier_0_data_qOutTask_bits,
	connArgumentNotifier_1_ctrl_serveStealReq_valid,
	connArgumentNotifier_1_ctrl_serveStealReq_ready,
	connArgumentNotifier_1_data_qOutTask_ready,
	connArgumentNotifier_1_data_qOutTask_valid,
	connArgumentNotifier_1_data_qOutTask_bits,
	connArgumentNotifier_2_ctrl_serveStealReq_valid,
	connArgumentNotifier_2_ctrl_serveStealReq_ready,
	connArgumentNotifier_2_data_qOutTask_ready,
	connArgumentNotifier_2_data_qOutTask_valid,
	connArgumentNotifier_2_data_qOutTask_bits,
	connArgumentNotifier_3_ctrl_serveStealReq_valid,
	connArgumentNotifier_3_ctrl_serveStealReq_ready,
	connArgumentNotifier_3_data_qOutTask_ready,
	connArgumentNotifier_3_data_qOutTask_valid,
	connArgumentNotifier_3_data_qOutTask_bits,
	connArgumentNotifier_4_ctrl_serveStealReq_valid,
	connArgumentNotifier_4_ctrl_serveStealReq_ready,
	connArgumentNotifier_4_data_qOutTask_ready,
	connArgumentNotifier_4_data_qOutTask_valid,
	connArgumentNotifier_4_data_qOutTask_bits,
	connArgumentNotifier_5_ctrl_serveStealReq_valid,
	connArgumentNotifier_5_ctrl_serveStealReq_ready,
	connArgumentNotifier_5_data_qOutTask_ready,
	connArgumentNotifier_5_data_qOutTask_valid,
	connArgumentNotifier_5_data_qOutTask_bits,
	connArgumentNotifier_6_ctrl_serveStealReq_valid,
	connArgumentNotifier_6_ctrl_serveStealReq_ready,
	connArgumentNotifier_6_data_qOutTask_ready,
	connArgumentNotifier_6_data_qOutTask_valid,
	connArgumentNotifier_6_data_qOutTask_bits,
	connArgumentNotifier_7_ctrl_serveStealReq_valid,
	connArgumentNotifier_7_ctrl_serveStealReq_ready,
	connArgumentNotifier_7_data_qOutTask_ready,
	connArgumentNotifier_7_data_qOutTask_valid,
	connArgumentNotifier_7_data_qOutTask_bits,
	connArgumentNotifier_8_ctrl_serveStealReq_valid,
	connArgumentNotifier_8_ctrl_serveStealReq_ready,
	connArgumentNotifier_8_data_qOutTask_ready,
	connArgumentNotifier_8_data_qOutTask_valid,
	connArgumentNotifier_8_data_qOutTask_bits,
	connArgumentNotifier_9_ctrl_serveStealReq_valid,
	connArgumentNotifier_9_ctrl_serveStealReq_ready,
	connArgumentNotifier_9_data_qOutTask_ready,
	connArgumentNotifier_9_data_qOutTask_valid,
	connArgumentNotifier_9_data_qOutTask_bits,
	connArgumentNotifier_10_ctrl_serveStealReq_valid,
	connArgumentNotifier_10_ctrl_serveStealReq_ready,
	connArgumentNotifier_10_data_qOutTask_ready,
	connArgumentNotifier_10_data_qOutTask_valid,
	connArgumentNotifier_10_data_qOutTask_bits,
	connArgumentNotifier_11_ctrl_serveStealReq_valid,
	connArgumentNotifier_11_ctrl_serveStealReq_ready,
	connArgumentNotifier_11_data_qOutTask_ready,
	connArgumentNotifier_11_data_qOutTask_valid,
	connArgumentNotifier_11_data_qOutTask_bits,
	connArgumentNotifier_12_ctrl_serveStealReq_valid,
	connArgumentNotifier_12_ctrl_serveStealReq_ready,
	connArgumentNotifier_12_data_qOutTask_ready,
	connArgumentNotifier_12_data_qOutTask_valid,
	connArgumentNotifier_12_data_qOutTask_bits,
	connArgumentNotifier_13_ctrl_serveStealReq_valid,
	connArgumentNotifier_13_ctrl_serveStealReq_ready,
	connArgumentNotifier_13_data_qOutTask_ready,
	connArgumentNotifier_13_data_qOutTask_valid,
	connArgumentNotifier_13_data_qOutTask_bits,
	connArgumentNotifier_14_ctrl_serveStealReq_valid,
	connArgumentNotifier_14_ctrl_serveStealReq_ready,
	connArgumentNotifier_14_data_qOutTask_ready,
	connArgumentNotifier_14_data_qOutTask_valid,
	connArgumentNotifier_14_data_qOutTask_bits,
	connArgumentNotifier_15_ctrl_serveStealReq_valid,
	connArgumentNotifier_15_ctrl_serveStealReq_ready,
	connArgumentNotifier_15_data_qOutTask_ready,
	connArgumentNotifier_15_data_qOutTask_valid,
	connArgumentNotifier_15_data_qOutTask_bits
);
	input clock;
	input reset;
	input io_export_taskOut_0_TREADY;
	output wire io_export_taskOut_0_TVALID;
	output wire [255:0] io_export_taskOut_0_TDATA;
	input io_export_taskOut_1_TREADY;
	output wire io_export_taskOut_1_TVALID;
	output wire [255:0] io_export_taskOut_1_TDATA;
	input io_export_taskOut_2_TREADY;
	output wire io_export_taskOut_2_TVALID;
	output wire [255:0] io_export_taskOut_2_TDATA;
	input io_export_taskOut_3_TREADY;
	output wire io_export_taskOut_3_TVALID;
	output wire [255:0] io_export_taskOut_3_TDATA;
	input io_export_taskOut_4_TREADY;
	output wire io_export_taskOut_4_TVALID;
	output wire [255:0] io_export_taskOut_4_TDATA;
	input io_export_taskOut_5_TREADY;
	output wire io_export_taskOut_5_TVALID;
	output wire [255:0] io_export_taskOut_5_TDATA;
	input io_export_taskOut_6_TREADY;
	output wire io_export_taskOut_6_TVALID;
	output wire [255:0] io_export_taskOut_6_TDATA;
	input io_export_taskOut_7_TREADY;
	output wire io_export_taskOut_7_TVALID;
	output wire [255:0] io_export_taskOut_7_TDATA;
	input io_export_taskOut_8_TREADY;
	output wire io_export_taskOut_8_TVALID;
	output wire [255:0] io_export_taskOut_8_TDATA;
	input io_export_taskOut_9_TREADY;
	output wire io_export_taskOut_9_TVALID;
	output wire [255:0] io_export_taskOut_9_TDATA;
	input io_export_taskOut_10_TREADY;
	output wire io_export_taskOut_10_TVALID;
	output wire [255:0] io_export_taskOut_10_TDATA;
	input io_export_taskOut_11_TREADY;
	output wire io_export_taskOut_11_TVALID;
	output wire [255:0] io_export_taskOut_11_TDATA;
	input io_export_taskOut_12_TREADY;
	output wire io_export_taskOut_12_TVALID;
	output wire [255:0] io_export_taskOut_12_TDATA;
	input io_export_taskOut_13_TREADY;
	output wire io_export_taskOut_13_TVALID;
	output wire [255:0] io_export_taskOut_13_TDATA;
	input io_export_taskOut_14_TREADY;
	output wire io_export_taskOut_14_TVALID;
	output wire [255:0] io_export_taskOut_14_TDATA;
	input io_export_taskOut_15_TREADY;
	output wire io_export_taskOut_15_TVALID;
	output wire [255:0] io_export_taskOut_15_TDATA;
	input io_export_taskOut_16_TREADY;
	output wire io_export_taskOut_16_TVALID;
	output wire [255:0] io_export_taskOut_16_TDATA;
	input io_export_taskOut_17_TREADY;
	output wire io_export_taskOut_17_TVALID;
	output wire [255:0] io_export_taskOut_17_TDATA;
	input io_export_taskOut_18_TREADY;
	output wire io_export_taskOut_18_TVALID;
	output wire [255:0] io_export_taskOut_18_TDATA;
	input io_export_taskOut_19_TREADY;
	output wire io_export_taskOut_19_TVALID;
	output wire [255:0] io_export_taskOut_19_TDATA;
	input io_export_taskOut_20_TREADY;
	output wire io_export_taskOut_20_TVALID;
	output wire [255:0] io_export_taskOut_20_TDATA;
	input io_export_taskOut_21_TREADY;
	output wire io_export_taskOut_21_TVALID;
	output wire [255:0] io_export_taskOut_21_TDATA;
	input io_export_taskOut_22_TREADY;
	output wire io_export_taskOut_22_TVALID;
	output wire [255:0] io_export_taskOut_22_TDATA;
	input io_export_taskOut_23_TREADY;
	output wire io_export_taskOut_23_TVALID;
	output wire [255:0] io_export_taskOut_23_TDATA;
	input io_export_taskOut_24_TREADY;
	output wire io_export_taskOut_24_TVALID;
	output wire [255:0] io_export_taskOut_24_TDATA;
	input io_export_taskOut_25_TREADY;
	output wire io_export_taskOut_25_TVALID;
	output wire [255:0] io_export_taskOut_25_TDATA;
	input io_export_taskOut_26_TREADY;
	output wire io_export_taskOut_26_TVALID;
	output wire [255:0] io_export_taskOut_26_TDATA;
	input io_export_taskOut_27_TREADY;
	output wire io_export_taskOut_27_TVALID;
	output wire [255:0] io_export_taskOut_27_TDATA;
	input io_export_taskOut_28_TREADY;
	output wire io_export_taskOut_28_TVALID;
	output wire [255:0] io_export_taskOut_28_TDATA;
	input io_export_taskOut_29_TREADY;
	output wire io_export_taskOut_29_TVALID;
	output wire [255:0] io_export_taskOut_29_TDATA;
	input io_export_taskOut_30_TREADY;
	output wire io_export_taskOut_30_TVALID;
	output wire [255:0] io_export_taskOut_30_TDATA;
	input io_export_taskOut_31_TREADY;
	output wire io_export_taskOut_31_TVALID;
	output wire [255:0] io_export_taskOut_31_TDATA;
	input io_export_taskOut_32_TREADY;
	output wire io_export_taskOut_32_TVALID;
	output wire [255:0] io_export_taskOut_32_TDATA;
	input io_export_taskOut_33_TREADY;
	output wire io_export_taskOut_33_TVALID;
	output wire [255:0] io_export_taskOut_33_TDATA;
	input io_export_taskOut_34_TREADY;
	output wire io_export_taskOut_34_TVALID;
	output wire [255:0] io_export_taskOut_34_TDATA;
	input io_export_taskOut_35_TREADY;
	output wire io_export_taskOut_35_TVALID;
	output wire [255:0] io_export_taskOut_35_TDATA;
	input io_export_taskOut_36_TREADY;
	output wire io_export_taskOut_36_TVALID;
	output wire [255:0] io_export_taskOut_36_TDATA;
	input io_export_taskOut_37_TREADY;
	output wire io_export_taskOut_37_TVALID;
	output wire [255:0] io_export_taskOut_37_TDATA;
	input io_export_taskOut_38_TREADY;
	output wire io_export_taskOut_38_TVALID;
	output wire [255:0] io_export_taskOut_38_TDATA;
	input io_export_taskOut_39_TREADY;
	output wire io_export_taskOut_39_TVALID;
	output wire [255:0] io_export_taskOut_39_TDATA;
	input io_export_taskOut_40_TREADY;
	output wire io_export_taskOut_40_TVALID;
	output wire [255:0] io_export_taskOut_40_TDATA;
	input io_export_taskOut_41_TREADY;
	output wire io_export_taskOut_41_TVALID;
	output wire [255:0] io_export_taskOut_41_TDATA;
	input io_export_taskOut_42_TREADY;
	output wire io_export_taskOut_42_TVALID;
	output wire [255:0] io_export_taskOut_42_TDATA;
	input io_export_taskOut_43_TREADY;
	output wire io_export_taskOut_43_TVALID;
	output wire [255:0] io_export_taskOut_43_TDATA;
	input io_export_taskOut_44_TREADY;
	output wire io_export_taskOut_44_TVALID;
	output wire [255:0] io_export_taskOut_44_TDATA;
	input io_export_taskOut_45_TREADY;
	output wire io_export_taskOut_45_TVALID;
	output wire [255:0] io_export_taskOut_45_TDATA;
	input io_export_taskOut_46_TREADY;
	output wire io_export_taskOut_46_TVALID;
	output wire [255:0] io_export_taskOut_46_TDATA;
	input io_export_taskOut_47_TREADY;
	output wire io_export_taskOut_47_TVALID;
	output wire [255:0] io_export_taskOut_47_TDATA;
	input io_export_taskOut_48_TREADY;
	output wire io_export_taskOut_48_TVALID;
	output wire [255:0] io_export_taskOut_48_TDATA;
	input io_export_taskOut_49_TREADY;
	output wire io_export_taskOut_49_TVALID;
	output wire [255:0] io_export_taskOut_49_TDATA;
	input io_export_taskOut_50_TREADY;
	output wire io_export_taskOut_50_TVALID;
	output wire [255:0] io_export_taskOut_50_TDATA;
	input io_export_taskOut_51_TREADY;
	output wire io_export_taskOut_51_TVALID;
	output wire [255:0] io_export_taskOut_51_TDATA;
	input io_export_taskOut_52_TREADY;
	output wire io_export_taskOut_52_TVALID;
	output wire [255:0] io_export_taskOut_52_TDATA;
	input io_export_taskOut_53_TREADY;
	output wire io_export_taskOut_53_TVALID;
	output wire [255:0] io_export_taskOut_53_TDATA;
	input io_export_taskOut_54_TREADY;
	output wire io_export_taskOut_54_TVALID;
	output wire [255:0] io_export_taskOut_54_TDATA;
	input io_export_taskOut_55_TREADY;
	output wire io_export_taskOut_55_TVALID;
	output wire [255:0] io_export_taskOut_55_TDATA;
	input io_export_taskOut_56_TREADY;
	output wire io_export_taskOut_56_TVALID;
	output wire [255:0] io_export_taskOut_56_TDATA;
	input io_export_taskOut_57_TREADY;
	output wire io_export_taskOut_57_TVALID;
	output wire [255:0] io_export_taskOut_57_TDATA;
	input io_export_taskOut_58_TREADY;
	output wire io_export_taskOut_58_TVALID;
	output wire [255:0] io_export_taskOut_58_TDATA;
	input io_export_taskOut_59_TREADY;
	output wire io_export_taskOut_59_TVALID;
	output wire [255:0] io_export_taskOut_59_TDATA;
	input io_export_taskOut_60_TREADY;
	output wire io_export_taskOut_60_TVALID;
	output wire [255:0] io_export_taskOut_60_TDATA;
	input io_export_taskOut_61_TREADY;
	output wire io_export_taskOut_61_TVALID;
	output wire [255:0] io_export_taskOut_61_TDATA;
	input io_export_taskOut_62_TREADY;
	output wire io_export_taskOut_62_TVALID;
	output wire [255:0] io_export_taskOut_62_TDATA;
	input io_export_taskOut_63_TREADY;
	output wire io_export_taskOut_63_TVALID;
	output wire [255:0] io_export_taskOut_63_TDATA;
	input io_internal_vss_axi_full_0_ar_ready;
	output wire io_internal_vss_axi_full_0_ar_valid;
	output wire [1:0] io_internal_vss_axi_full_0_ar_bits_id;
	output wire [63:0] io_internal_vss_axi_full_0_ar_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_ar_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_ar_bits_burst;
	output wire io_internal_vss_axi_full_0_ar_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_region;
	output wire io_internal_vss_axi_full_0_r_ready;
	input io_internal_vss_axi_full_0_r_valid;
	input [1:0] io_internal_vss_axi_full_0_r_bits_id;
	input [255:0] io_internal_vss_axi_full_0_r_bits_data;
	input [1:0] io_internal_vss_axi_full_0_r_bits_resp;
	input io_internal_vss_axi_full_0_r_bits_last;
	input io_internal_vss_axi_full_0_aw_ready;
	output wire io_internal_vss_axi_full_0_aw_valid;
	output wire [1:0] io_internal_vss_axi_full_0_aw_bits_id;
	output wire [63:0] io_internal_vss_axi_full_0_aw_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_aw_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_aw_bits_burst;
	output wire io_internal_vss_axi_full_0_aw_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_region;
	input io_internal_vss_axi_full_0_w_ready;
	output wire io_internal_vss_axi_full_0_w_valid;
	output wire [255:0] io_internal_vss_axi_full_0_w_bits_data;
	output wire [31:0] io_internal_vss_axi_full_0_w_bits_strb;
	output wire io_internal_vss_axi_full_0_w_bits_last;
	output wire io_internal_vss_axi_full_0_b_ready;
	input io_internal_vss_axi_full_0_b_valid;
	input [1:0] io_internal_vss_axi_full_0_b_bits_id;
	input [1:0] io_internal_vss_axi_full_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vss_0_ar_ready;
	input io_internal_axi_mgmt_vss_0_ar_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_ar_bits_prot;
	input io_internal_axi_mgmt_vss_0_r_ready;
	output wire io_internal_axi_mgmt_vss_0_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vss_0_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vss_0_r_bits_resp;
	output wire io_internal_axi_mgmt_vss_0_aw_ready;
	input io_internal_axi_mgmt_vss_0_aw_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_aw_bits_prot;
	output wire io_internal_axi_mgmt_vss_0_w_ready;
	input io_internal_axi_mgmt_vss_0_w_valid;
	input [63:0] io_internal_axi_mgmt_vss_0_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vss_0_w_bits_strb;
	input io_internal_axi_mgmt_vss_0_b_ready;
	output wire io_internal_axi_mgmt_vss_0_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vss_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vss_1_ar_ready;
	input io_internal_axi_mgmt_vss_1_ar_valid;
	input [5:0] io_internal_axi_mgmt_vss_1_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_1_ar_bits_prot;
	input io_internal_axi_mgmt_vss_1_r_ready;
	output wire io_internal_axi_mgmt_vss_1_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vss_1_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vss_1_r_bits_resp;
	output wire io_internal_axi_mgmt_vss_1_aw_ready;
	input io_internal_axi_mgmt_vss_1_aw_valid;
	input [5:0] io_internal_axi_mgmt_vss_1_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_1_aw_bits_prot;
	output wire io_internal_axi_mgmt_vss_1_w_ready;
	input io_internal_axi_mgmt_vss_1_w_valid;
	input [63:0] io_internal_axi_mgmt_vss_1_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vss_1_w_bits_strb;
	input io_internal_axi_mgmt_vss_1_b_ready;
	output wire io_internal_axi_mgmt_vss_1_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vss_1_b_bits_resp;
	input connArgumentNotifier_0_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_0_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_0_data_qOutTask_ready;
	input connArgumentNotifier_0_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_0_data_qOutTask_bits;
	input connArgumentNotifier_1_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_1_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_1_data_qOutTask_ready;
	input connArgumentNotifier_1_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_1_data_qOutTask_bits;
	input connArgumentNotifier_2_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_2_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_2_data_qOutTask_ready;
	input connArgumentNotifier_2_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_2_data_qOutTask_bits;
	input connArgumentNotifier_3_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_3_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_3_data_qOutTask_ready;
	input connArgumentNotifier_3_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_3_data_qOutTask_bits;
	input connArgumentNotifier_4_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_4_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_4_data_qOutTask_ready;
	input connArgumentNotifier_4_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_4_data_qOutTask_bits;
	input connArgumentNotifier_5_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_5_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_5_data_qOutTask_ready;
	input connArgumentNotifier_5_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_5_data_qOutTask_bits;
	input connArgumentNotifier_6_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_6_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_6_data_qOutTask_ready;
	input connArgumentNotifier_6_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_6_data_qOutTask_bits;
	input connArgumentNotifier_7_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_7_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_7_data_qOutTask_ready;
	input connArgumentNotifier_7_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_7_data_qOutTask_bits;
	input connArgumentNotifier_8_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_8_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_8_data_qOutTask_ready;
	input connArgumentNotifier_8_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_8_data_qOutTask_bits;
	input connArgumentNotifier_9_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_9_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_9_data_qOutTask_ready;
	input connArgumentNotifier_9_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_9_data_qOutTask_bits;
	input connArgumentNotifier_10_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_10_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_10_data_qOutTask_ready;
	input connArgumentNotifier_10_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_10_data_qOutTask_bits;
	input connArgumentNotifier_11_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_11_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_11_data_qOutTask_ready;
	input connArgumentNotifier_11_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_11_data_qOutTask_bits;
	input connArgumentNotifier_12_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_12_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_12_data_qOutTask_ready;
	input connArgumentNotifier_12_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_12_data_qOutTask_bits;
	input connArgumentNotifier_13_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_13_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_13_data_qOutTask_ready;
	input connArgumentNotifier_13_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_13_data_qOutTask_bits;
	input connArgumentNotifier_14_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_14_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_14_data_qOutTask_ready;
	input connArgumentNotifier_14_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_14_data_qOutTask_bits;
	input connArgumentNotifier_15_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_15_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_15_data_qOutTask_ready;
	input connArgumentNotifier_15_data_qOutTask_valid;
	input [255:0] connArgumentNotifier_15_data_qOutTask_bits;
	wire _axis_stream_converters_out_63_io_dataIn_TREADY;
	wire _axis_stream_converters_out_62_io_dataIn_TREADY;
	wire _axis_stream_converters_out_61_io_dataIn_TREADY;
	wire _axis_stream_converters_out_60_io_dataIn_TREADY;
	wire _axis_stream_converters_out_59_io_dataIn_TREADY;
	wire _axis_stream_converters_out_58_io_dataIn_TREADY;
	wire _axis_stream_converters_out_57_io_dataIn_TREADY;
	wire _axis_stream_converters_out_56_io_dataIn_TREADY;
	wire _axis_stream_converters_out_55_io_dataIn_TREADY;
	wire _axis_stream_converters_out_54_io_dataIn_TREADY;
	wire _axis_stream_converters_out_53_io_dataIn_TREADY;
	wire _axis_stream_converters_out_52_io_dataIn_TREADY;
	wire _axis_stream_converters_out_51_io_dataIn_TREADY;
	wire _axis_stream_converters_out_50_io_dataIn_TREADY;
	wire _axis_stream_converters_out_49_io_dataIn_TREADY;
	wire _axis_stream_converters_out_48_io_dataIn_TREADY;
	wire _axis_stream_converters_out_47_io_dataIn_TREADY;
	wire _axis_stream_converters_out_46_io_dataIn_TREADY;
	wire _axis_stream_converters_out_45_io_dataIn_TREADY;
	wire _axis_stream_converters_out_44_io_dataIn_TREADY;
	wire _axis_stream_converters_out_43_io_dataIn_TREADY;
	wire _axis_stream_converters_out_42_io_dataIn_TREADY;
	wire _axis_stream_converters_out_41_io_dataIn_TREADY;
	wire _axis_stream_converters_out_40_io_dataIn_TREADY;
	wire _axis_stream_converters_out_39_io_dataIn_TREADY;
	wire _axis_stream_converters_out_38_io_dataIn_TREADY;
	wire _axis_stream_converters_out_37_io_dataIn_TREADY;
	wire _axis_stream_converters_out_36_io_dataIn_TREADY;
	wire _axis_stream_converters_out_35_io_dataIn_TREADY;
	wire _axis_stream_converters_out_34_io_dataIn_TREADY;
	wire _axis_stream_converters_out_33_io_dataIn_TREADY;
	wire _axis_stream_converters_out_32_io_dataIn_TREADY;
	wire _axis_stream_converters_out_31_io_dataIn_TREADY;
	wire _axis_stream_converters_out_30_io_dataIn_TREADY;
	wire _axis_stream_converters_out_29_io_dataIn_TREADY;
	wire _axis_stream_converters_out_28_io_dataIn_TREADY;
	wire _axis_stream_converters_out_27_io_dataIn_TREADY;
	wire _axis_stream_converters_out_26_io_dataIn_TREADY;
	wire _axis_stream_converters_out_25_io_dataIn_TREADY;
	wire _axis_stream_converters_out_24_io_dataIn_TREADY;
	wire _axis_stream_converters_out_23_io_dataIn_TREADY;
	wire _axis_stream_converters_out_22_io_dataIn_TREADY;
	wire _axis_stream_converters_out_21_io_dataIn_TREADY;
	wire _axis_stream_converters_out_20_io_dataIn_TREADY;
	wire _axis_stream_converters_out_19_io_dataIn_TREADY;
	wire _axis_stream_converters_out_18_io_dataIn_TREADY;
	wire _axis_stream_converters_out_17_io_dataIn_TREADY;
	wire _axis_stream_converters_out_16_io_dataIn_TREADY;
	wire _axis_stream_converters_out_15_io_dataIn_TREADY;
	wire _axis_stream_converters_out_14_io_dataIn_TREADY;
	wire _axis_stream_converters_out_13_io_dataIn_TREADY;
	wire _axis_stream_converters_out_12_io_dataIn_TREADY;
	wire _axis_stream_converters_out_11_io_dataIn_TREADY;
	wire _axis_stream_converters_out_10_io_dataIn_TREADY;
	wire _axis_stream_converters_out_9_io_dataIn_TREADY;
	wire _axis_stream_converters_out_8_io_dataIn_TREADY;
	wire _axis_stream_converters_out_7_io_dataIn_TREADY;
	wire _axis_stream_converters_out_6_io_dataIn_TREADY;
	wire _axis_stream_converters_out_5_io_dataIn_TREADY;
	wire _axis_stream_converters_out_4_io_dataIn_TREADY;
	wire _axis_stream_converters_out_3_io_dataIn_TREADY;
	wire _axis_stream_converters_out_2_io_dataIn_TREADY;
	wire _axis_stream_converters_out_1_io_dataIn_TREADY;
	wire _axis_stream_converters_out_0_io_dataIn_TREADY;
	wire _module_1_s_axi_ar_ready;
	wire _module_1_s_axi_r_valid;
	wire [255:0] _module_1_s_axi_r_bits_data;
	wire _module_1_s_axi_aw_ready;
	wire _module_1_s_axi_w_ready;
	wire _module_1_s_axi_b_valid;
	wire _module_1_m_axi_ar_valid;
	wire [63:0] _module_1_m_axi_ar_bits_addr;
	wire [7:0] _module_1_m_axi_ar_bits_len;
	wire [2:0] _module_1_m_axi_ar_bits_size;
	wire [1:0] _module_1_m_axi_ar_bits_burst;
	wire _module_1_m_axi_ar_bits_lock;
	wire [3:0] _module_1_m_axi_ar_bits_cache;
	wire [2:0] _module_1_m_axi_ar_bits_prot;
	wire [3:0] _module_1_m_axi_ar_bits_qos;
	wire [3:0] _module_1_m_axi_ar_bits_region;
	wire _module_1_m_axi_r_ready;
	wire _module_1_m_axi_aw_valid;
	wire [63:0] _module_1_m_axi_aw_bits_addr;
	wire [7:0] _module_1_m_axi_aw_bits_len;
	wire [2:0] _module_1_m_axi_aw_bits_size;
	wire [1:0] _module_1_m_axi_aw_bits_burst;
	wire _module_1_m_axi_aw_bits_lock;
	wire [3:0] _module_1_m_axi_aw_bits_cache;
	wire [2:0] _module_1_m_axi_aw_bits_prot;
	wire [3:0] _module_1_m_axi_aw_bits_qos;
	wire [3:0] _module_1_m_axi_aw_bits_region;
	wire _module_1_m_axi_w_valid;
	wire [255:0] _module_1_m_axi_w_bits_data;
	wire _module_1_m_axi_w_bits_last;
	wire _module_s_axi_ar_ready;
	wire _module_s_axi_r_valid;
	wire [255:0] _module_s_axi_r_bits_data;
	wire _module_s_axi_aw_ready;
	wire _module_s_axi_w_ready;
	wire _module_s_axi_b_valid;
	wire _module_m_axi_ar_valid;
	wire [63:0] _module_m_axi_ar_bits_addr;
	wire [7:0] _module_m_axi_ar_bits_len;
	wire [2:0] _module_m_axi_ar_bits_size;
	wire [1:0] _module_m_axi_ar_bits_burst;
	wire _module_m_axi_ar_bits_lock;
	wire [3:0] _module_m_axi_ar_bits_cache;
	wire [2:0] _module_m_axi_ar_bits_prot;
	wire [3:0] _module_m_axi_ar_bits_qos;
	wire [3:0] _module_m_axi_ar_bits_region;
	wire _module_m_axi_r_ready;
	wire _module_m_axi_aw_valid;
	wire [63:0] _module_m_axi_aw_bits_addr;
	wire [7:0] _module_m_axi_aw_bits_len;
	wire [2:0] _module_m_axi_aw_bits_size;
	wire [1:0] _module_m_axi_aw_bits_burst;
	wire _module_m_axi_aw_bits_lock;
	wire [3:0] _module_m_axi_aw_bits_cache;
	wire [2:0] _module_m_axi_aw_bits_prot;
	wire [3:0] _module_m_axi_aw_bits_qos;
	wire [3:0] _module_m_axi_aw_bits_region;
	wire _module_m_axi_w_valid;
	wire [255:0] _module_m_axi_w_bits_data;
	wire _module_m_axi_w_bits_last;
	wire _mux_s_axi_0_ar_ready;
	wire _mux_s_axi_0_r_valid;
	wire [255:0] _mux_s_axi_0_r_bits_data;
	wire _mux_s_axi_0_aw_ready;
	wire _mux_s_axi_0_w_ready;
	wire _mux_s_axi_0_b_valid;
	wire _mux_s_axi_1_ar_ready;
	wire _mux_s_axi_1_r_valid;
	wire [255:0] _mux_s_axi_1_r_bits_data;
	wire _mux_s_axi_1_aw_ready;
	wire _mux_s_axi_1_w_ready;
	wire _mux_s_axi_1_b_valid;
	wire _vssRvm_1_io_read_address_ready;
	wire _vssRvm_1_io_read_data_valid;
	wire [255:0] _vssRvm_1_io_read_data_bits;
	wire _vssRvm_1_io_write_address_ready;
	wire _vssRvm_1_io_write_data_ready;
	wire _vssRvm_1_axi_ar_valid;
	wire [63:0] _vssRvm_1_axi_ar_bits_addr;
	wire [7:0] _vssRvm_1_axi_ar_bits_len;
	wire _vssRvm_1_axi_r_ready;
	wire _vssRvm_1_axi_aw_valid;
	wire [63:0] _vssRvm_1_axi_aw_bits_addr;
	wire [7:0] _vssRvm_1_axi_aw_bits_len;
	wire _vssRvm_1_axi_w_valid;
	wire [255:0] _vssRvm_1_axi_w_bits_data;
	wire _vssRvm_1_axi_w_bits_last;
	wire _vssRvm_0_io_read_address_ready;
	wire _vssRvm_0_io_read_data_valid;
	wire [255:0] _vssRvm_0_io_read_data_bits;
	wire _vssRvm_0_io_write_address_ready;
	wire _vssRvm_0_io_write_data_ready;
	wire _vssRvm_0_axi_ar_valid;
	wire [63:0] _vssRvm_0_axi_ar_bits_addr;
	wire [7:0] _vssRvm_0_axi_ar_bits_len;
	wire _vssRvm_0_axi_r_ready;
	wire _vssRvm_0_axi_aw_valid;
	wire [63:0] _vssRvm_0_axi_aw_bits_addr;
	wire [7:0] _vssRvm_0_axi_aw_bits_len;
	wire _vssRvm_0_axi_w_valid;
	wire [255:0] _vssRvm_0_axi_w_bits_data;
	wire _vssRvm_0_axi_w_bits_last;
	wire _virtualStealServers_1_io_connNetwork_ctrl_serveStealReq_valid;
	wire _virtualStealServers_1_io_connNetwork_data_availableTask_ready;
	wire _virtualStealServers_1_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _virtualStealServers_1_io_connNetwork_data_qOutTask_bits;
	wire _virtualStealServers_1_io_read_address_valid;
	wire [63:0] _virtualStealServers_1_io_read_address_bits;
	wire _virtualStealServers_1_io_read_data_ready;
	wire [3:0] _virtualStealServers_1_io_read_burst_len;
	wire _virtualStealServers_1_io_write_address_valid;
	wire [63:0] _virtualStealServers_1_io_write_address_bits;
	wire _virtualStealServers_1_io_write_data_valid;
	wire [255:0] _virtualStealServers_1_io_write_data_bits;
	wire [3:0] _virtualStealServers_1_io_write_burst_len;
	wire _virtualStealServers_1_io_write_last;
	wire _virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _virtualStealServers_0_io_connNetwork_data_availableTask_ready;
	wire _virtualStealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _virtualStealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _virtualStealServers_0_io_read_address_valid;
	wire [63:0] _virtualStealServers_0_io_read_address_bits;
	wire _virtualStealServers_0_io_read_data_ready;
	wire [3:0] _virtualStealServers_0_io_read_burst_len;
	wire _virtualStealServers_0_io_write_address_valid;
	wire [63:0] _virtualStealServers_0_io_write_address_bits;
	wire _virtualStealServers_0_io_write_data_valid;
	wire [255:0] _virtualStealServers_0_io_write_data_bits;
	wire [3:0] _virtualStealServers_0_io_write_burst_len;
	wire _virtualStealServers_0_io_write_last;
	wire _stealNW_TQ_io_connPE_0_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_0_pop_bits;
	wire _stealNW_TQ_io_connPE_1_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_1_pop_bits;
	wire _stealNW_TQ_io_connPE_2_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_2_pop_bits;
	wire _stealNW_TQ_io_connPE_3_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_3_pop_bits;
	wire _stealNW_TQ_io_connPE_4_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_4_pop_bits;
	wire _stealNW_TQ_io_connPE_5_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_5_pop_bits;
	wire _stealNW_TQ_io_connPE_6_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_6_pop_bits;
	wire _stealNW_TQ_io_connPE_7_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_7_pop_bits;
	wire _stealNW_TQ_io_connPE_8_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_8_pop_bits;
	wire _stealNW_TQ_io_connPE_9_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_9_pop_bits;
	wire _stealNW_TQ_io_connPE_10_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_10_pop_bits;
	wire _stealNW_TQ_io_connPE_11_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_11_pop_bits;
	wire _stealNW_TQ_io_connPE_12_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_12_pop_bits;
	wire _stealNW_TQ_io_connPE_13_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_13_pop_bits;
	wire _stealNW_TQ_io_connPE_14_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_14_pop_bits;
	wire _stealNW_TQ_io_connPE_15_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_15_pop_bits;
	wire _stealNW_TQ_io_connPE_16_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_16_pop_bits;
	wire _stealNW_TQ_io_connPE_17_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_17_pop_bits;
	wire _stealNW_TQ_io_connPE_18_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_18_pop_bits;
	wire _stealNW_TQ_io_connPE_19_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_19_pop_bits;
	wire _stealNW_TQ_io_connPE_20_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_20_pop_bits;
	wire _stealNW_TQ_io_connPE_21_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_21_pop_bits;
	wire _stealNW_TQ_io_connPE_22_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_22_pop_bits;
	wire _stealNW_TQ_io_connPE_23_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_23_pop_bits;
	wire _stealNW_TQ_io_connPE_24_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_24_pop_bits;
	wire _stealNW_TQ_io_connPE_25_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_25_pop_bits;
	wire _stealNW_TQ_io_connPE_26_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_26_pop_bits;
	wire _stealNW_TQ_io_connPE_27_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_27_pop_bits;
	wire _stealNW_TQ_io_connPE_28_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_28_pop_bits;
	wire _stealNW_TQ_io_connPE_29_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_29_pop_bits;
	wire _stealNW_TQ_io_connPE_30_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_30_pop_bits;
	wire _stealNW_TQ_io_connPE_31_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_31_pop_bits;
	wire _stealNW_TQ_io_connPE_32_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_32_pop_bits;
	wire _stealNW_TQ_io_connPE_33_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_33_pop_bits;
	wire _stealNW_TQ_io_connPE_34_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_34_pop_bits;
	wire _stealNW_TQ_io_connPE_35_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_35_pop_bits;
	wire _stealNW_TQ_io_connPE_36_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_36_pop_bits;
	wire _stealNW_TQ_io_connPE_37_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_37_pop_bits;
	wire _stealNW_TQ_io_connPE_38_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_38_pop_bits;
	wire _stealNW_TQ_io_connPE_39_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_39_pop_bits;
	wire _stealNW_TQ_io_connPE_40_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_40_pop_bits;
	wire _stealNW_TQ_io_connPE_41_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_41_pop_bits;
	wire _stealNW_TQ_io_connPE_42_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_42_pop_bits;
	wire _stealNW_TQ_io_connPE_43_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_43_pop_bits;
	wire _stealNW_TQ_io_connPE_44_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_44_pop_bits;
	wire _stealNW_TQ_io_connPE_45_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_45_pop_bits;
	wire _stealNW_TQ_io_connPE_46_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_46_pop_bits;
	wire _stealNW_TQ_io_connPE_47_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_47_pop_bits;
	wire _stealNW_TQ_io_connPE_48_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_48_pop_bits;
	wire _stealNW_TQ_io_connPE_49_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_49_pop_bits;
	wire _stealNW_TQ_io_connPE_50_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_50_pop_bits;
	wire _stealNW_TQ_io_connPE_51_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_51_pop_bits;
	wire _stealNW_TQ_io_connPE_52_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_52_pop_bits;
	wire _stealNW_TQ_io_connPE_53_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_53_pop_bits;
	wire _stealNW_TQ_io_connPE_54_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_54_pop_bits;
	wire _stealNW_TQ_io_connPE_55_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_55_pop_bits;
	wire _stealNW_TQ_io_connPE_56_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_56_pop_bits;
	wire _stealNW_TQ_io_connPE_57_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_57_pop_bits;
	wire _stealNW_TQ_io_connPE_58_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_58_pop_bits;
	wire _stealNW_TQ_io_connPE_59_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_59_pop_bits;
	wire _stealNW_TQ_io_connPE_60_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_60_pop_bits;
	wire _stealNW_TQ_io_connPE_61_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_61_pop_bits;
	wire _stealNW_TQ_io_connPE_62_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_62_pop_bits;
	wire _stealNW_TQ_io_connPE_63_pop_valid;
	wire [255:0] _stealNW_TQ_io_connPE_63_pop_bits;
	wire _stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready;
	wire _stealNW_TQ_io_connVSS_0_data_availableTask_valid;
	wire [255:0] _stealNW_TQ_io_connVSS_0_data_availableTask_bits;
	wire _stealNW_TQ_io_connVSS_0_data_qOutTask_ready;
	wire _stealNW_TQ_io_connVSS_1_ctrl_serveStealReq_ready;
	wire _stealNW_TQ_io_connVSS_1_data_availableTask_valid;
	wire [255:0] _stealNW_TQ_io_connVSS_1_data_availableTask_bits;
	wire _stealNW_TQ_io_connVSS_1_data_qOutTask_ready;
	wire _stealNW_TQ_io_ntwDataUnitOccupancyVSS_0;
	wire _stealNW_TQ_io_ntwDataUnitOccupancyVSS_1;
	SchedulerLocalNetwork_1 stealNW_TQ(
		.clock(clock),
		.reset(reset),
		.io_connPE_0_pop_ready(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_connPE_0_pop_valid(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_connPE_0_pop_bits(_stealNW_TQ_io_connPE_0_pop_bits),
		.io_connPE_1_pop_ready(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_connPE_1_pop_valid(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_connPE_1_pop_bits(_stealNW_TQ_io_connPE_1_pop_bits),
		.io_connPE_2_pop_ready(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_connPE_2_pop_valid(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_connPE_2_pop_bits(_stealNW_TQ_io_connPE_2_pop_bits),
		.io_connPE_3_pop_ready(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_connPE_3_pop_valid(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_connPE_3_pop_bits(_stealNW_TQ_io_connPE_3_pop_bits),
		.io_connPE_4_pop_ready(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_connPE_4_pop_valid(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_connPE_4_pop_bits(_stealNW_TQ_io_connPE_4_pop_bits),
		.io_connPE_5_pop_ready(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_connPE_5_pop_valid(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_connPE_5_pop_bits(_stealNW_TQ_io_connPE_5_pop_bits),
		.io_connPE_6_pop_ready(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_connPE_6_pop_valid(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_connPE_6_pop_bits(_stealNW_TQ_io_connPE_6_pop_bits),
		.io_connPE_7_pop_ready(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_connPE_7_pop_valid(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_connPE_7_pop_bits(_stealNW_TQ_io_connPE_7_pop_bits),
		.io_connPE_8_pop_ready(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_connPE_8_pop_valid(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_connPE_8_pop_bits(_stealNW_TQ_io_connPE_8_pop_bits),
		.io_connPE_9_pop_ready(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_connPE_9_pop_valid(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_connPE_9_pop_bits(_stealNW_TQ_io_connPE_9_pop_bits),
		.io_connPE_10_pop_ready(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_connPE_10_pop_valid(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_connPE_10_pop_bits(_stealNW_TQ_io_connPE_10_pop_bits),
		.io_connPE_11_pop_ready(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_connPE_11_pop_valid(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_connPE_11_pop_bits(_stealNW_TQ_io_connPE_11_pop_bits),
		.io_connPE_12_pop_ready(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_connPE_12_pop_valid(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_connPE_12_pop_bits(_stealNW_TQ_io_connPE_12_pop_bits),
		.io_connPE_13_pop_ready(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_connPE_13_pop_valid(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_connPE_13_pop_bits(_stealNW_TQ_io_connPE_13_pop_bits),
		.io_connPE_14_pop_ready(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_connPE_14_pop_valid(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_connPE_14_pop_bits(_stealNW_TQ_io_connPE_14_pop_bits),
		.io_connPE_15_pop_ready(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_connPE_15_pop_valid(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_connPE_15_pop_bits(_stealNW_TQ_io_connPE_15_pop_bits),
		.io_connPE_16_pop_ready(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_connPE_16_pop_valid(_stealNW_TQ_io_connPE_16_pop_valid),
		.io_connPE_16_pop_bits(_stealNW_TQ_io_connPE_16_pop_bits),
		.io_connPE_17_pop_ready(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_connPE_17_pop_valid(_stealNW_TQ_io_connPE_17_pop_valid),
		.io_connPE_17_pop_bits(_stealNW_TQ_io_connPE_17_pop_bits),
		.io_connPE_18_pop_ready(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_connPE_18_pop_valid(_stealNW_TQ_io_connPE_18_pop_valid),
		.io_connPE_18_pop_bits(_stealNW_TQ_io_connPE_18_pop_bits),
		.io_connPE_19_pop_ready(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_connPE_19_pop_valid(_stealNW_TQ_io_connPE_19_pop_valid),
		.io_connPE_19_pop_bits(_stealNW_TQ_io_connPE_19_pop_bits),
		.io_connPE_20_pop_ready(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_connPE_20_pop_valid(_stealNW_TQ_io_connPE_20_pop_valid),
		.io_connPE_20_pop_bits(_stealNW_TQ_io_connPE_20_pop_bits),
		.io_connPE_21_pop_ready(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_connPE_21_pop_valid(_stealNW_TQ_io_connPE_21_pop_valid),
		.io_connPE_21_pop_bits(_stealNW_TQ_io_connPE_21_pop_bits),
		.io_connPE_22_pop_ready(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_connPE_22_pop_valid(_stealNW_TQ_io_connPE_22_pop_valid),
		.io_connPE_22_pop_bits(_stealNW_TQ_io_connPE_22_pop_bits),
		.io_connPE_23_pop_ready(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_connPE_23_pop_valid(_stealNW_TQ_io_connPE_23_pop_valid),
		.io_connPE_23_pop_bits(_stealNW_TQ_io_connPE_23_pop_bits),
		.io_connPE_24_pop_ready(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_connPE_24_pop_valid(_stealNW_TQ_io_connPE_24_pop_valid),
		.io_connPE_24_pop_bits(_stealNW_TQ_io_connPE_24_pop_bits),
		.io_connPE_25_pop_ready(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_connPE_25_pop_valid(_stealNW_TQ_io_connPE_25_pop_valid),
		.io_connPE_25_pop_bits(_stealNW_TQ_io_connPE_25_pop_bits),
		.io_connPE_26_pop_ready(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_connPE_26_pop_valid(_stealNW_TQ_io_connPE_26_pop_valid),
		.io_connPE_26_pop_bits(_stealNW_TQ_io_connPE_26_pop_bits),
		.io_connPE_27_pop_ready(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_connPE_27_pop_valid(_stealNW_TQ_io_connPE_27_pop_valid),
		.io_connPE_27_pop_bits(_stealNW_TQ_io_connPE_27_pop_bits),
		.io_connPE_28_pop_ready(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_connPE_28_pop_valid(_stealNW_TQ_io_connPE_28_pop_valid),
		.io_connPE_28_pop_bits(_stealNW_TQ_io_connPE_28_pop_bits),
		.io_connPE_29_pop_ready(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_connPE_29_pop_valid(_stealNW_TQ_io_connPE_29_pop_valid),
		.io_connPE_29_pop_bits(_stealNW_TQ_io_connPE_29_pop_bits),
		.io_connPE_30_pop_ready(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_connPE_30_pop_valid(_stealNW_TQ_io_connPE_30_pop_valid),
		.io_connPE_30_pop_bits(_stealNW_TQ_io_connPE_30_pop_bits),
		.io_connPE_31_pop_ready(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_connPE_31_pop_valid(_stealNW_TQ_io_connPE_31_pop_valid),
		.io_connPE_31_pop_bits(_stealNW_TQ_io_connPE_31_pop_bits),
		.io_connPE_32_pop_ready(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_connPE_32_pop_valid(_stealNW_TQ_io_connPE_32_pop_valid),
		.io_connPE_32_pop_bits(_stealNW_TQ_io_connPE_32_pop_bits),
		.io_connPE_33_pop_ready(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_connPE_33_pop_valid(_stealNW_TQ_io_connPE_33_pop_valid),
		.io_connPE_33_pop_bits(_stealNW_TQ_io_connPE_33_pop_bits),
		.io_connPE_34_pop_ready(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_connPE_34_pop_valid(_stealNW_TQ_io_connPE_34_pop_valid),
		.io_connPE_34_pop_bits(_stealNW_TQ_io_connPE_34_pop_bits),
		.io_connPE_35_pop_ready(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_connPE_35_pop_valid(_stealNW_TQ_io_connPE_35_pop_valid),
		.io_connPE_35_pop_bits(_stealNW_TQ_io_connPE_35_pop_bits),
		.io_connPE_36_pop_ready(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_connPE_36_pop_valid(_stealNW_TQ_io_connPE_36_pop_valid),
		.io_connPE_36_pop_bits(_stealNW_TQ_io_connPE_36_pop_bits),
		.io_connPE_37_pop_ready(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_connPE_37_pop_valid(_stealNW_TQ_io_connPE_37_pop_valid),
		.io_connPE_37_pop_bits(_stealNW_TQ_io_connPE_37_pop_bits),
		.io_connPE_38_pop_ready(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_connPE_38_pop_valid(_stealNW_TQ_io_connPE_38_pop_valid),
		.io_connPE_38_pop_bits(_stealNW_TQ_io_connPE_38_pop_bits),
		.io_connPE_39_pop_ready(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_connPE_39_pop_valid(_stealNW_TQ_io_connPE_39_pop_valid),
		.io_connPE_39_pop_bits(_stealNW_TQ_io_connPE_39_pop_bits),
		.io_connPE_40_pop_ready(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_connPE_40_pop_valid(_stealNW_TQ_io_connPE_40_pop_valid),
		.io_connPE_40_pop_bits(_stealNW_TQ_io_connPE_40_pop_bits),
		.io_connPE_41_pop_ready(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_connPE_41_pop_valid(_stealNW_TQ_io_connPE_41_pop_valid),
		.io_connPE_41_pop_bits(_stealNW_TQ_io_connPE_41_pop_bits),
		.io_connPE_42_pop_ready(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_connPE_42_pop_valid(_stealNW_TQ_io_connPE_42_pop_valid),
		.io_connPE_42_pop_bits(_stealNW_TQ_io_connPE_42_pop_bits),
		.io_connPE_43_pop_ready(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_connPE_43_pop_valid(_stealNW_TQ_io_connPE_43_pop_valid),
		.io_connPE_43_pop_bits(_stealNW_TQ_io_connPE_43_pop_bits),
		.io_connPE_44_pop_ready(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_connPE_44_pop_valid(_stealNW_TQ_io_connPE_44_pop_valid),
		.io_connPE_44_pop_bits(_stealNW_TQ_io_connPE_44_pop_bits),
		.io_connPE_45_pop_ready(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_connPE_45_pop_valid(_stealNW_TQ_io_connPE_45_pop_valid),
		.io_connPE_45_pop_bits(_stealNW_TQ_io_connPE_45_pop_bits),
		.io_connPE_46_pop_ready(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_connPE_46_pop_valid(_stealNW_TQ_io_connPE_46_pop_valid),
		.io_connPE_46_pop_bits(_stealNW_TQ_io_connPE_46_pop_bits),
		.io_connPE_47_pop_ready(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_connPE_47_pop_valid(_stealNW_TQ_io_connPE_47_pop_valid),
		.io_connPE_47_pop_bits(_stealNW_TQ_io_connPE_47_pop_bits),
		.io_connPE_48_pop_ready(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_connPE_48_pop_valid(_stealNW_TQ_io_connPE_48_pop_valid),
		.io_connPE_48_pop_bits(_stealNW_TQ_io_connPE_48_pop_bits),
		.io_connPE_49_pop_ready(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_connPE_49_pop_valid(_stealNW_TQ_io_connPE_49_pop_valid),
		.io_connPE_49_pop_bits(_stealNW_TQ_io_connPE_49_pop_bits),
		.io_connPE_50_pop_ready(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_connPE_50_pop_valid(_stealNW_TQ_io_connPE_50_pop_valid),
		.io_connPE_50_pop_bits(_stealNW_TQ_io_connPE_50_pop_bits),
		.io_connPE_51_pop_ready(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_connPE_51_pop_valid(_stealNW_TQ_io_connPE_51_pop_valid),
		.io_connPE_51_pop_bits(_stealNW_TQ_io_connPE_51_pop_bits),
		.io_connPE_52_pop_ready(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_connPE_52_pop_valid(_stealNW_TQ_io_connPE_52_pop_valid),
		.io_connPE_52_pop_bits(_stealNW_TQ_io_connPE_52_pop_bits),
		.io_connPE_53_pop_ready(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_connPE_53_pop_valid(_stealNW_TQ_io_connPE_53_pop_valid),
		.io_connPE_53_pop_bits(_stealNW_TQ_io_connPE_53_pop_bits),
		.io_connPE_54_pop_ready(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_connPE_54_pop_valid(_stealNW_TQ_io_connPE_54_pop_valid),
		.io_connPE_54_pop_bits(_stealNW_TQ_io_connPE_54_pop_bits),
		.io_connPE_55_pop_ready(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_connPE_55_pop_valid(_stealNW_TQ_io_connPE_55_pop_valid),
		.io_connPE_55_pop_bits(_stealNW_TQ_io_connPE_55_pop_bits),
		.io_connPE_56_pop_ready(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_connPE_56_pop_valid(_stealNW_TQ_io_connPE_56_pop_valid),
		.io_connPE_56_pop_bits(_stealNW_TQ_io_connPE_56_pop_bits),
		.io_connPE_57_pop_ready(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_connPE_57_pop_valid(_stealNW_TQ_io_connPE_57_pop_valid),
		.io_connPE_57_pop_bits(_stealNW_TQ_io_connPE_57_pop_bits),
		.io_connPE_58_pop_ready(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_connPE_58_pop_valid(_stealNW_TQ_io_connPE_58_pop_valid),
		.io_connPE_58_pop_bits(_stealNW_TQ_io_connPE_58_pop_bits),
		.io_connPE_59_pop_ready(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_connPE_59_pop_valid(_stealNW_TQ_io_connPE_59_pop_valid),
		.io_connPE_59_pop_bits(_stealNW_TQ_io_connPE_59_pop_bits),
		.io_connPE_60_pop_ready(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_connPE_60_pop_valid(_stealNW_TQ_io_connPE_60_pop_valid),
		.io_connPE_60_pop_bits(_stealNW_TQ_io_connPE_60_pop_bits),
		.io_connPE_61_pop_ready(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_connPE_61_pop_valid(_stealNW_TQ_io_connPE_61_pop_valid),
		.io_connPE_61_pop_bits(_stealNW_TQ_io_connPE_61_pop_bits),
		.io_connPE_62_pop_ready(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_connPE_62_pop_valid(_stealNW_TQ_io_connPE_62_pop_valid),
		.io_connPE_62_pop_bits(_stealNW_TQ_io_connPE_62_pop_bits),
		.io_connPE_63_pop_ready(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_connPE_63_pop_valid(_stealNW_TQ_io_connPE_63_pop_valid),
		.io_connPE_63_pop_bits(_stealNW_TQ_io_connPE_63_pop_bits),
		.io_connVSS_0_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connVSS_0_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connVSS_0_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connVSS_0_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connVSS_0_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connVSS_0_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connVSS_0_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connVSS_0_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connVSS_1_ctrl_serveStealReq_valid(_virtualStealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connVSS_1_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_1_ctrl_serveStealReq_ready),
		.io_connVSS_1_data_availableTask_ready(_virtualStealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connVSS_1_data_availableTask_valid(_stealNW_TQ_io_connVSS_1_data_availableTask_valid),
		.io_connVSS_1_data_availableTask_bits(_stealNW_TQ_io_connVSS_1_data_availableTask_bits),
		.io_connVSS_1_data_qOutTask_ready(_stealNW_TQ_io_connVSS_1_data_qOutTask_ready),
		.io_connVSS_1_data_qOutTask_valid(_virtualStealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connVSS_1_data_qOutTask_bits(_virtualStealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connVAS_0_ctrl_serveStealReq_valid(connArgumentNotifier_0_ctrl_serveStealReq_valid),
		.io_connVAS_0_ctrl_serveStealReq_ready(connArgumentNotifier_0_ctrl_serveStealReq_ready),
		.io_connVAS_0_data_qOutTask_ready(connArgumentNotifier_0_data_qOutTask_ready),
		.io_connVAS_0_data_qOutTask_valid(connArgumentNotifier_0_data_qOutTask_valid),
		.io_connVAS_0_data_qOutTask_bits(connArgumentNotifier_0_data_qOutTask_bits),
		.io_connVAS_1_ctrl_serveStealReq_valid(connArgumentNotifier_1_ctrl_serveStealReq_valid),
		.io_connVAS_1_ctrl_serveStealReq_ready(connArgumentNotifier_1_ctrl_serveStealReq_ready),
		.io_connVAS_1_data_qOutTask_ready(connArgumentNotifier_1_data_qOutTask_ready),
		.io_connVAS_1_data_qOutTask_valid(connArgumentNotifier_1_data_qOutTask_valid),
		.io_connVAS_1_data_qOutTask_bits(connArgumentNotifier_1_data_qOutTask_bits),
		.io_connVAS_2_ctrl_serveStealReq_valid(connArgumentNotifier_2_ctrl_serveStealReq_valid),
		.io_connVAS_2_ctrl_serveStealReq_ready(connArgumentNotifier_2_ctrl_serveStealReq_ready),
		.io_connVAS_2_data_qOutTask_ready(connArgumentNotifier_2_data_qOutTask_ready),
		.io_connVAS_2_data_qOutTask_valid(connArgumentNotifier_2_data_qOutTask_valid),
		.io_connVAS_2_data_qOutTask_bits(connArgumentNotifier_2_data_qOutTask_bits),
		.io_connVAS_3_ctrl_serveStealReq_valid(connArgumentNotifier_3_ctrl_serveStealReq_valid),
		.io_connVAS_3_ctrl_serveStealReq_ready(connArgumentNotifier_3_ctrl_serveStealReq_ready),
		.io_connVAS_3_data_qOutTask_ready(connArgumentNotifier_3_data_qOutTask_ready),
		.io_connVAS_3_data_qOutTask_valid(connArgumentNotifier_3_data_qOutTask_valid),
		.io_connVAS_3_data_qOutTask_bits(connArgumentNotifier_3_data_qOutTask_bits),
		.io_connVAS_4_ctrl_serveStealReq_valid(connArgumentNotifier_4_ctrl_serveStealReq_valid),
		.io_connVAS_4_ctrl_serveStealReq_ready(connArgumentNotifier_4_ctrl_serveStealReq_ready),
		.io_connVAS_4_data_qOutTask_ready(connArgumentNotifier_4_data_qOutTask_ready),
		.io_connVAS_4_data_qOutTask_valid(connArgumentNotifier_4_data_qOutTask_valid),
		.io_connVAS_4_data_qOutTask_bits(connArgumentNotifier_4_data_qOutTask_bits),
		.io_connVAS_5_ctrl_serveStealReq_valid(connArgumentNotifier_5_ctrl_serveStealReq_valid),
		.io_connVAS_5_ctrl_serveStealReq_ready(connArgumentNotifier_5_ctrl_serveStealReq_ready),
		.io_connVAS_5_data_qOutTask_ready(connArgumentNotifier_5_data_qOutTask_ready),
		.io_connVAS_5_data_qOutTask_valid(connArgumentNotifier_5_data_qOutTask_valid),
		.io_connVAS_5_data_qOutTask_bits(connArgumentNotifier_5_data_qOutTask_bits),
		.io_connVAS_6_ctrl_serveStealReq_valid(connArgumentNotifier_6_ctrl_serveStealReq_valid),
		.io_connVAS_6_ctrl_serveStealReq_ready(connArgumentNotifier_6_ctrl_serveStealReq_ready),
		.io_connVAS_6_data_qOutTask_ready(connArgumentNotifier_6_data_qOutTask_ready),
		.io_connVAS_6_data_qOutTask_valid(connArgumentNotifier_6_data_qOutTask_valid),
		.io_connVAS_6_data_qOutTask_bits(connArgumentNotifier_6_data_qOutTask_bits),
		.io_connVAS_7_ctrl_serveStealReq_valid(connArgumentNotifier_7_ctrl_serveStealReq_valid),
		.io_connVAS_7_ctrl_serveStealReq_ready(connArgumentNotifier_7_ctrl_serveStealReq_ready),
		.io_connVAS_7_data_qOutTask_ready(connArgumentNotifier_7_data_qOutTask_ready),
		.io_connVAS_7_data_qOutTask_valid(connArgumentNotifier_7_data_qOutTask_valid),
		.io_connVAS_7_data_qOutTask_bits(connArgumentNotifier_7_data_qOutTask_bits),
		.io_connVAS_8_ctrl_serveStealReq_valid(connArgumentNotifier_8_ctrl_serveStealReq_valid),
		.io_connVAS_8_ctrl_serveStealReq_ready(connArgumentNotifier_8_ctrl_serveStealReq_ready),
		.io_connVAS_8_data_qOutTask_ready(connArgumentNotifier_8_data_qOutTask_ready),
		.io_connVAS_8_data_qOutTask_valid(connArgumentNotifier_8_data_qOutTask_valid),
		.io_connVAS_8_data_qOutTask_bits(connArgumentNotifier_8_data_qOutTask_bits),
		.io_connVAS_9_ctrl_serveStealReq_valid(connArgumentNotifier_9_ctrl_serveStealReq_valid),
		.io_connVAS_9_ctrl_serveStealReq_ready(connArgumentNotifier_9_ctrl_serveStealReq_ready),
		.io_connVAS_9_data_qOutTask_ready(connArgumentNotifier_9_data_qOutTask_ready),
		.io_connVAS_9_data_qOutTask_valid(connArgumentNotifier_9_data_qOutTask_valid),
		.io_connVAS_9_data_qOutTask_bits(connArgumentNotifier_9_data_qOutTask_bits),
		.io_connVAS_10_ctrl_serveStealReq_valid(connArgumentNotifier_10_ctrl_serveStealReq_valid),
		.io_connVAS_10_ctrl_serveStealReq_ready(connArgumentNotifier_10_ctrl_serveStealReq_ready),
		.io_connVAS_10_data_qOutTask_ready(connArgumentNotifier_10_data_qOutTask_ready),
		.io_connVAS_10_data_qOutTask_valid(connArgumentNotifier_10_data_qOutTask_valid),
		.io_connVAS_10_data_qOutTask_bits(connArgumentNotifier_10_data_qOutTask_bits),
		.io_connVAS_11_ctrl_serveStealReq_valid(connArgumentNotifier_11_ctrl_serveStealReq_valid),
		.io_connVAS_11_ctrl_serveStealReq_ready(connArgumentNotifier_11_ctrl_serveStealReq_ready),
		.io_connVAS_11_data_qOutTask_ready(connArgumentNotifier_11_data_qOutTask_ready),
		.io_connVAS_11_data_qOutTask_valid(connArgumentNotifier_11_data_qOutTask_valid),
		.io_connVAS_11_data_qOutTask_bits(connArgumentNotifier_11_data_qOutTask_bits),
		.io_connVAS_12_ctrl_serveStealReq_valid(connArgumentNotifier_12_ctrl_serveStealReq_valid),
		.io_connVAS_12_ctrl_serveStealReq_ready(connArgumentNotifier_12_ctrl_serveStealReq_ready),
		.io_connVAS_12_data_qOutTask_ready(connArgumentNotifier_12_data_qOutTask_ready),
		.io_connVAS_12_data_qOutTask_valid(connArgumentNotifier_12_data_qOutTask_valid),
		.io_connVAS_12_data_qOutTask_bits(connArgumentNotifier_12_data_qOutTask_bits),
		.io_connVAS_13_ctrl_serveStealReq_valid(connArgumentNotifier_13_ctrl_serveStealReq_valid),
		.io_connVAS_13_ctrl_serveStealReq_ready(connArgumentNotifier_13_ctrl_serveStealReq_ready),
		.io_connVAS_13_data_qOutTask_ready(connArgumentNotifier_13_data_qOutTask_ready),
		.io_connVAS_13_data_qOutTask_valid(connArgumentNotifier_13_data_qOutTask_valid),
		.io_connVAS_13_data_qOutTask_bits(connArgumentNotifier_13_data_qOutTask_bits),
		.io_connVAS_14_ctrl_serveStealReq_valid(connArgumentNotifier_14_ctrl_serveStealReq_valid),
		.io_connVAS_14_ctrl_serveStealReq_ready(connArgumentNotifier_14_ctrl_serveStealReq_ready),
		.io_connVAS_14_data_qOutTask_ready(connArgumentNotifier_14_data_qOutTask_ready),
		.io_connVAS_14_data_qOutTask_valid(connArgumentNotifier_14_data_qOutTask_valid),
		.io_connVAS_14_data_qOutTask_bits(connArgumentNotifier_14_data_qOutTask_bits),
		.io_connVAS_15_ctrl_serveStealReq_valid(connArgumentNotifier_15_ctrl_serveStealReq_valid),
		.io_connVAS_15_ctrl_serveStealReq_ready(connArgumentNotifier_15_ctrl_serveStealReq_ready),
		.io_connVAS_15_data_qOutTask_ready(connArgumentNotifier_15_data_qOutTask_ready),
		.io_connVAS_15_data_qOutTask_valid(connArgumentNotifier_15_data_qOutTask_valid),
		.io_connVAS_15_data_qOutTask_bits(connArgumentNotifier_15_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0),
		.io_ntwDataUnitOccupancyVSS_1(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_1)
	);
	SchedulerServer_2 virtualStealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connNetwork_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vss_0_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vss_0_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vss_0_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vss_0_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vss_0_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vss_0_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vss_0_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vss_0_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vss_0_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vss_0_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vss_0_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vss_0_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vss_0_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vss_0_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vss_0_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vss_0_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vss_0_b_bits_resp),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_read_burst_len(_virtualStealServers_0_io_read_burst_len),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_write_burst_len(_virtualStealServers_0_io_write_burst_len),
		.io_write_last(_virtualStealServers_0_io_write_last),
		.io_ntwDataUnitOccupancy(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerServer_2 virtualStealServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_virtualStealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_1_ctrl_serveStealReq_ready),
		.io_connNetwork_data_availableTask_ready(_virtualStealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNW_TQ_io_connVSS_1_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNW_TQ_io_connVSS_1_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNW_TQ_io_connVSS_1_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_virtualStealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_virtualStealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vss_1_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vss_1_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vss_1_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vss_1_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vss_1_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vss_1_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vss_1_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vss_1_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vss_1_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vss_1_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vss_1_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vss_1_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vss_1_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vss_1_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vss_1_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vss_1_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vss_1_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vss_1_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vss_1_b_bits_resp),
		.io_read_address_ready(_vssRvm_1_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_1_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_1_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_1_io_read_data_ready),
		.io_read_data_valid(_vssRvm_1_io_read_data_valid),
		.io_read_data_bits(_vssRvm_1_io_read_data_bits),
		.io_read_burst_len(_virtualStealServers_1_io_read_burst_len),
		.io_write_address_ready(_vssRvm_1_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_1_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_1_io_write_address_bits),
		.io_write_data_ready(_vssRvm_1_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_1_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_1_io_write_data_bits),
		.io_write_burst_len(_virtualStealServers_1_io_write_burst_len),
		.io_write_last(_virtualStealServers_1_io_write_last),
		.io_ntwDataUnitOccupancy(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_1)
	);
	RVtoAXIBridge_2 vssRvm_0(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_writeBurst_len(_virtualStealServers_0_io_write_burst_len),
		.io_writeBurst_last(_virtualStealServers_0_io_write_last),
		.io_readBurst_len(_virtualStealServers_0_io_read_burst_len),
		.axi_ar_ready(_module_s_axi_ar_ready),
		.axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.axi_r_ready(_vssRvm_0_axi_r_ready),
		.axi_r_valid(_module_s_axi_r_valid),
		.axi_r_bits_data(_module_s_axi_r_bits_data),
		.axi_aw_ready(_module_s_axi_aw_ready),
		.axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.axi_aw_bits_len(_vssRvm_0_axi_aw_bits_len),
		.axi_w_ready(_module_s_axi_w_ready),
		.axi_w_valid(_vssRvm_0_axi_w_valid),
		.axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.axi_b_valid(_module_s_axi_b_valid)
	);
	RVtoAXIBridge_2 vssRvm_1(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_vssRvm_1_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_1_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_1_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_1_io_read_data_ready),
		.io_read_data_valid(_vssRvm_1_io_read_data_valid),
		.io_read_data_bits(_vssRvm_1_io_read_data_bits),
		.io_write_address_ready(_vssRvm_1_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_1_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_1_io_write_address_bits),
		.io_write_data_ready(_vssRvm_1_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_1_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_1_io_write_data_bits),
		.io_writeBurst_len(_virtualStealServers_1_io_write_burst_len),
		.io_writeBurst_last(_virtualStealServers_1_io_write_last),
		.io_readBurst_len(_virtualStealServers_1_io_read_burst_len),
		.axi_ar_ready(_module_1_s_axi_ar_ready),
		.axi_ar_valid(_vssRvm_1_axi_ar_valid),
		.axi_ar_bits_addr(_vssRvm_1_axi_ar_bits_addr),
		.axi_ar_bits_len(_vssRvm_1_axi_ar_bits_len),
		.axi_r_ready(_vssRvm_1_axi_r_ready),
		.axi_r_valid(_module_1_s_axi_r_valid),
		.axi_r_bits_data(_module_1_s_axi_r_bits_data),
		.axi_aw_ready(_module_1_s_axi_aw_ready),
		.axi_aw_valid(_vssRvm_1_axi_aw_valid),
		.axi_aw_bits_addr(_vssRvm_1_axi_aw_bits_addr),
		.axi_aw_bits_len(_vssRvm_1_axi_aw_bits_len),
		.axi_w_ready(_module_1_s_axi_w_ready),
		.axi_w_valid(_vssRvm_1_axi_w_valid),
		.axi_w_bits_data(_vssRvm_1_axi_w_bits_data),
		.axi_w_bits_last(_vssRvm_1_axi_w_bits_last),
		.axi_b_valid(_module_1_s_axi_b_valid)
	);
	axi4FullMux_1 mux(
		.clock(clock),
		.reset(reset),
		.s_axi_0_ar_ready(_mux_s_axi_0_ar_ready),
		.s_axi_0_ar_valid(_module_m_axi_ar_valid),
		.s_axi_0_ar_bits_addr(_module_m_axi_ar_bits_addr),
		.s_axi_0_ar_bits_len(_module_m_axi_ar_bits_len),
		.s_axi_0_ar_bits_size(_module_m_axi_ar_bits_size),
		.s_axi_0_ar_bits_burst(_module_m_axi_ar_bits_burst),
		.s_axi_0_ar_bits_lock(_module_m_axi_ar_bits_lock),
		.s_axi_0_ar_bits_cache(_module_m_axi_ar_bits_cache),
		.s_axi_0_ar_bits_prot(_module_m_axi_ar_bits_prot),
		.s_axi_0_ar_bits_qos(_module_m_axi_ar_bits_qos),
		.s_axi_0_ar_bits_region(_module_m_axi_ar_bits_region),
		.s_axi_0_r_ready(_module_m_axi_r_ready),
		.s_axi_0_r_valid(_mux_s_axi_0_r_valid),
		.s_axi_0_r_bits_data(_mux_s_axi_0_r_bits_data),
		.s_axi_0_aw_ready(_mux_s_axi_0_aw_ready),
		.s_axi_0_aw_valid(_module_m_axi_aw_valid),
		.s_axi_0_aw_bits_addr(_module_m_axi_aw_bits_addr),
		.s_axi_0_aw_bits_len(_module_m_axi_aw_bits_len),
		.s_axi_0_aw_bits_size(_module_m_axi_aw_bits_size),
		.s_axi_0_aw_bits_burst(_module_m_axi_aw_bits_burst),
		.s_axi_0_aw_bits_lock(_module_m_axi_aw_bits_lock),
		.s_axi_0_aw_bits_cache(_module_m_axi_aw_bits_cache),
		.s_axi_0_aw_bits_prot(_module_m_axi_aw_bits_prot),
		.s_axi_0_aw_bits_qos(_module_m_axi_aw_bits_qos),
		.s_axi_0_aw_bits_region(_module_m_axi_aw_bits_region),
		.s_axi_0_w_ready(_mux_s_axi_0_w_ready),
		.s_axi_0_w_valid(_module_m_axi_w_valid),
		.s_axi_0_w_bits_data(_module_m_axi_w_bits_data),
		.s_axi_0_w_bits_last(_module_m_axi_w_bits_last),
		.s_axi_0_b_valid(_mux_s_axi_0_b_valid),
		.s_axi_1_ar_ready(_mux_s_axi_1_ar_ready),
		.s_axi_1_ar_valid(_module_1_m_axi_ar_valid),
		.s_axi_1_ar_bits_addr(_module_1_m_axi_ar_bits_addr),
		.s_axi_1_ar_bits_len(_module_1_m_axi_ar_bits_len),
		.s_axi_1_ar_bits_size(_module_1_m_axi_ar_bits_size),
		.s_axi_1_ar_bits_burst(_module_1_m_axi_ar_bits_burst),
		.s_axi_1_ar_bits_lock(_module_1_m_axi_ar_bits_lock),
		.s_axi_1_ar_bits_cache(_module_1_m_axi_ar_bits_cache),
		.s_axi_1_ar_bits_prot(_module_1_m_axi_ar_bits_prot),
		.s_axi_1_ar_bits_qos(_module_1_m_axi_ar_bits_qos),
		.s_axi_1_ar_bits_region(_module_1_m_axi_ar_bits_region),
		.s_axi_1_r_ready(_module_1_m_axi_r_ready),
		.s_axi_1_r_valid(_mux_s_axi_1_r_valid),
		.s_axi_1_r_bits_data(_mux_s_axi_1_r_bits_data),
		.s_axi_1_aw_ready(_mux_s_axi_1_aw_ready),
		.s_axi_1_aw_valid(_module_1_m_axi_aw_valid),
		.s_axi_1_aw_bits_addr(_module_1_m_axi_aw_bits_addr),
		.s_axi_1_aw_bits_len(_module_1_m_axi_aw_bits_len),
		.s_axi_1_aw_bits_size(_module_1_m_axi_aw_bits_size),
		.s_axi_1_aw_bits_burst(_module_1_m_axi_aw_bits_burst),
		.s_axi_1_aw_bits_lock(_module_1_m_axi_aw_bits_lock),
		.s_axi_1_aw_bits_cache(_module_1_m_axi_aw_bits_cache),
		.s_axi_1_aw_bits_prot(_module_1_m_axi_aw_bits_prot),
		.s_axi_1_aw_bits_qos(_module_1_m_axi_aw_bits_qos),
		.s_axi_1_aw_bits_region(_module_1_m_axi_aw_bits_region),
		.s_axi_1_w_ready(_mux_s_axi_1_w_ready),
		.s_axi_1_w_valid(_module_1_m_axi_w_valid),
		.s_axi_1_w_bits_data(_module_1_m_axi_w_bits_data),
		.s_axi_1_w_bits_last(_module_1_m_axi_w_bits_last),
		.s_axi_1_b_valid(_mux_s_axi_1_b_valid),
		.m_axi_ar_ready(io_internal_vss_axi_full_0_ar_ready),
		.m_axi_ar_valid(io_internal_vss_axi_full_0_ar_valid),
		.m_axi_ar_bits_id(io_internal_vss_axi_full_0_ar_bits_id),
		.m_axi_ar_bits_addr(io_internal_vss_axi_full_0_ar_bits_addr),
		.m_axi_ar_bits_len(io_internal_vss_axi_full_0_ar_bits_len),
		.m_axi_ar_bits_size(io_internal_vss_axi_full_0_ar_bits_size),
		.m_axi_ar_bits_burst(io_internal_vss_axi_full_0_ar_bits_burst),
		.m_axi_ar_bits_lock(io_internal_vss_axi_full_0_ar_bits_lock),
		.m_axi_ar_bits_cache(io_internal_vss_axi_full_0_ar_bits_cache),
		.m_axi_ar_bits_prot(io_internal_vss_axi_full_0_ar_bits_prot),
		.m_axi_ar_bits_qos(io_internal_vss_axi_full_0_ar_bits_qos),
		.m_axi_ar_bits_region(io_internal_vss_axi_full_0_ar_bits_region),
		.m_axi_r_ready(io_internal_vss_axi_full_0_r_ready),
		.m_axi_r_valid(io_internal_vss_axi_full_0_r_valid),
		.m_axi_r_bits_id(io_internal_vss_axi_full_0_r_bits_id),
		.m_axi_r_bits_data(io_internal_vss_axi_full_0_r_bits_data),
		.m_axi_r_bits_resp(io_internal_vss_axi_full_0_r_bits_resp),
		.m_axi_r_bits_last(io_internal_vss_axi_full_0_r_bits_last),
		.m_axi_aw_ready(io_internal_vss_axi_full_0_aw_ready),
		.m_axi_aw_valid(io_internal_vss_axi_full_0_aw_valid),
		.m_axi_aw_bits_id(io_internal_vss_axi_full_0_aw_bits_id),
		.m_axi_aw_bits_addr(io_internal_vss_axi_full_0_aw_bits_addr),
		.m_axi_aw_bits_len(io_internal_vss_axi_full_0_aw_bits_len),
		.m_axi_aw_bits_size(io_internal_vss_axi_full_0_aw_bits_size),
		.m_axi_aw_bits_burst(io_internal_vss_axi_full_0_aw_bits_burst),
		.m_axi_aw_bits_lock(io_internal_vss_axi_full_0_aw_bits_lock),
		.m_axi_aw_bits_cache(io_internal_vss_axi_full_0_aw_bits_cache),
		.m_axi_aw_bits_prot(io_internal_vss_axi_full_0_aw_bits_prot),
		.m_axi_aw_bits_qos(io_internal_vss_axi_full_0_aw_bits_qos),
		.m_axi_aw_bits_region(io_internal_vss_axi_full_0_aw_bits_region),
		.m_axi_w_ready(io_internal_vss_axi_full_0_w_ready),
		.m_axi_w_valid(io_internal_vss_axi_full_0_w_valid),
		.m_axi_w_bits_data(io_internal_vss_axi_full_0_w_bits_data),
		.m_axi_w_bits_strb(io_internal_vss_axi_full_0_w_bits_strb),
		.m_axi_w_bits_last(io_internal_vss_axi_full_0_w_bits_last),
		.m_axi_b_ready(io_internal_vss_axi_full_0_b_ready),
		.m_axi_b_valid(io_internal_vss_axi_full_0_b_valid),
		.m_axi_b_bits_id(io_internal_vss_axi_full_0_b_bits_id),
		.m_axi_b_bits_resp(io_internal_vss_axi_full_0_b_bits_resp)
	);
	AxiWriteBuffer_2 module_0(
		.clock(clock),
		.reset(reset),
		.s_axi_ar_ready(_module_s_axi_ar_ready),
		.s_axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.s_axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.s_axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.s_axi_r_ready(_vssRvm_0_axi_r_ready),
		.s_axi_r_valid(_module_s_axi_r_valid),
		.s_axi_r_bits_data(_module_s_axi_r_bits_data),
		.s_axi_aw_ready(_module_s_axi_aw_ready),
		.s_axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.s_axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.s_axi_aw_bits_len(_vssRvm_0_axi_aw_bits_len),
		.s_axi_w_ready(_module_s_axi_w_ready),
		.s_axi_w_valid(_vssRvm_0_axi_w_valid),
		.s_axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.s_axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.s_axi_b_valid(_module_s_axi_b_valid),
		.m_axi_ar_ready(_mux_s_axi_0_ar_ready),
		.m_axi_ar_valid(_module_m_axi_ar_valid),
		.m_axi_ar_bits_addr(_module_m_axi_ar_bits_addr),
		.m_axi_ar_bits_len(_module_m_axi_ar_bits_len),
		.m_axi_ar_bits_size(_module_m_axi_ar_bits_size),
		.m_axi_ar_bits_burst(_module_m_axi_ar_bits_burst),
		.m_axi_ar_bits_lock(_module_m_axi_ar_bits_lock),
		.m_axi_ar_bits_cache(_module_m_axi_ar_bits_cache),
		.m_axi_ar_bits_prot(_module_m_axi_ar_bits_prot),
		.m_axi_ar_bits_qos(_module_m_axi_ar_bits_qos),
		.m_axi_ar_bits_region(_module_m_axi_ar_bits_region),
		.m_axi_r_ready(_module_m_axi_r_ready),
		.m_axi_r_valid(_mux_s_axi_0_r_valid),
		.m_axi_r_bits_data(_mux_s_axi_0_r_bits_data),
		.m_axi_aw_ready(_mux_s_axi_0_aw_ready),
		.m_axi_aw_valid(_module_m_axi_aw_valid),
		.m_axi_aw_bits_addr(_module_m_axi_aw_bits_addr),
		.m_axi_aw_bits_len(_module_m_axi_aw_bits_len),
		.m_axi_aw_bits_size(_module_m_axi_aw_bits_size),
		.m_axi_aw_bits_burst(_module_m_axi_aw_bits_burst),
		.m_axi_aw_bits_lock(_module_m_axi_aw_bits_lock),
		.m_axi_aw_bits_cache(_module_m_axi_aw_bits_cache),
		.m_axi_aw_bits_prot(_module_m_axi_aw_bits_prot),
		.m_axi_aw_bits_qos(_module_m_axi_aw_bits_qos),
		.m_axi_aw_bits_region(_module_m_axi_aw_bits_region),
		.m_axi_w_ready(_mux_s_axi_0_w_ready),
		.m_axi_w_valid(_module_m_axi_w_valid),
		.m_axi_w_bits_data(_module_m_axi_w_bits_data),
		.m_axi_w_bits_last(_module_m_axi_w_bits_last),
		.m_axi_b_valid(_mux_s_axi_0_b_valid)
	);
	AxiWriteBuffer_2 module_1(
		.clock(clock),
		.reset(reset),
		.s_axi_ar_ready(_module_1_s_axi_ar_ready),
		.s_axi_ar_valid(_vssRvm_1_axi_ar_valid),
		.s_axi_ar_bits_addr(_vssRvm_1_axi_ar_bits_addr),
		.s_axi_ar_bits_len(_vssRvm_1_axi_ar_bits_len),
		.s_axi_r_ready(_vssRvm_1_axi_r_ready),
		.s_axi_r_valid(_module_1_s_axi_r_valid),
		.s_axi_r_bits_data(_module_1_s_axi_r_bits_data),
		.s_axi_aw_ready(_module_1_s_axi_aw_ready),
		.s_axi_aw_valid(_vssRvm_1_axi_aw_valid),
		.s_axi_aw_bits_addr(_vssRvm_1_axi_aw_bits_addr),
		.s_axi_aw_bits_len(_vssRvm_1_axi_aw_bits_len),
		.s_axi_w_ready(_module_1_s_axi_w_ready),
		.s_axi_w_valid(_vssRvm_1_axi_w_valid),
		.s_axi_w_bits_data(_vssRvm_1_axi_w_bits_data),
		.s_axi_w_bits_last(_vssRvm_1_axi_w_bits_last),
		.s_axi_b_valid(_module_1_s_axi_b_valid),
		.m_axi_ar_ready(_mux_s_axi_1_ar_ready),
		.m_axi_ar_valid(_module_1_m_axi_ar_valid),
		.m_axi_ar_bits_addr(_module_1_m_axi_ar_bits_addr),
		.m_axi_ar_bits_len(_module_1_m_axi_ar_bits_len),
		.m_axi_ar_bits_size(_module_1_m_axi_ar_bits_size),
		.m_axi_ar_bits_burst(_module_1_m_axi_ar_bits_burst),
		.m_axi_ar_bits_lock(_module_1_m_axi_ar_bits_lock),
		.m_axi_ar_bits_cache(_module_1_m_axi_ar_bits_cache),
		.m_axi_ar_bits_prot(_module_1_m_axi_ar_bits_prot),
		.m_axi_ar_bits_qos(_module_1_m_axi_ar_bits_qos),
		.m_axi_ar_bits_region(_module_1_m_axi_ar_bits_region),
		.m_axi_r_ready(_module_1_m_axi_r_ready),
		.m_axi_r_valid(_mux_s_axi_1_r_valid),
		.m_axi_r_bits_data(_mux_s_axi_1_r_bits_data),
		.m_axi_aw_ready(_mux_s_axi_1_aw_ready),
		.m_axi_aw_valid(_module_1_m_axi_aw_valid),
		.m_axi_aw_bits_addr(_module_1_m_axi_aw_bits_addr),
		.m_axi_aw_bits_len(_module_1_m_axi_aw_bits_len),
		.m_axi_aw_bits_size(_module_1_m_axi_aw_bits_size),
		.m_axi_aw_bits_burst(_module_1_m_axi_aw_bits_burst),
		.m_axi_aw_bits_lock(_module_1_m_axi_aw_bits_lock),
		.m_axi_aw_bits_cache(_module_1_m_axi_aw_bits_cache),
		.m_axi_aw_bits_prot(_module_1_m_axi_aw_bits_prot),
		.m_axi_aw_bits_qos(_module_1_m_axi_aw_bits_qos),
		.m_axi_aw_bits_region(_module_1_m_axi_aw_bits_region),
		.m_axi_w_ready(_mux_s_axi_1_w_ready),
		.m_axi_w_valid(_module_1_m_axi_w_valid),
		.m_axi_w_bits_data(_module_1_m_axi_w_bits_data),
		.m_axi_w_bits_last(_module_1_m_axi_w_bits_last),
		.m_axi_b_valid(_mux_s_axi_1_b_valid)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_0(
		.io_dataIn_TREADY(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_0_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_0_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_0_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_0_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_1(
		.io_dataIn_TREADY(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_1_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_1_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_1_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_1_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_2(
		.io_dataIn_TREADY(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_2_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_2_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_2_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_2_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_3(
		.io_dataIn_TREADY(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_3_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_3_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_3_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_3_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_4(
		.io_dataIn_TREADY(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_4_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_4_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_4_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_4_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_5(
		.io_dataIn_TREADY(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_5_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_5_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_5_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_5_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_6(
		.io_dataIn_TREADY(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_6_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_6_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_6_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_6_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_7(
		.io_dataIn_TREADY(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_7_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_7_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_7_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_7_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_8(
		.io_dataIn_TREADY(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_8_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_8_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_8_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_8_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_9(
		.io_dataIn_TREADY(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_9_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_9_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_9_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_9_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_10(
		.io_dataIn_TREADY(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_10_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_10_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_10_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_10_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_11(
		.io_dataIn_TREADY(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_11_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_11_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_11_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_11_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_12(
		.io_dataIn_TREADY(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_12_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_12_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_12_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_12_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_13(
		.io_dataIn_TREADY(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_13_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_13_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_13_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_13_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_14(
		.io_dataIn_TREADY(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_14_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_14_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_14_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_14_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_15(
		.io_dataIn_TREADY(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_15_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_15_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_15_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_15_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_16(
		.io_dataIn_TREADY(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_16_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_16_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_16_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_16_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_16_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_17(
		.io_dataIn_TREADY(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_17_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_17_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_17_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_17_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_17_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_18(
		.io_dataIn_TREADY(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_18_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_18_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_18_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_18_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_18_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_19(
		.io_dataIn_TREADY(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_19_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_19_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_19_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_19_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_19_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_20(
		.io_dataIn_TREADY(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_20_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_20_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_20_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_20_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_20_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_21(
		.io_dataIn_TREADY(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_21_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_21_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_21_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_21_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_21_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_22(
		.io_dataIn_TREADY(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_22_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_22_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_22_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_22_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_22_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_23(
		.io_dataIn_TREADY(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_23_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_23_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_23_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_23_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_23_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_24(
		.io_dataIn_TREADY(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_24_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_24_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_24_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_24_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_24_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_25(
		.io_dataIn_TREADY(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_25_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_25_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_25_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_25_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_25_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_26(
		.io_dataIn_TREADY(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_26_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_26_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_26_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_26_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_26_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_27(
		.io_dataIn_TREADY(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_27_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_27_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_27_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_27_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_27_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_28(
		.io_dataIn_TREADY(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_28_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_28_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_28_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_28_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_28_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_29(
		.io_dataIn_TREADY(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_29_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_29_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_29_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_29_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_29_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_30(
		.io_dataIn_TREADY(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_30_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_30_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_30_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_30_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_30_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_31(
		.io_dataIn_TREADY(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_31_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_31_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_31_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_31_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_31_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_32(
		.io_dataIn_TREADY(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_32_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_32_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_32_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_32_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_32_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_33(
		.io_dataIn_TREADY(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_33_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_33_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_33_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_33_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_33_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_34(
		.io_dataIn_TREADY(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_34_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_34_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_34_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_34_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_34_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_35(
		.io_dataIn_TREADY(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_35_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_35_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_35_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_35_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_35_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_36(
		.io_dataIn_TREADY(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_36_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_36_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_36_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_36_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_36_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_37(
		.io_dataIn_TREADY(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_37_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_37_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_37_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_37_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_37_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_38(
		.io_dataIn_TREADY(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_38_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_38_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_38_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_38_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_38_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_39(
		.io_dataIn_TREADY(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_39_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_39_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_39_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_39_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_39_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_40(
		.io_dataIn_TREADY(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_40_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_40_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_40_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_40_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_40_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_41(
		.io_dataIn_TREADY(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_41_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_41_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_41_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_41_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_41_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_42(
		.io_dataIn_TREADY(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_42_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_42_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_42_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_42_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_42_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_43(
		.io_dataIn_TREADY(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_43_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_43_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_43_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_43_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_43_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_44(
		.io_dataIn_TREADY(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_44_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_44_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_44_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_44_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_44_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_45(
		.io_dataIn_TREADY(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_45_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_45_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_45_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_45_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_45_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_46(
		.io_dataIn_TREADY(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_46_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_46_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_46_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_46_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_46_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_47(
		.io_dataIn_TREADY(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_47_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_47_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_47_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_47_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_47_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_48(
		.io_dataIn_TREADY(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_48_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_48_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_48_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_48_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_48_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_49(
		.io_dataIn_TREADY(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_49_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_49_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_49_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_49_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_49_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_50(
		.io_dataIn_TREADY(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_50_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_50_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_50_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_50_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_50_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_51(
		.io_dataIn_TREADY(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_51_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_51_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_51_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_51_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_51_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_52(
		.io_dataIn_TREADY(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_52_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_52_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_52_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_52_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_52_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_53(
		.io_dataIn_TREADY(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_53_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_53_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_53_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_53_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_53_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_54(
		.io_dataIn_TREADY(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_54_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_54_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_54_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_54_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_54_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_55(
		.io_dataIn_TREADY(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_55_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_55_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_55_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_55_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_55_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_56(
		.io_dataIn_TREADY(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_56_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_56_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_56_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_56_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_56_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_57(
		.io_dataIn_TREADY(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_57_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_57_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_57_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_57_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_57_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_58(
		.io_dataIn_TREADY(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_58_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_58_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_58_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_58_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_58_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_59(
		.io_dataIn_TREADY(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_59_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_59_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_59_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_59_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_59_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_60(
		.io_dataIn_TREADY(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_60_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_60_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_60_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_60_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_60_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_61(
		.io_dataIn_TREADY(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_61_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_61_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_61_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_61_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_61_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_62(
		.io_dataIn_TREADY(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_62_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_62_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_62_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_62_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_62_TDATA)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_63(
		.io_dataIn_TREADY(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_63_pop_valid),
		.io_dataIn_TDATA(_stealNW_TQ_io_connPE_63_pop_bits),
		.io_dataOut_TREADY(io_export_taskOut_63_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_63_TVALID),
		.io_dataOut_TDATA(io_export_taskOut_63_TDATA)
	);
endmodule
module AllocatorServerNetworkUnit (
	clock,
	reset,
	io_addressIn0_ready,
	io_addressIn0_valid,
	io_addressIn0_bits,
	io_addressIn1_ready,
	io_addressIn1_valid,
	io_addressIn1_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn0_ready;
	input io_addressIn0_valid;
	input [63:0] io_addressIn0_bits;
	output wire io_addressIn1_ready;
	input io_addressIn1_valid;
	input [63:0] io_addressIn1_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	reg priorityReg;
	wire io_addressIn0_ready_0 = stateReg == 2'h0;
	wire _GEN = stateReg == 2'h1;
	wire _GEN_0 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
			priorityReg <= 1'h1;
		end
		else if (io_addressIn0_ready_0) begin
			if (io_addressIn0_valid) begin
				stateReg <= 2'h2;
				addressReg <= io_addressIn0_bits;
				priorityReg <= ~priorityReg;
			end
			else begin
				if (io_addressIn1_valid)
					stateReg <= 2'h1;
				priorityReg <= io_addressIn1_valid ^ priorityReg;
			end
		end
		else begin
			if (_GEN) begin
				if (io_addressIn1_valid) begin
					stateReg <= 2'h2;
					priorityReg <= ~priorityReg;
				end
				else begin
					if (io_addressIn0_valid)
						stateReg <= 2'h0;
					priorityReg <= io_addressIn0_valid ^ priorityReg;
				end
			end
			else if (_GEN_0 & io_addressOut_ready)
				stateReg <= {1'h0, ~priorityReg};
			if (_GEN & io_addressIn1_valid)
				addressReg <= io_addressIn1_bits;
		end
	assign io_addressIn0_ready = io_addressIn0_ready_0;
	assign io_addressIn1_ready = ~io_addressIn0_ready_0 & _GEN;
	assign io_addressOut_valid = ~(io_addressIn0_ready_0 | _GEN) & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module AllocatorNetworkUnit (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits,
	io_casAddressOut_ready,
	io_casAddressOut_valid,
	io_casAddressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	input io_casAddressOut_ready;
	output wire io_casAddressOut_valid;
	output wire [63:0] io_casAddressOut_bits;
	reg stateReg;
	reg [63:0] addressReg;
	reg priorityReg;
	wire _GEN = io_addressOut_ready & io_casAddressOut_ready;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 1'h0;
			addressReg <= 64'h0000000000000000;
			priorityReg <= 1'h1;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_0;
			_GEN_0 = io_addressOut_ready | io_casAddressOut_ready;
			if (stateReg)
				stateReg <= stateReg & ~_GEN_0;
			else
				stateReg <= io_addressIn_valid | stateReg;
			if (~stateReg & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
			priorityReg <= (stateReg & _GEN_0) ^ priorityReg;
		end
	assign io_addressIn_ready = ~stateReg;
	assign io_addressOut_valid = stateReg & (_GEN ? ~priorityReg & io_addressOut_ready : ~io_casAddressOut_ready & io_addressOut_ready);
	assign io_addressOut_bits = addressReg;
	assign io_casAddressOut_valid = (stateReg & (~_GEN | priorityReg)) & io_casAddressOut_ready;
	assign io_casAddressOut_bits = addressReg;
endmodule
module AllocatorClient (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg stateReg;
	reg [63:0] addressReg;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 1'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (stateReg)
				stateReg <= stateReg & ~io_addressOut_ready;
			else
				stateReg <= io_addressIn_valid | stateReg;
			if (~stateReg & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = ~stateReg;
	assign io_addressOut_valid = stateReg;
	assign io_addressOut_bits = addressReg;
endmodule
module ram_16x64 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [3:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [63:0] R0_data;
	input [3:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [63:0] W0_data;
	reg [63:0] Memory [0:15];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue16_UInt_4 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits;
	reg [3:0] enq_ptr_value;
	reg [3:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 4'h0;
			deq_ptr_value <= 4'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 4'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 4'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_16x64 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module AllocatorBuffer (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	Queue16_UInt_4 q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_addressIn_ready),
		.io_enq_valid(io_addressIn_valid),
		.io_enq_bits(io_addressIn_bits),
		.io_deq_ready(io_addressOut_ready),
		.io_deq_valid(io_addressOut_valid),
		.io_deq_bits(io_addressOut_bits)
	);
endmodule
module AllocatorNetwork (
	clock,
	reset,
	io_connVCAS_0_ready,
	io_connVCAS_0_valid,
	io_connVCAS_0_bits,
	io_connVCAS_1_ready,
	io_connVCAS_1_valid,
	io_connVCAS_1_bits,
	io_connVCAS_2_ready,
	io_connVCAS_2_valid,
	io_connVCAS_2_bits,
	io_connVCAS_3_ready,
	io_connVCAS_3_valid,
	io_connVCAS_3_bits,
	io_connPE_0_ready,
	io_connPE_0_valid,
	io_connPE_0_bits,
	io_connPE_1_ready,
	io_connPE_1_valid,
	io_connPE_1_bits,
	io_connPE_2_ready,
	io_connPE_2_valid,
	io_connPE_2_bits,
	io_connPE_3_ready,
	io_connPE_3_valid,
	io_connPE_3_bits,
	io_connPE_4_ready,
	io_connPE_4_valid,
	io_connPE_4_bits,
	io_connPE_5_ready,
	io_connPE_5_valid,
	io_connPE_5_bits,
	io_connPE_6_ready,
	io_connPE_6_valid,
	io_connPE_6_bits,
	io_connPE_7_ready,
	io_connPE_7_valid,
	io_connPE_7_bits,
	io_connPE_8_ready,
	io_connPE_8_valid,
	io_connPE_8_bits,
	io_connPE_9_ready,
	io_connPE_9_valid,
	io_connPE_9_bits,
	io_connPE_10_ready,
	io_connPE_10_valid,
	io_connPE_10_bits,
	io_connPE_11_ready,
	io_connPE_11_valid,
	io_connPE_11_bits,
	io_connPE_12_ready,
	io_connPE_12_valid,
	io_connPE_12_bits,
	io_connPE_13_ready,
	io_connPE_13_valid,
	io_connPE_13_bits,
	io_connPE_14_ready,
	io_connPE_14_valid,
	io_connPE_14_bits,
	io_connPE_15_ready,
	io_connPE_15_valid,
	io_connPE_15_bits,
	io_connPE_16_ready,
	io_connPE_16_valid,
	io_connPE_16_bits,
	io_connPE_17_ready,
	io_connPE_17_valid,
	io_connPE_17_bits,
	io_connPE_18_ready,
	io_connPE_18_valid,
	io_connPE_18_bits,
	io_connPE_19_ready,
	io_connPE_19_valid,
	io_connPE_19_bits,
	io_connPE_20_ready,
	io_connPE_20_valid,
	io_connPE_20_bits,
	io_connPE_21_ready,
	io_connPE_21_valid,
	io_connPE_21_bits,
	io_connPE_22_ready,
	io_connPE_22_valid,
	io_connPE_22_bits,
	io_connPE_23_ready,
	io_connPE_23_valid,
	io_connPE_23_bits,
	io_connPE_24_ready,
	io_connPE_24_valid,
	io_connPE_24_bits,
	io_connPE_25_ready,
	io_connPE_25_valid,
	io_connPE_25_bits,
	io_connPE_26_ready,
	io_connPE_26_valid,
	io_connPE_26_bits,
	io_connPE_27_ready,
	io_connPE_27_valid,
	io_connPE_27_bits,
	io_connPE_28_ready,
	io_connPE_28_valid,
	io_connPE_28_bits,
	io_connPE_29_ready,
	io_connPE_29_valid,
	io_connPE_29_bits,
	io_connPE_30_ready,
	io_connPE_30_valid,
	io_connPE_30_bits,
	io_connPE_31_ready,
	io_connPE_31_valid,
	io_connPE_31_bits,
	io_connPE_32_ready,
	io_connPE_32_valid,
	io_connPE_32_bits,
	io_connPE_33_ready,
	io_connPE_33_valid,
	io_connPE_33_bits,
	io_connPE_34_ready,
	io_connPE_34_valid,
	io_connPE_34_bits,
	io_connPE_35_ready,
	io_connPE_35_valid,
	io_connPE_35_bits,
	io_connPE_36_ready,
	io_connPE_36_valid,
	io_connPE_36_bits,
	io_connPE_37_ready,
	io_connPE_37_valid,
	io_connPE_37_bits,
	io_connPE_38_ready,
	io_connPE_38_valid,
	io_connPE_38_bits,
	io_connPE_39_ready,
	io_connPE_39_valid,
	io_connPE_39_bits,
	io_connPE_40_ready,
	io_connPE_40_valid,
	io_connPE_40_bits,
	io_connPE_41_ready,
	io_connPE_41_valid,
	io_connPE_41_bits,
	io_connPE_42_ready,
	io_connPE_42_valid,
	io_connPE_42_bits,
	io_connPE_43_ready,
	io_connPE_43_valid,
	io_connPE_43_bits,
	io_connPE_44_ready,
	io_connPE_44_valid,
	io_connPE_44_bits,
	io_connPE_45_ready,
	io_connPE_45_valid,
	io_connPE_45_bits,
	io_connPE_46_ready,
	io_connPE_46_valid,
	io_connPE_46_bits,
	io_connPE_47_ready,
	io_connPE_47_valid,
	io_connPE_47_bits,
	io_connPE_48_ready,
	io_connPE_48_valid,
	io_connPE_48_bits,
	io_connPE_49_ready,
	io_connPE_49_valid,
	io_connPE_49_bits,
	io_connPE_50_ready,
	io_connPE_50_valid,
	io_connPE_50_bits,
	io_connPE_51_ready,
	io_connPE_51_valid,
	io_connPE_51_bits,
	io_connPE_52_ready,
	io_connPE_52_valid,
	io_connPE_52_bits,
	io_connPE_53_ready,
	io_connPE_53_valid,
	io_connPE_53_bits,
	io_connPE_54_ready,
	io_connPE_54_valid,
	io_connPE_54_bits,
	io_connPE_55_ready,
	io_connPE_55_valid,
	io_connPE_55_bits,
	io_connPE_56_ready,
	io_connPE_56_valid,
	io_connPE_56_bits,
	io_connPE_57_ready,
	io_connPE_57_valid,
	io_connPE_57_bits,
	io_connPE_58_ready,
	io_connPE_58_valid,
	io_connPE_58_bits,
	io_connPE_59_ready,
	io_connPE_59_valid,
	io_connPE_59_bits,
	io_connPE_60_ready,
	io_connPE_60_valid,
	io_connPE_60_bits,
	io_connPE_61_ready,
	io_connPE_61_valid,
	io_connPE_61_bits,
	io_connPE_62_ready,
	io_connPE_62_valid,
	io_connPE_62_bits,
	io_connPE_63_ready,
	io_connPE_63_valid,
	io_connPE_63_bits
);
	input clock;
	input reset;
	output wire io_connVCAS_0_ready;
	input io_connVCAS_0_valid;
	input [63:0] io_connVCAS_0_bits;
	output wire io_connVCAS_1_ready;
	input io_connVCAS_1_valid;
	input [63:0] io_connVCAS_1_bits;
	output wire io_connVCAS_2_ready;
	input io_connVCAS_2_valid;
	input [63:0] io_connVCAS_2_bits;
	output wire io_connVCAS_3_ready;
	input io_connVCAS_3_valid;
	input [63:0] io_connVCAS_3_bits;
	input io_connPE_0_ready;
	output wire io_connPE_0_valid;
	output wire [63:0] io_connPE_0_bits;
	input io_connPE_1_ready;
	output wire io_connPE_1_valid;
	output wire [63:0] io_connPE_1_bits;
	input io_connPE_2_ready;
	output wire io_connPE_2_valid;
	output wire [63:0] io_connPE_2_bits;
	input io_connPE_3_ready;
	output wire io_connPE_3_valid;
	output wire [63:0] io_connPE_3_bits;
	input io_connPE_4_ready;
	output wire io_connPE_4_valid;
	output wire [63:0] io_connPE_4_bits;
	input io_connPE_5_ready;
	output wire io_connPE_5_valid;
	output wire [63:0] io_connPE_5_bits;
	input io_connPE_6_ready;
	output wire io_connPE_6_valid;
	output wire [63:0] io_connPE_6_bits;
	input io_connPE_7_ready;
	output wire io_connPE_7_valid;
	output wire [63:0] io_connPE_7_bits;
	input io_connPE_8_ready;
	output wire io_connPE_8_valid;
	output wire [63:0] io_connPE_8_bits;
	input io_connPE_9_ready;
	output wire io_connPE_9_valid;
	output wire [63:0] io_connPE_9_bits;
	input io_connPE_10_ready;
	output wire io_connPE_10_valid;
	output wire [63:0] io_connPE_10_bits;
	input io_connPE_11_ready;
	output wire io_connPE_11_valid;
	output wire [63:0] io_connPE_11_bits;
	input io_connPE_12_ready;
	output wire io_connPE_12_valid;
	output wire [63:0] io_connPE_12_bits;
	input io_connPE_13_ready;
	output wire io_connPE_13_valid;
	output wire [63:0] io_connPE_13_bits;
	input io_connPE_14_ready;
	output wire io_connPE_14_valid;
	output wire [63:0] io_connPE_14_bits;
	input io_connPE_15_ready;
	output wire io_connPE_15_valid;
	output wire [63:0] io_connPE_15_bits;
	input io_connPE_16_ready;
	output wire io_connPE_16_valid;
	output wire [63:0] io_connPE_16_bits;
	input io_connPE_17_ready;
	output wire io_connPE_17_valid;
	output wire [63:0] io_connPE_17_bits;
	input io_connPE_18_ready;
	output wire io_connPE_18_valid;
	output wire [63:0] io_connPE_18_bits;
	input io_connPE_19_ready;
	output wire io_connPE_19_valid;
	output wire [63:0] io_connPE_19_bits;
	input io_connPE_20_ready;
	output wire io_connPE_20_valid;
	output wire [63:0] io_connPE_20_bits;
	input io_connPE_21_ready;
	output wire io_connPE_21_valid;
	output wire [63:0] io_connPE_21_bits;
	input io_connPE_22_ready;
	output wire io_connPE_22_valid;
	output wire [63:0] io_connPE_22_bits;
	input io_connPE_23_ready;
	output wire io_connPE_23_valid;
	output wire [63:0] io_connPE_23_bits;
	input io_connPE_24_ready;
	output wire io_connPE_24_valid;
	output wire [63:0] io_connPE_24_bits;
	input io_connPE_25_ready;
	output wire io_connPE_25_valid;
	output wire [63:0] io_connPE_25_bits;
	input io_connPE_26_ready;
	output wire io_connPE_26_valid;
	output wire [63:0] io_connPE_26_bits;
	input io_connPE_27_ready;
	output wire io_connPE_27_valid;
	output wire [63:0] io_connPE_27_bits;
	input io_connPE_28_ready;
	output wire io_connPE_28_valid;
	output wire [63:0] io_connPE_28_bits;
	input io_connPE_29_ready;
	output wire io_connPE_29_valid;
	output wire [63:0] io_connPE_29_bits;
	input io_connPE_30_ready;
	output wire io_connPE_30_valid;
	output wire [63:0] io_connPE_30_bits;
	input io_connPE_31_ready;
	output wire io_connPE_31_valid;
	output wire [63:0] io_connPE_31_bits;
	input io_connPE_32_ready;
	output wire io_connPE_32_valid;
	output wire [63:0] io_connPE_32_bits;
	input io_connPE_33_ready;
	output wire io_connPE_33_valid;
	output wire [63:0] io_connPE_33_bits;
	input io_connPE_34_ready;
	output wire io_connPE_34_valid;
	output wire [63:0] io_connPE_34_bits;
	input io_connPE_35_ready;
	output wire io_connPE_35_valid;
	output wire [63:0] io_connPE_35_bits;
	input io_connPE_36_ready;
	output wire io_connPE_36_valid;
	output wire [63:0] io_connPE_36_bits;
	input io_connPE_37_ready;
	output wire io_connPE_37_valid;
	output wire [63:0] io_connPE_37_bits;
	input io_connPE_38_ready;
	output wire io_connPE_38_valid;
	output wire [63:0] io_connPE_38_bits;
	input io_connPE_39_ready;
	output wire io_connPE_39_valid;
	output wire [63:0] io_connPE_39_bits;
	input io_connPE_40_ready;
	output wire io_connPE_40_valid;
	output wire [63:0] io_connPE_40_bits;
	input io_connPE_41_ready;
	output wire io_connPE_41_valid;
	output wire [63:0] io_connPE_41_bits;
	input io_connPE_42_ready;
	output wire io_connPE_42_valid;
	output wire [63:0] io_connPE_42_bits;
	input io_connPE_43_ready;
	output wire io_connPE_43_valid;
	output wire [63:0] io_connPE_43_bits;
	input io_connPE_44_ready;
	output wire io_connPE_44_valid;
	output wire [63:0] io_connPE_44_bits;
	input io_connPE_45_ready;
	output wire io_connPE_45_valid;
	output wire [63:0] io_connPE_45_bits;
	input io_connPE_46_ready;
	output wire io_connPE_46_valid;
	output wire [63:0] io_connPE_46_bits;
	input io_connPE_47_ready;
	output wire io_connPE_47_valid;
	output wire [63:0] io_connPE_47_bits;
	input io_connPE_48_ready;
	output wire io_connPE_48_valid;
	output wire [63:0] io_connPE_48_bits;
	input io_connPE_49_ready;
	output wire io_connPE_49_valid;
	output wire [63:0] io_connPE_49_bits;
	input io_connPE_50_ready;
	output wire io_connPE_50_valid;
	output wire [63:0] io_connPE_50_bits;
	input io_connPE_51_ready;
	output wire io_connPE_51_valid;
	output wire [63:0] io_connPE_51_bits;
	input io_connPE_52_ready;
	output wire io_connPE_52_valid;
	output wire [63:0] io_connPE_52_bits;
	input io_connPE_53_ready;
	output wire io_connPE_53_valid;
	output wire [63:0] io_connPE_53_bits;
	input io_connPE_54_ready;
	output wire io_connPE_54_valid;
	output wire [63:0] io_connPE_54_bits;
	input io_connPE_55_ready;
	output wire io_connPE_55_valid;
	output wire [63:0] io_connPE_55_bits;
	input io_connPE_56_ready;
	output wire io_connPE_56_valid;
	output wire [63:0] io_connPE_56_bits;
	input io_connPE_57_ready;
	output wire io_connPE_57_valid;
	output wire [63:0] io_connPE_57_bits;
	input io_connPE_58_ready;
	output wire io_connPE_58_valid;
	output wire [63:0] io_connPE_58_bits;
	input io_connPE_59_ready;
	output wire io_connPE_59_valid;
	output wire [63:0] io_connPE_59_bits;
	input io_connPE_60_ready;
	output wire io_connPE_60_valid;
	output wire [63:0] io_connPE_60_bits;
	input io_connPE_61_ready;
	output wire io_connPE_61_valid;
	output wire [63:0] io_connPE_61_bits;
	input io_connPE_62_ready;
	output wire io_connPE_62_valid;
	output wire [63:0] io_connPE_62_bits;
	input io_connPE_63_ready;
	output wire io_connPE_63_valid;
	output wire [63:0] io_connPE_63_bits;
	wire _queues_63_io_addressIn_ready;
	wire _queues_62_io_addressIn_ready;
	wire _queues_61_io_addressIn_ready;
	wire _queues_60_io_addressIn_ready;
	wire _queues_59_io_addressIn_ready;
	wire _queues_58_io_addressIn_ready;
	wire _queues_57_io_addressIn_ready;
	wire _queues_56_io_addressIn_ready;
	wire _queues_55_io_addressIn_ready;
	wire _queues_54_io_addressIn_ready;
	wire _queues_53_io_addressIn_ready;
	wire _queues_52_io_addressIn_ready;
	wire _queues_51_io_addressIn_ready;
	wire _queues_50_io_addressIn_ready;
	wire _queues_49_io_addressIn_ready;
	wire _queues_48_io_addressIn_ready;
	wire _queues_47_io_addressIn_ready;
	wire _queues_46_io_addressIn_ready;
	wire _queues_45_io_addressIn_ready;
	wire _queues_44_io_addressIn_ready;
	wire _queues_43_io_addressIn_ready;
	wire _queues_42_io_addressIn_ready;
	wire _queues_41_io_addressIn_ready;
	wire _queues_40_io_addressIn_ready;
	wire _queues_39_io_addressIn_ready;
	wire _queues_38_io_addressIn_ready;
	wire _queues_37_io_addressIn_ready;
	wire _queues_36_io_addressIn_ready;
	wire _queues_35_io_addressIn_ready;
	wire _queues_34_io_addressIn_ready;
	wire _queues_33_io_addressIn_ready;
	wire _queues_32_io_addressIn_ready;
	wire _queues_31_io_addressIn_ready;
	wire _queues_30_io_addressIn_ready;
	wire _queues_29_io_addressIn_ready;
	wire _queues_28_io_addressIn_ready;
	wire _queues_27_io_addressIn_ready;
	wire _queues_26_io_addressIn_ready;
	wire _queues_25_io_addressIn_ready;
	wire _queues_24_io_addressIn_ready;
	wire _queues_23_io_addressIn_ready;
	wire _queues_22_io_addressIn_ready;
	wire _queues_21_io_addressIn_ready;
	wire _queues_20_io_addressIn_ready;
	wire _queues_19_io_addressIn_ready;
	wire _queues_18_io_addressIn_ready;
	wire _queues_17_io_addressIn_ready;
	wire _queues_16_io_addressIn_ready;
	wire _queues_15_io_addressIn_ready;
	wire _queues_14_io_addressIn_ready;
	wire _queues_13_io_addressIn_ready;
	wire _queues_12_io_addressIn_ready;
	wire _queues_11_io_addressIn_ready;
	wire _queues_10_io_addressIn_ready;
	wire _queues_9_io_addressIn_ready;
	wire _queues_8_io_addressIn_ready;
	wire _queues_7_io_addressIn_ready;
	wire _queues_6_io_addressIn_ready;
	wire _queues_5_io_addressIn_ready;
	wire _queues_4_io_addressIn_ready;
	wire _queues_3_io_addressIn_ready;
	wire _queues_2_io_addressIn_ready;
	wire _queues_1_io_addressIn_ready;
	wire _queues_0_io_addressIn_ready;
	wire _casServers_63_io_addressIn_ready;
	wire _casServers_63_io_addressOut_valid;
	wire [63:0] _casServers_63_io_addressOut_bits;
	wire _casServers_62_io_addressIn_ready;
	wire _casServers_62_io_addressOut_valid;
	wire [63:0] _casServers_62_io_addressOut_bits;
	wire _casServers_61_io_addressIn_ready;
	wire _casServers_61_io_addressOut_valid;
	wire [63:0] _casServers_61_io_addressOut_bits;
	wire _casServers_60_io_addressIn_ready;
	wire _casServers_60_io_addressOut_valid;
	wire [63:0] _casServers_60_io_addressOut_bits;
	wire _casServers_59_io_addressIn_ready;
	wire _casServers_59_io_addressOut_valid;
	wire [63:0] _casServers_59_io_addressOut_bits;
	wire _casServers_58_io_addressIn_ready;
	wire _casServers_58_io_addressOut_valid;
	wire [63:0] _casServers_58_io_addressOut_bits;
	wire _casServers_57_io_addressIn_ready;
	wire _casServers_57_io_addressOut_valid;
	wire [63:0] _casServers_57_io_addressOut_bits;
	wire _casServers_56_io_addressIn_ready;
	wire _casServers_56_io_addressOut_valid;
	wire [63:0] _casServers_56_io_addressOut_bits;
	wire _casServers_55_io_addressIn_ready;
	wire _casServers_55_io_addressOut_valid;
	wire [63:0] _casServers_55_io_addressOut_bits;
	wire _casServers_54_io_addressIn_ready;
	wire _casServers_54_io_addressOut_valid;
	wire [63:0] _casServers_54_io_addressOut_bits;
	wire _casServers_53_io_addressIn_ready;
	wire _casServers_53_io_addressOut_valid;
	wire [63:0] _casServers_53_io_addressOut_bits;
	wire _casServers_52_io_addressIn_ready;
	wire _casServers_52_io_addressOut_valid;
	wire [63:0] _casServers_52_io_addressOut_bits;
	wire _casServers_51_io_addressIn_ready;
	wire _casServers_51_io_addressOut_valid;
	wire [63:0] _casServers_51_io_addressOut_bits;
	wire _casServers_50_io_addressIn_ready;
	wire _casServers_50_io_addressOut_valid;
	wire [63:0] _casServers_50_io_addressOut_bits;
	wire _casServers_49_io_addressIn_ready;
	wire _casServers_49_io_addressOut_valid;
	wire [63:0] _casServers_49_io_addressOut_bits;
	wire _casServers_48_io_addressIn_ready;
	wire _casServers_48_io_addressOut_valid;
	wire [63:0] _casServers_48_io_addressOut_bits;
	wire _casServers_47_io_addressIn_ready;
	wire _casServers_47_io_addressOut_valid;
	wire [63:0] _casServers_47_io_addressOut_bits;
	wire _casServers_46_io_addressIn_ready;
	wire _casServers_46_io_addressOut_valid;
	wire [63:0] _casServers_46_io_addressOut_bits;
	wire _casServers_45_io_addressIn_ready;
	wire _casServers_45_io_addressOut_valid;
	wire [63:0] _casServers_45_io_addressOut_bits;
	wire _casServers_44_io_addressIn_ready;
	wire _casServers_44_io_addressOut_valid;
	wire [63:0] _casServers_44_io_addressOut_bits;
	wire _casServers_43_io_addressIn_ready;
	wire _casServers_43_io_addressOut_valid;
	wire [63:0] _casServers_43_io_addressOut_bits;
	wire _casServers_42_io_addressIn_ready;
	wire _casServers_42_io_addressOut_valid;
	wire [63:0] _casServers_42_io_addressOut_bits;
	wire _casServers_41_io_addressIn_ready;
	wire _casServers_41_io_addressOut_valid;
	wire [63:0] _casServers_41_io_addressOut_bits;
	wire _casServers_40_io_addressIn_ready;
	wire _casServers_40_io_addressOut_valid;
	wire [63:0] _casServers_40_io_addressOut_bits;
	wire _casServers_39_io_addressIn_ready;
	wire _casServers_39_io_addressOut_valid;
	wire [63:0] _casServers_39_io_addressOut_bits;
	wire _casServers_38_io_addressIn_ready;
	wire _casServers_38_io_addressOut_valid;
	wire [63:0] _casServers_38_io_addressOut_bits;
	wire _casServers_37_io_addressIn_ready;
	wire _casServers_37_io_addressOut_valid;
	wire [63:0] _casServers_37_io_addressOut_bits;
	wire _casServers_36_io_addressIn_ready;
	wire _casServers_36_io_addressOut_valid;
	wire [63:0] _casServers_36_io_addressOut_bits;
	wire _casServers_35_io_addressIn_ready;
	wire _casServers_35_io_addressOut_valid;
	wire [63:0] _casServers_35_io_addressOut_bits;
	wire _casServers_34_io_addressIn_ready;
	wire _casServers_34_io_addressOut_valid;
	wire [63:0] _casServers_34_io_addressOut_bits;
	wire _casServers_33_io_addressIn_ready;
	wire _casServers_33_io_addressOut_valid;
	wire [63:0] _casServers_33_io_addressOut_bits;
	wire _casServers_32_io_addressIn_ready;
	wire _casServers_32_io_addressOut_valid;
	wire [63:0] _casServers_32_io_addressOut_bits;
	wire _casServers_31_io_addressIn_ready;
	wire _casServers_31_io_addressOut_valid;
	wire [63:0] _casServers_31_io_addressOut_bits;
	wire _casServers_30_io_addressIn_ready;
	wire _casServers_30_io_addressOut_valid;
	wire [63:0] _casServers_30_io_addressOut_bits;
	wire _casServers_29_io_addressIn_ready;
	wire _casServers_29_io_addressOut_valid;
	wire [63:0] _casServers_29_io_addressOut_bits;
	wire _casServers_28_io_addressIn_ready;
	wire _casServers_28_io_addressOut_valid;
	wire [63:0] _casServers_28_io_addressOut_bits;
	wire _casServers_27_io_addressIn_ready;
	wire _casServers_27_io_addressOut_valid;
	wire [63:0] _casServers_27_io_addressOut_bits;
	wire _casServers_26_io_addressIn_ready;
	wire _casServers_26_io_addressOut_valid;
	wire [63:0] _casServers_26_io_addressOut_bits;
	wire _casServers_25_io_addressIn_ready;
	wire _casServers_25_io_addressOut_valid;
	wire [63:0] _casServers_25_io_addressOut_bits;
	wire _casServers_24_io_addressIn_ready;
	wire _casServers_24_io_addressOut_valid;
	wire [63:0] _casServers_24_io_addressOut_bits;
	wire _casServers_23_io_addressIn_ready;
	wire _casServers_23_io_addressOut_valid;
	wire [63:0] _casServers_23_io_addressOut_bits;
	wire _casServers_22_io_addressIn_ready;
	wire _casServers_22_io_addressOut_valid;
	wire [63:0] _casServers_22_io_addressOut_bits;
	wire _casServers_21_io_addressIn_ready;
	wire _casServers_21_io_addressOut_valid;
	wire [63:0] _casServers_21_io_addressOut_bits;
	wire _casServers_20_io_addressIn_ready;
	wire _casServers_20_io_addressOut_valid;
	wire [63:0] _casServers_20_io_addressOut_bits;
	wire _casServers_19_io_addressIn_ready;
	wire _casServers_19_io_addressOut_valid;
	wire [63:0] _casServers_19_io_addressOut_bits;
	wire _casServers_18_io_addressIn_ready;
	wire _casServers_18_io_addressOut_valid;
	wire [63:0] _casServers_18_io_addressOut_bits;
	wire _casServers_17_io_addressIn_ready;
	wire _casServers_17_io_addressOut_valid;
	wire [63:0] _casServers_17_io_addressOut_bits;
	wire _casServers_16_io_addressIn_ready;
	wire _casServers_16_io_addressOut_valid;
	wire [63:0] _casServers_16_io_addressOut_bits;
	wire _casServers_15_io_addressIn_ready;
	wire _casServers_15_io_addressOut_valid;
	wire [63:0] _casServers_15_io_addressOut_bits;
	wire _casServers_14_io_addressIn_ready;
	wire _casServers_14_io_addressOut_valid;
	wire [63:0] _casServers_14_io_addressOut_bits;
	wire _casServers_13_io_addressIn_ready;
	wire _casServers_13_io_addressOut_valid;
	wire [63:0] _casServers_13_io_addressOut_bits;
	wire _casServers_12_io_addressIn_ready;
	wire _casServers_12_io_addressOut_valid;
	wire [63:0] _casServers_12_io_addressOut_bits;
	wire _casServers_11_io_addressIn_ready;
	wire _casServers_11_io_addressOut_valid;
	wire [63:0] _casServers_11_io_addressOut_bits;
	wire _casServers_10_io_addressIn_ready;
	wire _casServers_10_io_addressOut_valid;
	wire [63:0] _casServers_10_io_addressOut_bits;
	wire _casServers_9_io_addressIn_ready;
	wire _casServers_9_io_addressOut_valid;
	wire [63:0] _casServers_9_io_addressOut_bits;
	wire _casServers_8_io_addressIn_ready;
	wire _casServers_8_io_addressOut_valid;
	wire [63:0] _casServers_8_io_addressOut_bits;
	wire _casServers_7_io_addressIn_ready;
	wire _casServers_7_io_addressOut_valid;
	wire [63:0] _casServers_7_io_addressOut_bits;
	wire _casServers_6_io_addressIn_ready;
	wire _casServers_6_io_addressOut_valid;
	wire [63:0] _casServers_6_io_addressOut_bits;
	wire _casServers_5_io_addressIn_ready;
	wire _casServers_5_io_addressOut_valid;
	wire [63:0] _casServers_5_io_addressOut_bits;
	wire _casServers_4_io_addressIn_ready;
	wire _casServers_4_io_addressOut_valid;
	wire [63:0] _casServers_4_io_addressOut_bits;
	wire _casServers_3_io_addressIn_ready;
	wire _casServers_3_io_addressOut_valid;
	wire [63:0] _casServers_3_io_addressOut_bits;
	wire _casServers_2_io_addressIn_ready;
	wire _casServers_2_io_addressOut_valid;
	wire [63:0] _casServers_2_io_addressOut_bits;
	wire _casServers_1_io_addressIn_ready;
	wire _casServers_1_io_addressOut_valid;
	wire [63:0] _casServers_1_io_addressOut_bits;
	wire _casServers_0_io_addressIn_ready;
	wire _casServers_0_io_addressOut_valid;
	wire [63:0] _casServers_0_io_addressOut_bits;
	wire _networkUnits_63_io_addressIn_ready;
	wire _networkUnits_63_io_casAddressOut_valid;
	wire [63:0] _networkUnits_63_io_casAddressOut_bits;
	wire _networkUnits_62_io_addressIn_ready;
	wire _networkUnits_62_io_addressOut_valid;
	wire [63:0] _networkUnits_62_io_addressOut_bits;
	wire _networkUnits_62_io_casAddressOut_valid;
	wire [63:0] _networkUnits_62_io_casAddressOut_bits;
	wire _networkUnits_61_io_addressIn_ready;
	wire _networkUnits_61_io_addressOut_valid;
	wire [63:0] _networkUnits_61_io_addressOut_bits;
	wire _networkUnits_61_io_casAddressOut_valid;
	wire [63:0] _networkUnits_61_io_casAddressOut_bits;
	wire _networkUnits_60_io_addressIn_ready;
	wire _networkUnits_60_io_addressOut_valid;
	wire [63:0] _networkUnits_60_io_addressOut_bits;
	wire _networkUnits_60_io_casAddressOut_valid;
	wire [63:0] _networkUnits_60_io_casAddressOut_bits;
	wire _networkUnits_59_io_addressIn_ready;
	wire _networkUnits_59_io_addressOut_valid;
	wire [63:0] _networkUnits_59_io_addressOut_bits;
	wire _networkUnits_59_io_casAddressOut_valid;
	wire [63:0] _networkUnits_59_io_casAddressOut_bits;
	wire _networkUnits_58_io_addressIn_ready;
	wire _networkUnits_58_io_addressOut_valid;
	wire [63:0] _networkUnits_58_io_addressOut_bits;
	wire _networkUnits_58_io_casAddressOut_valid;
	wire [63:0] _networkUnits_58_io_casAddressOut_bits;
	wire _networkUnits_57_io_addressIn_ready;
	wire _networkUnits_57_io_addressOut_valid;
	wire [63:0] _networkUnits_57_io_addressOut_bits;
	wire _networkUnits_57_io_casAddressOut_valid;
	wire [63:0] _networkUnits_57_io_casAddressOut_bits;
	wire _networkUnits_56_io_addressIn_ready;
	wire _networkUnits_56_io_addressOut_valid;
	wire [63:0] _networkUnits_56_io_addressOut_bits;
	wire _networkUnits_56_io_casAddressOut_valid;
	wire [63:0] _networkUnits_56_io_casAddressOut_bits;
	wire _networkUnits_55_io_addressIn_ready;
	wire _networkUnits_55_io_addressOut_valid;
	wire [63:0] _networkUnits_55_io_addressOut_bits;
	wire _networkUnits_55_io_casAddressOut_valid;
	wire [63:0] _networkUnits_55_io_casAddressOut_bits;
	wire _networkUnits_54_io_addressIn_ready;
	wire _networkUnits_54_io_addressOut_valid;
	wire [63:0] _networkUnits_54_io_addressOut_bits;
	wire _networkUnits_54_io_casAddressOut_valid;
	wire [63:0] _networkUnits_54_io_casAddressOut_bits;
	wire _networkUnits_53_io_addressIn_ready;
	wire _networkUnits_53_io_addressOut_valid;
	wire [63:0] _networkUnits_53_io_addressOut_bits;
	wire _networkUnits_53_io_casAddressOut_valid;
	wire [63:0] _networkUnits_53_io_casAddressOut_bits;
	wire _networkUnits_52_io_addressIn_ready;
	wire _networkUnits_52_io_addressOut_valid;
	wire [63:0] _networkUnits_52_io_addressOut_bits;
	wire _networkUnits_52_io_casAddressOut_valid;
	wire [63:0] _networkUnits_52_io_casAddressOut_bits;
	wire _networkUnits_51_io_addressIn_ready;
	wire _networkUnits_51_io_addressOut_valid;
	wire [63:0] _networkUnits_51_io_addressOut_bits;
	wire _networkUnits_51_io_casAddressOut_valid;
	wire [63:0] _networkUnits_51_io_casAddressOut_bits;
	wire _networkUnits_50_io_addressIn_ready;
	wire _networkUnits_50_io_addressOut_valid;
	wire [63:0] _networkUnits_50_io_addressOut_bits;
	wire _networkUnits_50_io_casAddressOut_valid;
	wire [63:0] _networkUnits_50_io_casAddressOut_bits;
	wire _networkUnits_49_io_addressIn_ready;
	wire _networkUnits_49_io_addressOut_valid;
	wire [63:0] _networkUnits_49_io_addressOut_bits;
	wire _networkUnits_49_io_casAddressOut_valid;
	wire [63:0] _networkUnits_49_io_casAddressOut_bits;
	wire _networkUnits_48_io_addressIn_ready;
	wire _networkUnits_48_io_addressOut_valid;
	wire [63:0] _networkUnits_48_io_addressOut_bits;
	wire _networkUnits_48_io_casAddressOut_valid;
	wire [63:0] _networkUnits_48_io_casAddressOut_bits;
	wire _networkUnits_47_io_addressIn_ready;
	wire _networkUnits_47_io_addressOut_valid;
	wire [63:0] _networkUnits_47_io_addressOut_bits;
	wire _networkUnits_47_io_casAddressOut_valid;
	wire [63:0] _networkUnits_47_io_casAddressOut_bits;
	wire _networkUnits_46_io_addressIn_ready;
	wire _networkUnits_46_io_addressOut_valid;
	wire [63:0] _networkUnits_46_io_addressOut_bits;
	wire _networkUnits_46_io_casAddressOut_valid;
	wire [63:0] _networkUnits_46_io_casAddressOut_bits;
	wire _networkUnits_45_io_addressIn_ready;
	wire _networkUnits_45_io_addressOut_valid;
	wire [63:0] _networkUnits_45_io_addressOut_bits;
	wire _networkUnits_45_io_casAddressOut_valid;
	wire [63:0] _networkUnits_45_io_casAddressOut_bits;
	wire _networkUnits_44_io_addressIn_ready;
	wire _networkUnits_44_io_addressOut_valid;
	wire [63:0] _networkUnits_44_io_addressOut_bits;
	wire _networkUnits_44_io_casAddressOut_valid;
	wire [63:0] _networkUnits_44_io_casAddressOut_bits;
	wire _networkUnits_43_io_addressIn_ready;
	wire _networkUnits_43_io_addressOut_valid;
	wire [63:0] _networkUnits_43_io_addressOut_bits;
	wire _networkUnits_43_io_casAddressOut_valid;
	wire [63:0] _networkUnits_43_io_casAddressOut_bits;
	wire _networkUnits_42_io_addressIn_ready;
	wire _networkUnits_42_io_addressOut_valid;
	wire [63:0] _networkUnits_42_io_addressOut_bits;
	wire _networkUnits_42_io_casAddressOut_valid;
	wire [63:0] _networkUnits_42_io_casAddressOut_bits;
	wire _networkUnits_41_io_addressIn_ready;
	wire _networkUnits_41_io_addressOut_valid;
	wire [63:0] _networkUnits_41_io_addressOut_bits;
	wire _networkUnits_41_io_casAddressOut_valid;
	wire [63:0] _networkUnits_41_io_casAddressOut_bits;
	wire _networkUnits_40_io_addressIn_ready;
	wire _networkUnits_40_io_addressOut_valid;
	wire [63:0] _networkUnits_40_io_addressOut_bits;
	wire _networkUnits_40_io_casAddressOut_valid;
	wire [63:0] _networkUnits_40_io_casAddressOut_bits;
	wire _networkUnits_39_io_addressIn_ready;
	wire _networkUnits_39_io_addressOut_valid;
	wire [63:0] _networkUnits_39_io_addressOut_bits;
	wire _networkUnits_39_io_casAddressOut_valid;
	wire [63:0] _networkUnits_39_io_casAddressOut_bits;
	wire _networkUnits_38_io_addressIn_ready;
	wire _networkUnits_38_io_addressOut_valid;
	wire [63:0] _networkUnits_38_io_addressOut_bits;
	wire _networkUnits_38_io_casAddressOut_valid;
	wire [63:0] _networkUnits_38_io_casAddressOut_bits;
	wire _networkUnits_37_io_addressIn_ready;
	wire _networkUnits_37_io_addressOut_valid;
	wire [63:0] _networkUnits_37_io_addressOut_bits;
	wire _networkUnits_37_io_casAddressOut_valid;
	wire [63:0] _networkUnits_37_io_casAddressOut_bits;
	wire _networkUnits_36_io_addressIn_ready;
	wire _networkUnits_36_io_addressOut_valid;
	wire [63:0] _networkUnits_36_io_addressOut_bits;
	wire _networkUnits_36_io_casAddressOut_valid;
	wire [63:0] _networkUnits_36_io_casAddressOut_bits;
	wire _networkUnits_35_io_addressIn_ready;
	wire _networkUnits_35_io_addressOut_valid;
	wire [63:0] _networkUnits_35_io_addressOut_bits;
	wire _networkUnits_35_io_casAddressOut_valid;
	wire [63:0] _networkUnits_35_io_casAddressOut_bits;
	wire _networkUnits_34_io_addressIn_ready;
	wire _networkUnits_34_io_addressOut_valid;
	wire [63:0] _networkUnits_34_io_addressOut_bits;
	wire _networkUnits_34_io_casAddressOut_valid;
	wire [63:0] _networkUnits_34_io_casAddressOut_bits;
	wire _networkUnits_33_io_addressIn_ready;
	wire _networkUnits_33_io_addressOut_valid;
	wire [63:0] _networkUnits_33_io_addressOut_bits;
	wire _networkUnits_33_io_casAddressOut_valid;
	wire [63:0] _networkUnits_33_io_casAddressOut_bits;
	wire _networkUnits_32_io_addressIn_ready;
	wire _networkUnits_32_io_addressOut_valid;
	wire [63:0] _networkUnits_32_io_addressOut_bits;
	wire _networkUnits_32_io_casAddressOut_valid;
	wire [63:0] _networkUnits_32_io_casAddressOut_bits;
	wire _networkUnits_31_io_addressIn_ready;
	wire _networkUnits_31_io_addressOut_valid;
	wire [63:0] _networkUnits_31_io_addressOut_bits;
	wire _networkUnits_31_io_casAddressOut_valid;
	wire [63:0] _networkUnits_31_io_casAddressOut_bits;
	wire _networkUnits_30_io_addressIn_ready;
	wire _networkUnits_30_io_addressOut_valid;
	wire [63:0] _networkUnits_30_io_addressOut_bits;
	wire _networkUnits_30_io_casAddressOut_valid;
	wire [63:0] _networkUnits_30_io_casAddressOut_bits;
	wire _networkUnits_29_io_addressIn_ready;
	wire _networkUnits_29_io_addressOut_valid;
	wire [63:0] _networkUnits_29_io_addressOut_bits;
	wire _networkUnits_29_io_casAddressOut_valid;
	wire [63:0] _networkUnits_29_io_casAddressOut_bits;
	wire _networkUnits_28_io_addressIn_ready;
	wire _networkUnits_28_io_addressOut_valid;
	wire [63:0] _networkUnits_28_io_addressOut_bits;
	wire _networkUnits_28_io_casAddressOut_valid;
	wire [63:0] _networkUnits_28_io_casAddressOut_bits;
	wire _networkUnits_27_io_addressIn_ready;
	wire _networkUnits_27_io_addressOut_valid;
	wire [63:0] _networkUnits_27_io_addressOut_bits;
	wire _networkUnits_27_io_casAddressOut_valid;
	wire [63:0] _networkUnits_27_io_casAddressOut_bits;
	wire _networkUnits_26_io_addressIn_ready;
	wire _networkUnits_26_io_addressOut_valid;
	wire [63:0] _networkUnits_26_io_addressOut_bits;
	wire _networkUnits_26_io_casAddressOut_valid;
	wire [63:0] _networkUnits_26_io_casAddressOut_bits;
	wire _networkUnits_25_io_addressIn_ready;
	wire _networkUnits_25_io_addressOut_valid;
	wire [63:0] _networkUnits_25_io_addressOut_bits;
	wire _networkUnits_25_io_casAddressOut_valid;
	wire [63:0] _networkUnits_25_io_casAddressOut_bits;
	wire _networkUnits_24_io_addressIn_ready;
	wire _networkUnits_24_io_addressOut_valid;
	wire [63:0] _networkUnits_24_io_addressOut_bits;
	wire _networkUnits_24_io_casAddressOut_valid;
	wire [63:0] _networkUnits_24_io_casAddressOut_bits;
	wire _networkUnits_23_io_addressIn_ready;
	wire _networkUnits_23_io_addressOut_valid;
	wire [63:0] _networkUnits_23_io_addressOut_bits;
	wire _networkUnits_23_io_casAddressOut_valid;
	wire [63:0] _networkUnits_23_io_casAddressOut_bits;
	wire _networkUnits_22_io_addressIn_ready;
	wire _networkUnits_22_io_addressOut_valid;
	wire [63:0] _networkUnits_22_io_addressOut_bits;
	wire _networkUnits_22_io_casAddressOut_valid;
	wire [63:0] _networkUnits_22_io_casAddressOut_bits;
	wire _networkUnits_21_io_addressIn_ready;
	wire _networkUnits_21_io_addressOut_valid;
	wire [63:0] _networkUnits_21_io_addressOut_bits;
	wire _networkUnits_21_io_casAddressOut_valid;
	wire [63:0] _networkUnits_21_io_casAddressOut_bits;
	wire _networkUnits_20_io_addressIn_ready;
	wire _networkUnits_20_io_addressOut_valid;
	wire [63:0] _networkUnits_20_io_addressOut_bits;
	wire _networkUnits_20_io_casAddressOut_valid;
	wire [63:0] _networkUnits_20_io_casAddressOut_bits;
	wire _networkUnits_19_io_addressIn_ready;
	wire _networkUnits_19_io_addressOut_valid;
	wire [63:0] _networkUnits_19_io_addressOut_bits;
	wire _networkUnits_19_io_casAddressOut_valid;
	wire [63:0] _networkUnits_19_io_casAddressOut_bits;
	wire _networkUnits_18_io_addressIn_ready;
	wire _networkUnits_18_io_addressOut_valid;
	wire [63:0] _networkUnits_18_io_addressOut_bits;
	wire _networkUnits_18_io_casAddressOut_valid;
	wire [63:0] _networkUnits_18_io_casAddressOut_bits;
	wire _networkUnits_17_io_addressIn_ready;
	wire _networkUnits_17_io_addressOut_valid;
	wire [63:0] _networkUnits_17_io_addressOut_bits;
	wire _networkUnits_17_io_casAddressOut_valid;
	wire [63:0] _networkUnits_17_io_casAddressOut_bits;
	wire _networkUnits_16_io_addressIn_ready;
	wire _networkUnits_16_io_addressOut_valid;
	wire [63:0] _networkUnits_16_io_addressOut_bits;
	wire _networkUnits_16_io_casAddressOut_valid;
	wire [63:0] _networkUnits_16_io_casAddressOut_bits;
	wire _networkUnits_15_io_addressIn_ready;
	wire _networkUnits_15_io_addressOut_valid;
	wire [63:0] _networkUnits_15_io_addressOut_bits;
	wire _networkUnits_15_io_casAddressOut_valid;
	wire [63:0] _networkUnits_15_io_casAddressOut_bits;
	wire _networkUnits_14_io_addressIn_ready;
	wire _networkUnits_14_io_addressOut_valid;
	wire [63:0] _networkUnits_14_io_addressOut_bits;
	wire _networkUnits_14_io_casAddressOut_valid;
	wire [63:0] _networkUnits_14_io_casAddressOut_bits;
	wire _networkUnits_13_io_addressIn_ready;
	wire _networkUnits_13_io_addressOut_valid;
	wire [63:0] _networkUnits_13_io_addressOut_bits;
	wire _networkUnits_13_io_casAddressOut_valid;
	wire [63:0] _networkUnits_13_io_casAddressOut_bits;
	wire _networkUnits_12_io_addressIn_ready;
	wire _networkUnits_12_io_addressOut_valid;
	wire [63:0] _networkUnits_12_io_addressOut_bits;
	wire _networkUnits_12_io_casAddressOut_valid;
	wire [63:0] _networkUnits_12_io_casAddressOut_bits;
	wire _networkUnits_11_io_addressIn_ready;
	wire _networkUnits_11_io_addressOut_valid;
	wire [63:0] _networkUnits_11_io_addressOut_bits;
	wire _networkUnits_11_io_casAddressOut_valid;
	wire [63:0] _networkUnits_11_io_casAddressOut_bits;
	wire _networkUnits_10_io_addressIn_ready;
	wire _networkUnits_10_io_addressOut_valid;
	wire [63:0] _networkUnits_10_io_addressOut_bits;
	wire _networkUnits_10_io_casAddressOut_valid;
	wire [63:0] _networkUnits_10_io_casAddressOut_bits;
	wire _networkUnits_9_io_addressIn_ready;
	wire _networkUnits_9_io_addressOut_valid;
	wire [63:0] _networkUnits_9_io_addressOut_bits;
	wire _networkUnits_9_io_casAddressOut_valid;
	wire [63:0] _networkUnits_9_io_casAddressOut_bits;
	wire _networkUnits_8_io_addressIn_ready;
	wire _networkUnits_8_io_addressOut_valid;
	wire [63:0] _networkUnits_8_io_addressOut_bits;
	wire _networkUnits_8_io_casAddressOut_valid;
	wire [63:0] _networkUnits_8_io_casAddressOut_bits;
	wire _networkUnits_7_io_addressIn_ready;
	wire _networkUnits_7_io_addressOut_valid;
	wire [63:0] _networkUnits_7_io_addressOut_bits;
	wire _networkUnits_7_io_casAddressOut_valid;
	wire [63:0] _networkUnits_7_io_casAddressOut_bits;
	wire _networkUnits_6_io_addressIn_ready;
	wire _networkUnits_6_io_addressOut_valid;
	wire [63:0] _networkUnits_6_io_addressOut_bits;
	wire _networkUnits_6_io_casAddressOut_valid;
	wire [63:0] _networkUnits_6_io_casAddressOut_bits;
	wire _networkUnits_5_io_addressIn_ready;
	wire _networkUnits_5_io_addressOut_valid;
	wire [63:0] _networkUnits_5_io_addressOut_bits;
	wire _networkUnits_5_io_casAddressOut_valid;
	wire [63:0] _networkUnits_5_io_casAddressOut_bits;
	wire _networkUnits_4_io_addressIn_ready;
	wire _networkUnits_4_io_addressOut_valid;
	wire [63:0] _networkUnits_4_io_addressOut_bits;
	wire _networkUnits_4_io_casAddressOut_valid;
	wire [63:0] _networkUnits_4_io_casAddressOut_bits;
	wire _networkUnits_3_io_addressIn_ready;
	wire _networkUnits_3_io_addressOut_valid;
	wire [63:0] _networkUnits_3_io_addressOut_bits;
	wire _networkUnits_3_io_casAddressOut_valid;
	wire [63:0] _networkUnits_3_io_casAddressOut_bits;
	wire _networkUnits_2_io_addressIn_ready;
	wire _networkUnits_2_io_addressOut_valid;
	wire [63:0] _networkUnits_2_io_addressOut_bits;
	wire _networkUnits_2_io_casAddressOut_valid;
	wire [63:0] _networkUnits_2_io_casAddressOut_bits;
	wire _networkUnits_1_io_addressIn_ready;
	wire _networkUnits_1_io_addressOut_valid;
	wire [63:0] _networkUnits_1_io_addressOut_bits;
	wire _networkUnits_1_io_casAddressOut_valid;
	wire [63:0] _networkUnits_1_io_casAddressOut_bits;
	wire _networkUnits_0_io_addressIn_ready;
	wire _networkUnits_0_io_addressOut_valid;
	wire [63:0] _networkUnits_0_io_addressOut_bits;
	wire _networkUnits_0_io_casAddressOut_valid;
	wire [63:0] _networkUnits_0_io_casAddressOut_bits;
	wire _vcasNetworkUnits_3_io_addressIn0_ready;
	wire _vcasNetworkUnits_3_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_3_io_addressOut_bits;
	wire _vcasNetworkUnits_2_io_addressIn0_ready;
	wire _vcasNetworkUnits_2_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_2_io_addressOut_bits;
	wire _vcasNetworkUnits_1_io_addressIn0_ready;
	wire _vcasNetworkUnits_1_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_1_io_addressOut_bits;
	wire _vcasNetworkUnits_0_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_0_io_addressOut_bits;
	AllocatorServerNetworkUnit vcasNetworkUnits_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(),
		.io_addressIn0_valid(1'h0),
		.io_addressIn0_bits(64'h0000000000000000),
		.io_addressIn1_ready(io_connVCAS_0_ready),
		.io_addressIn1_valid(io_connVCAS_0_valid),
		.io_addressIn1_bits(io_connVCAS_0_bits),
		.io_addressOut_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_0_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_0_io_addressOut_bits)
	);
	AllocatorServerNetworkUnit vcasNetworkUnits_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(_vcasNetworkUnits_1_io_addressIn0_ready),
		.io_addressIn0_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressIn0_bits(_networkUnits_15_io_addressOut_bits),
		.io_addressIn1_ready(io_connVCAS_1_ready),
		.io_addressIn1_valid(io_connVCAS_1_valid),
		.io_addressIn1_bits(io_connVCAS_1_bits),
		.io_addressOut_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_1_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_1_io_addressOut_bits)
	);
	AllocatorServerNetworkUnit vcasNetworkUnits_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(_vcasNetworkUnits_2_io_addressIn0_ready),
		.io_addressIn0_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressIn0_bits(_networkUnits_31_io_addressOut_bits),
		.io_addressIn1_ready(io_connVCAS_2_ready),
		.io_addressIn1_valid(io_connVCAS_2_valid),
		.io_addressIn1_bits(io_connVCAS_2_bits),
		.io_addressOut_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_2_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_2_io_addressOut_bits)
	);
	AllocatorServerNetworkUnit vcasNetworkUnits_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(_vcasNetworkUnits_3_io_addressIn0_ready),
		.io_addressIn0_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressIn0_bits(_networkUnits_47_io_addressOut_bits),
		.io_addressIn1_ready(io_connVCAS_3_ready),
		.io_addressIn1_valid(io_connVCAS_3_valid),
		.io_addressIn1_bits(io_connVCAS_3_bits),
		.io_addressOut_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_3_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_3_io_addressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_0_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_0_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_0_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_0_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_0_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_0_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_0_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_1_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_1_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_1_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_1_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_1_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_2_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_2_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_2_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_2_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_2_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_3_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_3_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_3_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_3_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_3_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_4_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_4_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_4_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_4_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_4_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_5_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_5_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_5_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_5_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_5_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_6_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_6_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_6_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_6_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_6_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_7_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_7_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_7_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_7_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_7_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_8_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_8_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_8_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_8_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_8_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_9_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_9_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_9_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_9_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_9_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_10_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_10_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_10_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_10_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_10_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_11_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_11_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_11_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_11_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_11_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_12_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_12_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_12_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_12_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_12_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_13_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_13_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_13_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_13_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_13_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_14_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_14_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_14_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_14_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_14_io_addressOut_bits),
		.io_addressOut_ready(_vcasNetworkUnits_1_io_addressIn0_ready),
		.io_addressOut_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_15_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_15_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_15_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_15_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_1_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_1_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_16_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_16_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_16_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_16_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_16_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_17_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_17_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_17_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_17_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_17_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_18_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_18_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_18_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_18_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_18_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_19_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_19_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_19_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_19_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_19_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_20_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_20_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_20_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_20_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_20_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_21_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_21_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_21_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_21_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_21_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_22_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_22_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_22_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_22_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_22_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_23_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_23_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_23_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_23_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_23_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_24_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_24_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_24_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_24_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_24_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_25_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_25_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_25_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_25_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_25_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_26_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_26_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_26_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_26_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_26_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_27_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_27_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_27_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_27_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_27_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_28_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_28_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_28_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_28_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_28_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_29_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_29_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_29_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_29_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_29_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_30_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_30_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_30_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_30_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_30_io_addressOut_bits),
		.io_addressOut_ready(_vcasNetworkUnits_2_io_addressIn0_ready),
		.io_addressOut_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_31_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_31_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_31_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_31_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_2_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_2_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_32_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_32_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_32_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_32_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_32_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_33_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_33_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_33_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_33_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_33_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_34_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_34_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_34_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_34_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_34_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_35_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_35_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_35_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_35_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_35_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_36_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_36_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_36_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_36_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_36_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_37_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_37_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_37_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_37_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_37_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_38_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_38_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_38_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_38_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_38_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_39_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_39_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_39_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_39_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_39_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_40_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_40_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_40_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_40_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_40_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_41_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_41_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_41_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_41_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_41_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_42_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_42_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_42_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_42_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_42_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_43_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_43_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_43_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_43_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_43_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_44_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_44_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_44_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_44_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_44_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_45_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_45_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_45_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_45_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_45_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_46_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_46_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_46_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_46_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_46_io_addressOut_bits),
		.io_addressOut_ready(_vcasNetworkUnits_3_io_addressIn0_ready),
		.io_addressOut_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_47_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_47_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_47_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_47_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_3_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_3_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_48_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_48_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_48_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_48_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_48_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_49_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_49_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_49_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_49_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_49_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_50_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_50_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_50_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_50_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_50_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_51_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_51_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_51_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_51_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_51_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_52_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_52_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_52_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_52_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_52_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_53_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_53_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_53_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_53_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_53_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_54_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_54_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_54_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_54_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_54_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_55_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_55_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_55_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_55_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_55_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_56_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_56_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_56_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_56_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_56_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_57_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_57_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_57_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_57_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_57_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_58_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_58_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_58_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_58_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_58_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_59_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_59_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_59_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_59_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_59_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_60_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_60_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_60_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_60_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_60_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_61_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_61_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_61_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_61_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_61_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_62_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_62_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_62_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_62_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_62_io_addressOut_bits),
		.io_addressOut_ready(1'h0),
		.io_addressOut_valid(),
		.io_addressOut_bits(),
		.io_casAddressOut_ready(_casServers_63_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_63_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_63_io_casAddressOut_bits)
	);
	AllocatorClient casServers_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_0_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_0_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_0_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_0_io_addressIn_ready),
		.io_addressOut_valid(_casServers_0_io_addressOut_valid),
		.io_addressOut_bits(_casServers_0_io_addressOut_bits)
	);
	AllocatorClient casServers_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_1_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_1_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_1_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_1_io_addressIn_ready),
		.io_addressOut_valid(_casServers_1_io_addressOut_valid),
		.io_addressOut_bits(_casServers_1_io_addressOut_bits)
	);
	AllocatorClient casServers_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_2_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_2_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_2_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_2_io_addressIn_ready),
		.io_addressOut_valid(_casServers_2_io_addressOut_valid),
		.io_addressOut_bits(_casServers_2_io_addressOut_bits)
	);
	AllocatorClient casServers_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_3_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_3_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_3_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_3_io_addressIn_ready),
		.io_addressOut_valid(_casServers_3_io_addressOut_valid),
		.io_addressOut_bits(_casServers_3_io_addressOut_bits)
	);
	AllocatorClient casServers_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_4_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_4_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_4_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_4_io_addressIn_ready),
		.io_addressOut_valid(_casServers_4_io_addressOut_valid),
		.io_addressOut_bits(_casServers_4_io_addressOut_bits)
	);
	AllocatorClient casServers_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_5_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_5_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_5_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_5_io_addressIn_ready),
		.io_addressOut_valid(_casServers_5_io_addressOut_valid),
		.io_addressOut_bits(_casServers_5_io_addressOut_bits)
	);
	AllocatorClient casServers_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_6_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_6_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_6_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_6_io_addressIn_ready),
		.io_addressOut_valid(_casServers_6_io_addressOut_valid),
		.io_addressOut_bits(_casServers_6_io_addressOut_bits)
	);
	AllocatorClient casServers_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_7_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_7_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_7_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_7_io_addressIn_ready),
		.io_addressOut_valid(_casServers_7_io_addressOut_valid),
		.io_addressOut_bits(_casServers_7_io_addressOut_bits)
	);
	AllocatorClient casServers_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_8_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_8_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_8_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_8_io_addressIn_ready),
		.io_addressOut_valid(_casServers_8_io_addressOut_valid),
		.io_addressOut_bits(_casServers_8_io_addressOut_bits)
	);
	AllocatorClient casServers_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_9_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_9_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_9_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_9_io_addressIn_ready),
		.io_addressOut_valid(_casServers_9_io_addressOut_valid),
		.io_addressOut_bits(_casServers_9_io_addressOut_bits)
	);
	AllocatorClient casServers_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_10_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_10_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_10_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_10_io_addressIn_ready),
		.io_addressOut_valid(_casServers_10_io_addressOut_valid),
		.io_addressOut_bits(_casServers_10_io_addressOut_bits)
	);
	AllocatorClient casServers_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_11_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_11_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_11_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_11_io_addressIn_ready),
		.io_addressOut_valid(_casServers_11_io_addressOut_valid),
		.io_addressOut_bits(_casServers_11_io_addressOut_bits)
	);
	AllocatorClient casServers_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_12_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_12_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_12_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_12_io_addressIn_ready),
		.io_addressOut_valid(_casServers_12_io_addressOut_valid),
		.io_addressOut_bits(_casServers_12_io_addressOut_bits)
	);
	AllocatorClient casServers_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_13_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_13_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_13_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_13_io_addressIn_ready),
		.io_addressOut_valid(_casServers_13_io_addressOut_valid),
		.io_addressOut_bits(_casServers_13_io_addressOut_bits)
	);
	AllocatorClient casServers_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_14_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_14_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_14_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_14_io_addressIn_ready),
		.io_addressOut_valid(_casServers_14_io_addressOut_valid),
		.io_addressOut_bits(_casServers_14_io_addressOut_bits)
	);
	AllocatorClient casServers_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_15_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_15_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_15_io_addressIn_ready),
		.io_addressOut_valid(_casServers_15_io_addressOut_valid),
		.io_addressOut_bits(_casServers_15_io_addressOut_bits)
	);
	AllocatorClient casServers_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_16_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_16_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_16_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_16_io_addressIn_ready),
		.io_addressOut_valid(_casServers_16_io_addressOut_valid),
		.io_addressOut_bits(_casServers_16_io_addressOut_bits)
	);
	AllocatorClient casServers_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_17_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_17_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_17_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_17_io_addressIn_ready),
		.io_addressOut_valid(_casServers_17_io_addressOut_valid),
		.io_addressOut_bits(_casServers_17_io_addressOut_bits)
	);
	AllocatorClient casServers_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_18_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_18_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_18_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_18_io_addressIn_ready),
		.io_addressOut_valid(_casServers_18_io_addressOut_valid),
		.io_addressOut_bits(_casServers_18_io_addressOut_bits)
	);
	AllocatorClient casServers_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_19_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_19_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_19_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_19_io_addressIn_ready),
		.io_addressOut_valid(_casServers_19_io_addressOut_valid),
		.io_addressOut_bits(_casServers_19_io_addressOut_bits)
	);
	AllocatorClient casServers_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_20_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_20_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_20_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_20_io_addressIn_ready),
		.io_addressOut_valid(_casServers_20_io_addressOut_valid),
		.io_addressOut_bits(_casServers_20_io_addressOut_bits)
	);
	AllocatorClient casServers_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_21_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_21_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_21_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_21_io_addressIn_ready),
		.io_addressOut_valid(_casServers_21_io_addressOut_valid),
		.io_addressOut_bits(_casServers_21_io_addressOut_bits)
	);
	AllocatorClient casServers_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_22_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_22_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_22_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_22_io_addressIn_ready),
		.io_addressOut_valid(_casServers_22_io_addressOut_valid),
		.io_addressOut_bits(_casServers_22_io_addressOut_bits)
	);
	AllocatorClient casServers_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_23_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_23_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_23_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_23_io_addressIn_ready),
		.io_addressOut_valid(_casServers_23_io_addressOut_valid),
		.io_addressOut_bits(_casServers_23_io_addressOut_bits)
	);
	AllocatorClient casServers_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_24_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_24_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_24_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_24_io_addressIn_ready),
		.io_addressOut_valid(_casServers_24_io_addressOut_valid),
		.io_addressOut_bits(_casServers_24_io_addressOut_bits)
	);
	AllocatorClient casServers_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_25_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_25_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_25_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_25_io_addressIn_ready),
		.io_addressOut_valid(_casServers_25_io_addressOut_valid),
		.io_addressOut_bits(_casServers_25_io_addressOut_bits)
	);
	AllocatorClient casServers_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_26_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_26_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_26_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_26_io_addressIn_ready),
		.io_addressOut_valid(_casServers_26_io_addressOut_valid),
		.io_addressOut_bits(_casServers_26_io_addressOut_bits)
	);
	AllocatorClient casServers_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_27_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_27_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_27_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_27_io_addressIn_ready),
		.io_addressOut_valid(_casServers_27_io_addressOut_valid),
		.io_addressOut_bits(_casServers_27_io_addressOut_bits)
	);
	AllocatorClient casServers_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_28_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_28_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_28_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_28_io_addressIn_ready),
		.io_addressOut_valid(_casServers_28_io_addressOut_valid),
		.io_addressOut_bits(_casServers_28_io_addressOut_bits)
	);
	AllocatorClient casServers_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_29_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_29_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_29_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_29_io_addressIn_ready),
		.io_addressOut_valid(_casServers_29_io_addressOut_valid),
		.io_addressOut_bits(_casServers_29_io_addressOut_bits)
	);
	AllocatorClient casServers_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_30_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_30_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_30_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_30_io_addressIn_ready),
		.io_addressOut_valid(_casServers_30_io_addressOut_valid),
		.io_addressOut_bits(_casServers_30_io_addressOut_bits)
	);
	AllocatorClient casServers_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_31_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_31_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_31_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_31_io_addressIn_ready),
		.io_addressOut_valid(_casServers_31_io_addressOut_valid),
		.io_addressOut_bits(_casServers_31_io_addressOut_bits)
	);
	AllocatorClient casServers_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_32_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_32_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_32_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_32_io_addressIn_ready),
		.io_addressOut_valid(_casServers_32_io_addressOut_valid),
		.io_addressOut_bits(_casServers_32_io_addressOut_bits)
	);
	AllocatorClient casServers_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_33_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_33_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_33_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_33_io_addressIn_ready),
		.io_addressOut_valid(_casServers_33_io_addressOut_valid),
		.io_addressOut_bits(_casServers_33_io_addressOut_bits)
	);
	AllocatorClient casServers_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_34_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_34_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_34_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_34_io_addressIn_ready),
		.io_addressOut_valid(_casServers_34_io_addressOut_valid),
		.io_addressOut_bits(_casServers_34_io_addressOut_bits)
	);
	AllocatorClient casServers_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_35_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_35_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_35_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_35_io_addressIn_ready),
		.io_addressOut_valid(_casServers_35_io_addressOut_valid),
		.io_addressOut_bits(_casServers_35_io_addressOut_bits)
	);
	AllocatorClient casServers_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_36_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_36_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_36_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_36_io_addressIn_ready),
		.io_addressOut_valid(_casServers_36_io_addressOut_valid),
		.io_addressOut_bits(_casServers_36_io_addressOut_bits)
	);
	AllocatorClient casServers_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_37_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_37_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_37_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_37_io_addressIn_ready),
		.io_addressOut_valid(_casServers_37_io_addressOut_valid),
		.io_addressOut_bits(_casServers_37_io_addressOut_bits)
	);
	AllocatorClient casServers_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_38_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_38_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_38_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_38_io_addressIn_ready),
		.io_addressOut_valid(_casServers_38_io_addressOut_valid),
		.io_addressOut_bits(_casServers_38_io_addressOut_bits)
	);
	AllocatorClient casServers_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_39_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_39_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_39_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_39_io_addressIn_ready),
		.io_addressOut_valid(_casServers_39_io_addressOut_valid),
		.io_addressOut_bits(_casServers_39_io_addressOut_bits)
	);
	AllocatorClient casServers_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_40_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_40_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_40_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_40_io_addressIn_ready),
		.io_addressOut_valid(_casServers_40_io_addressOut_valid),
		.io_addressOut_bits(_casServers_40_io_addressOut_bits)
	);
	AllocatorClient casServers_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_41_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_41_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_41_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_41_io_addressIn_ready),
		.io_addressOut_valid(_casServers_41_io_addressOut_valid),
		.io_addressOut_bits(_casServers_41_io_addressOut_bits)
	);
	AllocatorClient casServers_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_42_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_42_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_42_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_42_io_addressIn_ready),
		.io_addressOut_valid(_casServers_42_io_addressOut_valid),
		.io_addressOut_bits(_casServers_42_io_addressOut_bits)
	);
	AllocatorClient casServers_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_43_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_43_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_43_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_43_io_addressIn_ready),
		.io_addressOut_valid(_casServers_43_io_addressOut_valid),
		.io_addressOut_bits(_casServers_43_io_addressOut_bits)
	);
	AllocatorClient casServers_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_44_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_44_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_44_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_44_io_addressIn_ready),
		.io_addressOut_valid(_casServers_44_io_addressOut_valid),
		.io_addressOut_bits(_casServers_44_io_addressOut_bits)
	);
	AllocatorClient casServers_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_45_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_45_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_45_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_45_io_addressIn_ready),
		.io_addressOut_valid(_casServers_45_io_addressOut_valid),
		.io_addressOut_bits(_casServers_45_io_addressOut_bits)
	);
	AllocatorClient casServers_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_46_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_46_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_46_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_46_io_addressIn_ready),
		.io_addressOut_valid(_casServers_46_io_addressOut_valid),
		.io_addressOut_bits(_casServers_46_io_addressOut_bits)
	);
	AllocatorClient casServers_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_47_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_47_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_47_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_47_io_addressIn_ready),
		.io_addressOut_valid(_casServers_47_io_addressOut_valid),
		.io_addressOut_bits(_casServers_47_io_addressOut_bits)
	);
	AllocatorClient casServers_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_48_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_48_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_48_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_48_io_addressIn_ready),
		.io_addressOut_valid(_casServers_48_io_addressOut_valid),
		.io_addressOut_bits(_casServers_48_io_addressOut_bits)
	);
	AllocatorClient casServers_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_49_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_49_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_49_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_49_io_addressIn_ready),
		.io_addressOut_valid(_casServers_49_io_addressOut_valid),
		.io_addressOut_bits(_casServers_49_io_addressOut_bits)
	);
	AllocatorClient casServers_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_50_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_50_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_50_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_50_io_addressIn_ready),
		.io_addressOut_valid(_casServers_50_io_addressOut_valid),
		.io_addressOut_bits(_casServers_50_io_addressOut_bits)
	);
	AllocatorClient casServers_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_51_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_51_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_51_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_51_io_addressIn_ready),
		.io_addressOut_valid(_casServers_51_io_addressOut_valid),
		.io_addressOut_bits(_casServers_51_io_addressOut_bits)
	);
	AllocatorClient casServers_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_52_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_52_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_52_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_52_io_addressIn_ready),
		.io_addressOut_valid(_casServers_52_io_addressOut_valid),
		.io_addressOut_bits(_casServers_52_io_addressOut_bits)
	);
	AllocatorClient casServers_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_53_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_53_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_53_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_53_io_addressIn_ready),
		.io_addressOut_valid(_casServers_53_io_addressOut_valid),
		.io_addressOut_bits(_casServers_53_io_addressOut_bits)
	);
	AllocatorClient casServers_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_54_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_54_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_54_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_54_io_addressIn_ready),
		.io_addressOut_valid(_casServers_54_io_addressOut_valid),
		.io_addressOut_bits(_casServers_54_io_addressOut_bits)
	);
	AllocatorClient casServers_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_55_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_55_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_55_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_55_io_addressIn_ready),
		.io_addressOut_valid(_casServers_55_io_addressOut_valid),
		.io_addressOut_bits(_casServers_55_io_addressOut_bits)
	);
	AllocatorClient casServers_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_56_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_56_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_56_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_56_io_addressIn_ready),
		.io_addressOut_valid(_casServers_56_io_addressOut_valid),
		.io_addressOut_bits(_casServers_56_io_addressOut_bits)
	);
	AllocatorClient casServers_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_57_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_57_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_57_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_57_io_addressIn_ready),
		.io_addressOut_valid(_casServers_57_io_addressOut_valid),
		.io_addressOut_bits(_casServers_57_io_addressOut_bits)
	);
	AllocatorClient casServers_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_58_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_58_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_58_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_58_io_addressIn_ready),
		.io_addressOut_valid(_casServers_58_io_addressOut_valid),
		.io_addressOut_bits(_casServers_58_io_addressOut_bits)
	);
	AllocatorClient casServers_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_59_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_59_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_59_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_59_io_addressIn_ready),
		.io_addressOut_valid(_casServers_59_io_addressOut_valid),
		.io_addressOut_bits(_casServers_59_io_addressOut_bits)
	);
	AllocatorClient casServers_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_60_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_60_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_60_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_60_io_addressIn_ready),
		.io_addressOut_valid(_casServers_60_io_addressOut_valid),
		.io_addressOut_bits(_casServers_60_io_addressOut_bits)
	);
	AllocatorClient casServers_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_61_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_61_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_61_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_61_io_addressIn_ready),
		.io_addressOut_valid(_casServers_61_io_addressOut_valid),
		.io_addressOut_bits(_casServers_61_io_addressOut_bits)
	);
	AllocatorClient casServers_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_62_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_62_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_62_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_62_io_addressIn_ready),
		.io_addressOut_valid(_casServers_62_io_addressOut_valid),
		.io_addressOut_bits(_casServers_62_io_addressOut_bits)
	);
	AllocatorClient casServers_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_63_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_63_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_63_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_63_io_addressIn_ready),
		.io_addressOut_valid(_casServers_63_io_addressOut_valid),
		.io_addressOut_bits(_casServers_63_io_addressOut_bits)
	);
	AllocatorBuffer queues_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_0_io_addressIn_ready),
		.io_addressIn_valid(_casServers_0_io_addressOut_valid),
		.io_addressIn_bits(_casServers_0_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_0_ready),
		.io_addressOut_valid(io_connPE_0_valid),
		.io_addressOut_bits(io_connPE_0_bits)
	);
	AllocatorBuffer queues_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_1_io_addressIn_ready),
		.io_addressIn_valid(_casServers_1_io_addressOut_valid),
		.io_addressIn_bits(_casServers_1_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_1_ready),
		.io_addressOut_valid(io_connPE_1_valid),
		.io_addressOut_bits(io_connPE_1_bits)
	);
	AllocatorBuffer queues_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_2_io_addressIn_ready),
		.io_addressIn_valid(_casServers_2_io_addressOut_valid),
		.io_addressIn_bits(_casServers_2_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_2_ready),
		.io_addressOut_valid(io_connPE_2_valid),
		.io_addressOut_bits(io_connPE_2_bits)
	);
	AllocatorBuffer queues_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_3_io_addressIn_ready),
		.io_addressIn_valid(_casServers_3_io_addressOut_valid),
		.io_addressIn_bits(_casServers_3_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_3_ready),
		.io_addressOut_valid(io_connPE_3_valid),
		.io_addressOut_bits(io_connPE_3_bits)
	);
	AllocatorBuffer queues_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_4_io_addressIn_ready),
		.io_addressIn_valid(_casServers_4_io_addressOut_valid),
		.io_addressIn_bits(_casServers_4_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_4_ready),
		.io_addressOut_valid(io_connPE_4_valid),
		.io_addressOut_bits(io_connPE_4_bits)
	);
	AllocatorBuffer queues_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_5_io_addressIn_ready),
		.io_addressIn_valid(_casServers_5_io_addressOut_valid),
		.io_addressIn_bits(_casServers_5_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_5_ready),
		.io_addressOut_valid(io_connPE_5_valid),
		.io_addressOut_bits(io_connPE_5_bits)
	);
	AllocatorBuffer queues_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_6_io_addressIn_ready),
		.io_addressIn_valid(_casServers_6_io_addressOut_valid),
		.io_addressIn_bits(_casServers_6_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_6_ready),
		.io_addressOut_valid(io_connPE_6_valid),
		.io_addressOut_bits(io_connPE_6_bits)
	);
	AllocatorBuffer queues_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_7_io_addressIn_ready),
		.io_addressIn_valid(_casServers_7_io_addressOut_valid),
		.io_addressIn_bits(_casServers_7_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_7_ready),
		.io_addressOut_valid(io_connPE_7_valid),
		.io_addressOut_bits(io_connPE_7_bits)
	);
	AllocatorBuffer queues_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_8_io_addressIn_ready),
		.io_addressIn_valid(_casServers_8_io_addressOut_valid),
		.io_addressIn_bits(_casServers_8_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_8_ready),
		.io_addressOut_valid(io_connPE_8_valid),
		.io_addressOut_bits(io_connPE_8_bits)
	);
	AllocatorBuffer queues_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_9_io_addressIn_ready),
		.io_addressIn_valid(_casServers_9_io_addressOut_valid),
		.io_addressIn_bits(_casServers_9_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_9_ready),
		.io_addressOut_valid(io_connPE_9_valid),
		.io_addressOut_bits(io_connPE_9_bits)
	);
	AllocatorBuffer queues_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_10_io_addressIn_ready),
		.io_addressIn_valid(_casServers_10_io_addressOut_valid),
		.io_addressIn_bits(_casServers_10_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_10_ready),
		.io_addressOut_valid(io_connPE_10_valid),
		.io_addressOut_bits(io_connPE_10_bits)
	);
	AllocatorBuffer queues_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_11_io_addressIn_ready),
		.io_addressIn_valid(_casServers_11_io_addressOut_valid),
		.io_addressIn_bits(_casServers_11_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_11_ready),
		.io_addressOut_valid(io_connPE_11_valid),
		.io_addressOut_bits(io_connPE_11_bits)
	);
	AllocatorBuffer queues_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_12_io_addressIn_ready),
		.io_addressIn_valid(_casServers_12_io_addressOut_valid),
		.io_addressIn_bits(_casServers_12_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_12_ready),
		.io_addressOut_valid(io_connPE_12_valid),
		.io_addressOut_bits(io_connPE_12_bits)
	);
	AllocatorBuffer queues_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_13_io_addressIn_ready),
		.io_addressIn_valid(_casServers_13_io_addressOut_valid),
		.io_addressIn_bits(_casServers_13_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_13_ready),
		.io_addressOut_valid(io_connPE_13_valid),
		.io_addressOut_bits(io_connPE_13_bits)
	);
	AllocatorBuffer queues_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_14_io_addressIn_ready),
		.io_addressIn_valid(_casServers_14_io_addressOut_valid),
		.io_addressIn_bits(_casServers_14_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_14_ready),
		.io_addressOut_valid(io_connPE_14_valid),
		.io_addressOut_bits(io_connPE_14_bits)
	);
	AllocatorBuffer queues_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_15_io_addressIn_ready),
		.io_addressIn_valid(_casServers_15_io_addressOut_valid),
		.io_addressIn_bits(_casServers_15_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_15_ready),
		.io_addressOut_valid(io_connPE_15_valid),
		.io_addressOut_bits(io_connPE_15_bits)
	);
	AllocatorBuffer queues_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_16_io_addressIn_ready),
		.io_addressIn_valid(_casServers_16_io_addressOut_valid),
		.io_addressIn_bits(_casServers_16_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_16_ready),
		.io_addressOut_valid(io_connPE_16_valid),
		.io_addressOut_bits(io_connPE_16_bits)
	);
	AllocatorBuffer queues_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_17_io_addressIn_ready),
		.io_addressIn_valid(_casServers_17_io_addressOut_valid),
		.io_addressIn_bits(_casServers_17_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_17_ready),
		.io_addressOut_valid(io_connPE_17_valid),
		.io_addressOut_bits(io_connPE_17_bits)
	);
	AllocatorBuffer queues_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_18_io_addressIn_ready),
		.io_addressIn_valid(_casServers_18_io_addressOut_valid),
		.io_addressIn_bits(_casServers_18_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_18_ready),
		.io_addressOut_valid(io_connPE_18_valid),
		.io_addressOut_bits(io_connPE_18_bits)
	);
	AllocatorBuffer queues_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_19_io_addressIn_ready),
		.io_addressIn_valid(_casServers_19_io_addressOut_valid),
		.io_addressIn_bits(_casServers_19_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_19_ready),
		.io_addressOut_valid(io_connPE_19_valid),
		.io_addressOut_bits(io_connPE_19_bits)
	);
	AllocatorBuffer queues_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_20_io_addressIn_ready),
		.io_addressIn_valid(_casServers_20_io_addressOut_valid),
		.io_addressIn_bits(_casServers_20_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_20_ready),
		.io_addressOut_valid(io_connPE_20_valid),
		.io_addressOut_bits(io_connPE_20_bits)
	);
	AllocatorBuffer queues_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_21_io_addressIn_ready),
		.io_addressIn_valid(_casServers_21_io_addressOut_valid),
		.io_addressIn_bits(_casServers_21_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_21_ready),
		.io_addressOut_valid(io_connPE_21_valid),
		.io_addressOut_bits(io_connPE_21_bits)
	);
	AllocatorBuffer queues_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_22_io_addressIn_ready),
		.io_addressIn_valid(_casServers_22_io_addressOut_valid),
		.io_addressIn_bits(_casServers_22_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_22_ready),
		.io_addressOut_valid(io_connPE_22_valid),
		.io_addressOut_bits(io_connPE_22_bits)
	);
	AllocatorBuffer queues_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_23_io_addressIn_ready),
		.io_addressIn_valid(_casServers_23_io_addressOut_valid),
		.io_addressIn_bits(_casServers_23_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_23_ready),
		.io_addressOut_valid(io_connPE_23_valid),
		.io_addressOut_bits(io_connPE_23_bits)
	);
	AllocatorBuffer queues_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_24_io_addressIn_ready),
		.io_addressIn_valid(_casServers_24_io_addressOut_valid),
		.io_addressIn_bits(_casServers_24_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_24_ready),
		.io_addressOut_valid(io_connPE_24_valid),
		.io_addressOut_bits(io_connPE_24_bits)
	);
	AllocatorBuffer queues_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_25_io_addressIn_ready),
		.io_addressIn_valid(_casServers_25_io_addressOut_valid),
		.io_addressIn_bits(_casServers_25_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_25_ready),
		.io_addressOut_valid(io_connPE_25_valid),
		.io_addressOut_bits(io_connPE_25_bits)
	);
	AllocatorBuffer queues_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_26_io_addressIn_ready),
		.io_addressIn_valid(_casServers_26_io_addressOut_valid),
		.io_addressIn_bits(_casServers_26_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_26_ready),
		.io_addressOut_valid(io_connPE_26_valid),
		.io_addressOut_bits(io_connPE_26_bits)
	);
	AllocatorBuffer queues_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_27_io_addressIn_ready),
		.io_addressIn_valid(_casServers_27_io_addressOut_valid),
		.io_addressIn_bits(_casServers_27_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_27_ready),
		.io_addressOut_valid(io_connPE_27_valid),
		.io_addressOut_bits(io_connPE_27_bits)
	);
	AllocatorBuffer queues_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_28_io_addressIn_ready),
		.io_addressIn_valid(_casServers_28_io_addressOut_valid),
		.io_addressIn_bits(_casServers_28_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_28_ready),
		.io_addressOut_valid(io_connPE_28_valid),
		.io_addressOut_bits(io_connPE_28_bits)
	);
	AllocatorBuffer queues_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_29_io_addressIn_ready),
		.io_addressIn_valid(_casServers_29_io_addressOut_valid),
		.io_addressIn_bits(_casServers_29_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_29_ready),
		.io_addressOut_valid(io_connPE_29_valid),
		.io_addressOut_bits(io_connPE_29_bits)
	);
	AllocatorBuffer queues_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_30_io_addressIn_ready),
		.io_addressIn_valid(_casServers_30_io_addressOut_valid),
		.io_addressIn_bits(_casServers_30_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_30_ready),
		.io_addressOut_valid(io_connPE_30_valid),
		.io_addressOut_bits(io_connPE_30_bits)
	);
	AllocatorBuffer queues_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_31_io_addressIn_ready),
		.io_addressIn_valid(_casServers_31_io_addressOut_valid),
		.io_addressIn_bits(_casServers_31_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_31_ready),
		.io_addressOut_valid(io_connPE_31_valid),
		.io_addressOut_bits(io_connPE_31_bits)
	);
	AllocatorBuffer queues_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_32_io_addressIn_ready),
		.io_addressIn_valid(_casServers_32_io_addressOut_valid),
		.io_addressIn_bits(_casServers_32_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_32_ready),
		.io_addressOut_valid(io_connPE_32_valid),
		.io_addressOut_bits(io_connPE_32_bits)
	);
	AllocatorBuffer queues_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_33_io_addressIn_ready),
		.io_addressIn_valid(_casServers_33_io_addressOut_valid),
		.io_addressIn_bits(_casServers_33_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_33_ready),
		.io_addressOut_valid(io_connPE_33_valid),
		.io_addressOut_bits(io_connPE_33_bits)
	);
	AllocatorBuffer queues_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_34_io_addressIn_ready),
		.io_addressIn_valid(_casServers_34_io_addressOut_valid),
		.io_addressIn_bits(_casServers_34_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_34_ready),
		.io_addressOut_valid(io_connPE_34_valid),
		.io_addressOut_bits(io_connPE_34_bits)
	);
	AllocatorBuffer queues_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_35_io_addressIn_ready),
		.io_addressIn_valid(_casServers_35_io_addressOut_valid),
		.io_addressIn_bits(_casServers_35_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_35_ready),
		.io_addressOut_valid(io_connPE_35_valid),
		.io_addressOut_bits(io_connPE_35_bits)
	);
	AllocatorBuffer queues_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_36_io_addressIn_ready),
		.io_addressIn_valid(_casServers_36_io_addressOut_valid),
		.io_addressIn_bits(_casServers_36_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_36_ready),
		.io_addressOut_valid(io_connPE_36_valid),
		.io_addressOut_bits(io_connPE_36_bits)
	);
	AllocatorBuffer queues_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_37_io_addressIn_ready),
		.io_addressIn_valid(_casServers_37_io_addressOut_valid),
		.io_addressIn_bits(_casServers_37_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_37_ready),
		.io_addressOut_valid(io_connPE_37_valid),
		.io_addressOut_bits(io_connPE_37_bits)
	);
	AllocatorBuffer queues_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_38_io_addressIn_ready),
		.io_addressIn_valid(_casServers_38_io_addressOut_valid),
		.io_addressIn_bits(_casServers_38_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_38_ready),
		.io_addressOut_valid(io_connPE_38_valid),
		.io_addressOut_bits(io_connPE_38_bits)
	);
	AllocatorBuffer queues_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_39_io_addressIn_ready),
		.io_addressIn_valid(_casServers_39_io_addressOut_valid),
		.io_addressIn_bits(_casServers_39_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_39_ready),
		.io_addressOut_valid(io_connPE_39_valid),
		.io_addressOut_bits(io_connPE_39_bits)
	);
	AllocatorBuffer queues_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_40_io_addressIn_ready),
		.io_addressIn_valid(_casServers_40_io_addressOut_valid),
		.io_addressIn_bits(_casServers_40_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_40_ready),
		.io_addressOut_valid(io_connPE_40_valid),
		.io_addressOut_bits(io_connPE_40_bits)
	);
	AllocatorBuffer queues_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_41_io_addressIn_ready),
		.io_addressIn_valid(_casServers_41_io_addressOut_valid),
		.io_addressIn_bits(_casServers_41_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_41_ready),
		.io_addressOut_valid(io_connPE_41_valid),
		.io_addressOut_bits(io_connPE_41_bits)
	);
	AllocatorBuffer queues_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_42_io_addressIn_ready),
		.io_addressIn_valid(_casServers_42_io_addressOut_valid),
		.io_addressIn_bits(_casServers_42_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_42_ready),
		.io_addressOut_valid(io_connPE_42_valid),
		.io_addressOut_bits(io_connPE_42_bits)
	);
	AllocatorBuffer queues_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_43_io_addressIn_ready),
		.io_addressIn_valid(_casServers_43_io_addressOut_valid),
		.io_addressIn_bits(_casServers_43_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_43_ready),
		.io_addressOut_valid(io_connPE_43_valid),
		.io_addressOut_bits(io_connPE_43_bits)
	);
	AllocatorBuffer queues_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_44_io_addressIn_ready),
		.io_addressIn_valid(_casServers_44_io_addressOut_valid),
		.io_addressIn_bits(_casServers_44_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_44_ready),
		.io_addressOut_valid(io_connPE_44_valid),
		.io_addressOut_bits(io_connPE_44_bits)
	);
	AllocatorBuffer queues_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_45_io_addressIn_ready),
		.io_addressIn_valid(_casServers_45_io_addressOut_valid),
		.io_addressIn_bits(_casServers_45_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_45_ready),
		.io_addressOut_valid(io_connPE_45_valid),
		.io_addressOut_bits(io_connPE_45_bits)
	);
	AllocatorBuffer queues_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_46_io_addressIn_ready),
		.io_addressIn_valid(_casServers_46_io_addressOut_valid),
		.io_addressIn_bits(_casServers_46_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_46_ready),
		.io_addressOut_valid(io_connPE_46_valid),
		.io_addressOut_bits(io_connPE_46_bits)
	);
	AllocatorBuffer queues_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_47_io_addressIn_ready),
		.io_addressIn_valid(_casServers_47_io_addressOut_valid),
		.io_addressIn_bits(_casServers_47_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_47_ready),
		.io_addressOut_valid(io_connPE_47_valid),
		.io_addressOut_bits(io_connPE_47_bits)
	);
	AllocatorBuffer queues_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_48_io_addressIn_ready),
		.io_addressIn_valid(_casServers_48_io_addressOut_valid),
		.io_addressIn_bits(_casServers_48_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_48_ready),
		.io_addressOut_valid(io_connPE_48_valid),
		.io_addressOut_bits(io_connPE_48_bits)
	);
	AllocatorBuffer queues_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_49_io_addressIn_ready),
		.io_addressIn_valid(_casServers_49_io_addressOut_valid),
		.io_addressIn_bits(_casServers_49_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_49_ready),
		.io_addressOut_valid(io_connPE_49_valid),
		.io_addressOut_bits(io_connPE_49_bits)
	);
	AllocatorBuffer queues_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_50_io_addressIn_ready),
		.io_addressIn_valid(_casServers_50_io_addressOut_valid),
		.io_addressIn_bits(_casServers_50_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_50_ready),
		.io_addressOut_valid(io_connPE_50_valid),
		.io_addressOut_bits(io_connPE_50_bits)
	);
	AllocatorBuffer queues_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_51_io_addressIn_ready),
		.io_addressIn_valid(_casServers_51_io_addressOut_valid),
		.io_addressIn_bits(_casServers_51_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_51_ready),
		.io_addressOut_valid(io_connPE_51_valid),
		.io_addressOut_bits(io_connPE_51_bits)
	);
	AllocatorBuffer queues_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_52_io_addressIn_ready),
		.io_addressIn_valid(_casServers_52_io_addressOut_valid),
		.io_addressIn_bits(_casServers_52_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_52_ready),
		.io_addressOut_valid(io_connPE_52_valid),
		.io_addressOut_bits(io_connPE_52_bits)
	);
	AllocatorBuffer queues_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_53_io_addressIn_ready),
		.io_addressIn_valid(_casServers_53_io_addressOut_valid),
		.io_addressIn_bits(_casServers_53_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_53_ready),
		.io_addressOut_valid(io_connPE_53_valid),
		.io_addressOut_bits(io_connPE_53_bits)
	);
	AllocatorBuffer queues_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_54_io_addressIn_ready),
		.io_addressIn_valid(_casServers_54_io_addressOut_valid),
		.io_addressIn_bits(_casServers_54_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_54_ready),
		.io_addressOut_valid(io_connPE_54_valid),
		.io_addressOut_bits(io_connPE_54_bits)
	);
	AllocatorBuffer queues_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_55_io_addressIn_ready),
		.io_addressIn_valid(_casServers_55_io_addressOut_valid),
		.io_addressIn_bits(_casServers_55_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_55_ready),
		.io_addressOut_valid(io_connPE_55_valid),
		.io_addressOut_bits(io_connPE_55_bits)
	);
	AllocatorBuffer queues_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_56_io_addressIn_ready),
		.io_addressIn_valid(_casServers_56_io_addressOut_valid),
		.io_addressIn_bits(_casServers_56_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_56_ready),
		.io_addressOut_valid(io_connPE_56_valid),
		.io_addressOut_bits(io_connPE_56_bits)
	);
	AllocatorBuffer queues_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_57_io_addressIn_ready),
		.io_addressIn_valid(_casServers_57_io_addressOut_valid),
		.io_addressIn_bits(_casServers_57_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_57_ready),
		.io_addressOut_valid(io_connPE_57_valid),
		.io_addressOut_bits(io_connPE_57_bits)
	);
	AllocatorBuffer queues_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_58_io_addressIn_ready),
		.io_addressIn_valid(_casServers_58_io_addressOut_valid),
		.io_addressIn_bits(_casServers_58_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_58_ready),
		.io_addressOut_valid(io_connPE_58_valid),
		.io_addressOut_bits(io_connPE_58_bits)
	);
	AllocatorBuffer queues_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_59_io_addressIn_ready),
		.io_addressIn_valid(_casServers_59_io_addressOut_valid),
		.io_addressIn_bits(_casServers_59_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_59_ready),
		.io_addressOut_valid(io_connPE_59_valid),
		.io_addressOut_bits(io_connPE_59_bits)
	);
	AllocatorBuffer queues_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_60_io_addressIn_ready),
		.io_addressIn_valid(_casServers_60_io_addressOut_valid),
		.io_addressIn_bits(_casServers_60_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_60_ready),
		.io_addressOut_valid(io_connPE_60_valid),
		.io_addressOut_bits(io_connPE_60_bits)
	);
	AllocatorBuffer queues_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_61_io_addressIn_ready),
		.io_addressIn_valid(_casServers_61_io_addressOut_valid),
		.io_addressIn_bits(_casServers_61_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_61_ready),
		.io_addressOut_valid(io_connPE_61_valid),
		.io_addressOut_bits(io_connPE_61_bits)
	);
	AllocatorBuffer queues_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_62_io_addressIn_ready),
		.io_addressIn_valid(_casServers_62_io_addressOut_valid),
		.io_addressIn_bits(_casServers_62_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_62_ready),
		.io_addressOut_valid(io_connPE_62_valid),
		.io_addressOut_bits(io_connPE_62_bits)
	);
	AllocatorBuffer queues_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_63_io_addressIn_ready),
		.io_addressIn_valid(_casServers_63_io_addressOut_valid),
		.io_addressIn_bits(_casServers_63_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_63_ready),
		.io_addressOut_valid(io_connPE_63_valid),
		.io_addressOut_bits(io_connPE_63_bits)
	);
endmodule
module AllocatorServer (
	clock,
	reset,
	io_dataOut_ready,
	io_dataOut_valid,
	io_dataOut_bits,
	io_axi_mgmt_ar_ready,
	io_axi_mgmt_ar_valid,
	io_axi_mgmt_ar_bits_addr,
	io_axi_mgmt_ar_bits_prot,
	io_axi_mgmt_r_ready,
	io_axi_mgmt_r_valid,
	io_axi_mgmt_r_bits_data,
	io_axi_mgmt_r_bits_resp,
	io_axi_mgmt_aw_ready,
	io_axi_mgmt_aw_valid,
	io_axi_mgmt_aw_bits_addr,
	io_axi_mgmt_aw_bits_prot,
	io_axi_mgmt_w_ready,
	io_axi_mgmt_w_valid,
	io_axi_mgmt_w_bits_data,
	io_axi_mgmt_w_bits_strb,
	io_axi_mgmt_b_ready,
	io_axi_mgmt_b_valid,
	io_axi_mgmt_b_bits_resp,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits
);
	input clock;
	input reset;
	input io_dataOut_ready;
	output wire io_dataOut_valid;
	output wire [63:0] io_dataOut_bits;
	output wire io_axi_mgmt_ar_ready;
	input io_axi_mgmt_ar_valid;
	input [5:0] io_axi_mgmt_ar_bits_addr;
	input [2:0] io_axi_mgmt_ar_bits_prot;
	input io_axi_mgmt_r_ready;
	output wire io_axi_mgmt_r_valid;
	output wire [63:0] io_axi_mgmt_r_bits_data;
	output wire [1:0] io_axi_mgmt_r_bits_resp;
	output wire io_axi_mgmt_aw_ready;
	input io_axi_mgmt_aw_valid;
	input [5:0] io_axi_mgmt_aw_bits_addr;
	input [2:0] io_axi_mgmt_aw_bits_prot;
	output wire io_axi_mgmt_w_ready;
	input io_axi_mgmt_w_valid;
	input [63:0] io_axi_mgmt_w_bits_data;
	input [7:0] io_axi_mgmt_w_bits_strb;
	input io_axi_mgmt_b_ready;
	output wire io_axi_mgmt_b_valid;
	output wire [1:0] io_axi_mgmt_b_bits_resp;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [63:0] io_read_data_bits;
	wire _wrRespQueue__io_enq_ready;
	wire _wrRespQueue__io_deq_valid;
	wire _wrReqData__deq_q_io_enq_ready;
	wire _wrReqData__deq_q_io_deq_valid;
	wire [63:0] _wrReqData__deq_q_io_deq_bits_data;
	wire [7:0] _wrReqData__deq_q_io_deq_bits_strb;
	wire _wrReq__deq_q_io_enq_ready;
	wire _wrReq__deq_q_io_deq_valid;
	wire [5:0] _wrReq__deq_q_io_deq_bits_addr;
	wire _rdRespQueue__io_enq_ready;
	wire _rdRespQueue__io_deq_valid;
	wire [63:0] _rdRespQueue__io_deq_bits_data;
	wire [1:0] _rdRespQueue__io_deq_bits_resp;
	wire _rdReq__deq_q_io_enq_ready;
	wire _rdReq__deq_q_io_deq_valid;
	wire [5:0] _rdReq__deq_q_io_deq_bits_addr;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	wire rdReq = _rdReq__deq_q_io_deq_valid & _rdRespQueue__io_enq_ready;
	wire wrReq = (_wrReq__deq_q_io_deq_valid & _wrReqData__deq_q_io_deq_valid) & _wrRespQueue__io_enq_ready;
	reg [63:0] rAddr;
	reg [63:0] rPause;
	reg [63:0] avaialbleSize;
	reg [2:0] stateReg;
	reg [63:0] continuationsRegisters_0;
	reg [63:0] continuationsRegisters_1;
	reg [63:0] continuationsRegisters_2;
	reg [63:0] continuationsRegisters_3;
	reg [63:0] continuationsRegisters_4;
	reg [63:0] continuationsRegisters_5;
	reg [63:0] continuationsRegisters_6;
	reg [63:0] continuationsRegisters_7;
	reg [63:0] continuationsRegisters_8;
	reg [63:0] continuationsRegisters_9;
	reg [63:0] continuationsRegisters_10;
	reg [63:0] continuationsRegisters_11;
	reg [63:0] continuationsRegisters_12;
	reg [63:0] continuationsRegisters_13;
	reg [63:0] continuationsRegisters_14;
	reg [63:0] continuationsRegisters_15;
	reg [3:0] burstCounter;
	wire io_read_address_valid_0 = stateReg == 3'h1;
	wire _GEN = stateReg == 3'h2;
	wire _GEN_0 = stateReg == 3'h3;
	wire [1023:0] _GEN_1 = {continuationsRegisters_15, continuationsRegisters_14, continuationsRegisters_13, continuationsRegisters_12, continuationsRegisters_11, continuationsRegisters_10, continuationsRegisters_9, continuationsRegisters_8, continuationsRegisters_7, continuationsRegisters_6, continuationsRegisters_5, continuationsRegisters_4, continuationsRegisters_3, continuationsRegisters_2, continuationsRegisters_1, continuationsRegisters_0};
	always @(posedge clock)
		if (reset) begin
			rAddr <= 64'h0000000000000000;
			rPause <= 64'h0000000000000000;
			avaialbleSize <= 64'h0000000000000000;
			stateReg <= 3'h0;
			continuationsRegisters_0 <= 64'h0000000000000000;
			continuationsRegisters_1 <= 64'h0000000000000000;
			continuationsRegisters_2 <= 64'h0000000000000000;
			continuationsRegisters_3 <= 64'h0000000000000000;
			continuationsRegisters_4 <= 64'h0000000000000000;
			continuationsRegisters_5 <= 64'h0000000000000000;
			continuationsRegisters_6 <= 64'h0000000000000000;
			continuationsRegisters_7 <= 64'h0000000000000000;
			continuationsRegisters_8 <= 64'h0000000000000000;
			continuationsRegisters_9 <= 64'h0000000000000000;
			continuationsRegisters_10 <= 64'h0000000000000000;
			continuationsRegisters_11 <= 64'h0000000000000000;
			continuationsRegisters_12 <= 64'h0000000000000000;
			continuationsRegisters_13 <= 64'h0000000000000000;
			continuationsRegisters_14 <= 64'h0000000000000000;
			continuationsRegisters_15 <= 64'h0000000000000000;
			burstCounter <= 4'hf;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_2;
			reg _GEN_3;
			reg _GEN_4;
			reg _GEN_5;
			_GEN_2 = stateReg == 3'h0;
			_GEN_3 = burstCounter == 4'h0;
			_GEN_4 = _GEN_2 | io_read_address_valid_0;
			_GEN_5 = _GEN_3 & io_read_data_valid;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h1))
				rAddr <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rAddr[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rAddr[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rAddr[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rAddr[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rAddr[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rAddr[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rAddr[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rAddr[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h0))
				rPause <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rPause[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rPause[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rPause[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rPause[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rPause[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rPause[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rPause[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rPause[7:0])};
			else if (~_GEN_2 | (|avaialbleSize[63:4]))
				;
			else
				rPause <= 64'hffffffffffffffff;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h2))
				avaialbleSize <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : avaialbleSize[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : avaialbleSize[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : avaialbleSize[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : avaialbleSize[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : avaialbleSize[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : avaialbleSize[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : avaialbleSize[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : avaialbleSize[7:0])};
			else if (_GEN_4 | ~_GEN)
				;
			else if (_GEN_5)
				avaialbleSize <= avaialbleSize - 64'h0000000000000001;
			else if (io_read_data_valid)
				avaialbleSize <= avaialbleSize - 64'h0000000000000001;
			if (_GEN_2)
				stateReg <= (|avaialbleSize[63:4] ? 3'h1 : 3'h4);
			else if (io_read_address_valid_0) begin
				if (io_read_address_ready) begin
					stateReg <= 3'h2;
					burstCounter <= 4'hf;
				end
			end
			else if (_GEN) begin
				if (_GEN_5) begin
					stateReg <= 3'h3;
					burstCounter <= 4'hf;
				end
				else if (io_read_data_valid)
					burstCounter <= burstCounter - 4'h1;
			end
			else begin
				if ((_GEN_0 ? _GEN_3 & io_dataOut_ready : (stateReg == 3'h4) & (rPause == 64'h0000000000000000)))
					stateReg <= 3'h0;
				if (_GEN_0 & io_dataOut_ready)
					burstCounter <= burstCounter - 4'h1;
			end
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & _GEN_3))
				;
			else
				continuationsRegisters_0 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h1)))
				;
			else
				continuationsRegisters_1 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h2)))
				;
			else
				continuationsRegisters_2 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h3)))
				;
			else
				continuationsRegisters_3 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h4)))
				;
			else
				continuationsRegisters_4 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h5)))
				;
			else
				continuationsRegisters_5 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h6)))
				;
			else
				continuationsRegisters_6 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h7)))
				;
			else
				continuationsRegisters_7 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h8)))
				;
			else
				continuationsRegisters_8 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h9)))
				;
			else
				continuationsRegisters_9 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'ha)))
				;
			else
				continuationsRegisters_10 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'hb)))
				;
			else
				continuationsRegisters_11 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'hc)))
				;
			else
				continuationsRegisters_12 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'hd)))
				;
			else
				continuationsRegisters_13 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'he)))
				;
			else
				continuationsRegisters_14 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (&burstCounter)))
				;
			else
				continuationsRegisters_15 <= io_read_data_bits;
		end
	Queue2_AddressChannel_2 s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_ar_ready),
		.io_enq_valid(io_axi_mgmt_ar_valid),
		.io_enq_bits_addr(io_axi_mgmt_ar_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_ar_bits_prot),
		.io_deq_ready(_rdReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_rdRespQueue__io_deq_valid),
		.io_enq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_enq_bits_resp(_rdRespQueue__io_deq_bits_resp),
		.io_deq_ready(io_axi_mgmt_r_ready),
		.io_deq_valid(io_axi_mgmt_r_valid),
		.io_deq_bits_data(io_axi_mgmt_r_bits_data),
		.io_deq_bits_resp(io_axi_mgmt_r_bits_resp)
	);
	Queue2_AddressChannel_2 s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_aw_ready),
		.io_enq_valid(io_axi_mgmt_aw_valid),
		.io_enq_bits_addr(io_axi_mgmt_aw_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_aw_bits_prot),
		.io_deq_ready(_wrReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_w_ready),
		.io_enq_valid(io_axi_mgmt_w_valid),
		.io_enq_bits_data(io_axi_mgmt_w_bits_data),
		.io_enq_bits_strb(io_axi_mgmt_w_bits_strb),
		.io_deq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_wrRespQueue__io_deq_valid),
		.io_enq_bits_resp(2'h0),
		.io_deq_ready(io_axi_mgmt_b_ready),
		.io_deq_valid(io_axi_mgmt_b_valid),
		.io_deq_bits_resp(io_axi_mgmt_b_bits_resp)
	);
	Queue1_AddressChannel rdReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_deq_ready(rdReq),
		.io_deq_valid(_rdReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_rdReq__deq_q_io_deq_bits_addr)
	);
	Queue1_ReadDataChannel rdRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdRespQueue__io_enq_ready),
		.io_enq_valid(rdReq),
		.io_enq_bits_data((_rdReq__deq_q_io_deq_bits_addr[5:3] == 3'h2 ? avaialbleSize : (_rdReq__deq_q_io_deq_bits_addr[5:3] == 3'h1 ? rAddr : (_rdReq__deq_q_io_deq_bits_addr[5:3] == 3'h0 ? rPause : 64'hffffffffffffffff)))),
		.io_deq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_deq_valid(_rdRespQueue__io_deq_valid),
		.io_deq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_deq_bits_resp(_rdRespQueue__io_deq_bits_resp)
	);
	Queue1_AddressChannel wrReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_wrReq__deq_q_io_deq_bits_addr)
	);
	Queue1_WriteDataChannel wrReqData__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_enq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_enq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReqData__deq_q_io_deq_valid),
		.io_deq_bits_data(_wrReqData__deq_q_io_deq_bits_data),
		.io_deq_bits_strb(_wrReqData__deq_q_io_deq_bits_strb)
	);
	Queue1_WriteResponseChannel wrRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrRespQueue__io_enq_ready),
		.io_enq_valid(wrReq),
		.io_deq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_deq_valid(_wrRespQueue__io_deq_valid)
	);
	assign io_dataOut_valid = ~(io_read_address_valid_0 | _GEN) & _GEN_0;
	assign io_dataOut_bits = _GEN_1[burstCounter * 64+:64];
	assign io_read_address_valid = io_read_address_valid_0;
	assign io_read_address_bits = rAddr + {avaialbleSize[60:0] - 61'h0000000000000010, 3'h0};
	assign io_read_data_ready = ~io_read_address_valid_0 & _GEN;
endmodule
module RVtoAXIBridge_4 (
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data
);
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [63:0] io_read_data_bits;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire axi_r_ready;
	input axi_r_valid;
	input [63:0] axi_r_bits_data;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_r_ready = io_read_data_ready;
endmodule
module ram_2x94 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [93:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [93:0] W0_data;
	reg [93:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 94'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadAddressChannel_6 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [93:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x94 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({29'h00000b0f, io_enq_bits_addr, 1'h0})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[0];
	assign io_deq_bits_addr = _ram_ext_R0_data[64:1];
	assign io_deq_bits_len = _ram_ext_R0_data[72:65];
	assign io_deq_bits_size = _ram_ext_R0_data[75:73];
	assign io_deq_bits_burst = _ram_ext_R0_data[77:76];
	assign io_deq_bits_lock = _ram_ext_R0_data[78];
	assign io_deq_bits_cache = _ram_ext_R0_data[82:79];
	assign io_deq_bits_prot = _ram_ext_R0_data[85:83];
	assign io_deq_bits_qos = _ram_ext_R0_data[89:86];
	assign io_deq_bits_region = _ram_ext_R0_data[93:90];
endmodule
module ram_2x64 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [63:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [63:0] W0_data;
	reg [63:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel_11 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits_id;
	input [63:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x64 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_data)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module Queue2_WriteAddressChannel_6 (
	clock,
	reset,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	reg wrap_1;
	always @(posedge clock)
		if (reset)
			wrap_1 <= 1'h0;
		else if (io_deq_ready & wrap_1)
			wrap_1 <= wrap_1 - 1'h1;
	assign io_deq_valid = wrap_1;
	assign io_deq_bits_id = 1'h0;
	assign io_deq_bits_addr = 64'h0000000000000000;
	assign io_deq_bits_len = 8'h00;
	assign io_deq_bits_size = 3'h0;
	assign io_deq_bits_burst = 2'h0;
	assign io_deq_bits_lock = 1'h0;
	assign io_deq_bits_cache = 4'h0;
	assign io_deq_bits_prot = 3'h0;
	assign io_deq_bits_qos = 4'h0;
	assign io_deq_bits_region = 4'h0;
endmodule
module ram_2x73 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [72:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [72:0] W0_data;
	reg [72:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 73'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteDataChannel_11 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [7:0] io_enq_bits_strb;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [7:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	wire [72:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x73 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_strb, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[63:0];
	assign io_deq_bits_strb = _ram_ext_R0_data[71:64];
	assign io_deq_bits_last = _ram_ext_R0_data[72];
endmodule
module Queue2_WriteResponseChannel_11 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	reg wrap;
	reg maybe_full;
	wire full = ~wrap & maybe_full;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_enq;
			do_enq = ~full & io_enq_valid;
			if (do_enq) begin
				wrap <= wrap - 1'h1;
				maybe_full <= do_enq;
			end
		end
	assign io_enq_ready = ~full;
endmodule
module ram_2x96 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [95:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [95:0] W0_data;
	reg [95:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 96'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadAddressChannel_10 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_id;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [95:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x96 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[2:0];
	assign io_deq_bits_addr = _ram_ext_R0_data[66:3];
	assign io_deq_bits_len = _ram_ext_R0_data[74:67];
	assign io_deq_bits_size = _ram_ext_R0_data[77:75];
	assign io_deq_bits_burst = _ram_ext_R0_data[79:78];
	assign io_deq_bits_lock = _ram_ext_R0_data[80];
	assign io_deq_bits_cache = _ram_ext_R0_data[84:81];
	assign io_deq_bits_prot = _ram_ext_R0_data[87:85];
	assign io_deq_bits_qos = _ram_ext_R0_data[91:88];
	assign io_deq_bits_region = _ram_ext_R0_data[95:92];
endmodule
module ram_2x70 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [69:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [69:0] W0_data;
	reg [69:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 70'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel_15 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_data,
	io_deq_bits_resp,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_id;
	input [63:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	output wire io_deq_bits_last;
	wire [69:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x70 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_resp, io_enq_bits_data, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[2:0];
	assign io_deq_bits_data = _ram_ext_R0_data[66:3];
	assign io_deq_bits_resp = _ram_ext_R0_data[68:67];
	assign io_deq_bits_last = _ram_ext_R0_data[69];
endmodule
module Queue2_WriteAddressChannel_10 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_id;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [95:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x96 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[2:0];
	assign io_deq_bits_addr = _ram_ext_R0_data[66:3];
	assign io_deq_bits_len = _ram_ext_R0_data[74:67];
	assign io_deq_bits_size = _ram_ext_R0_data[77:75];
	assign io_deq_bits_burst = _ram_ext_R0_data[79:78];
	assign io_deq_bits_lock = _ram_ext_R0_data[80];
	assign io_deq_bits_cache = _ram_ext_R0_data[84:81];
	assign io_deq_bits_prot = _ram_ext_R0_data[87:85];
	assign io_deq_bits_qos = _ram_ext_R0_data[91:88];
	assign io_deq_bits_region = _ram_ext_R0_data[95:92];
endmodule
module ram_2x3 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [2:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [2:0] W0_data;
	reg [2:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 3'bxxx);
endmodule
module Queue2_WriteResponseChannel_15 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_id;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_id;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x3 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_id),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_id)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module elasticArbiter_4 (
	clock,
	reset,
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_id,
	io_sources_0_bits_addr,
	io_sources_0_bits_len,
	io_sources_0_bits_size,
	io_sources_0_bits_burst,
	io_sources_0_bits_lock,
	io_sources_0_bits_cache,
	io_sources_0_bits_prot,
	io_sources_0_bits_qos,
	io_sources_0_bits_region,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_id,
	io_sources_1_bits_addr,
	io_sources_1_bits_len,
	io_sources_1_bits_size,
	io_sources_1_bits_burst,
	io_sources_1_bits_lock,
	io_sources_1_bits_cache,
	io_sources_1_bits_prot,
	io_sources_1_bits_qos,
	io_sources_1_bits_region,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_id,
	io_sources_2_bits_addr,
	io_sources_2_bits_len,
	io_sources_2_bits_size,
	io_sources_2_bits_burst,
	io_sources_2_bits_lock,
	io_sources_2_bits_cache,
	io_sources_2_bits_prot,
	io_sources_2_bits_qos,
	io_sources_2_bits_region,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_id,
	io_sources_3_bits_addr,
	io_sources_3_bits_len,
	io_sources_3_bits_size,
	io_sources_3_bits_burst,
	io_sources_3_bits_lock,
	io_sources_3_bits_cache,
	io_sources_3_bits_prot,
	io_sources_3_bits_qos,
	io_sources_3_bits_region,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_id,
	io_sink_bits_addr,
	io_sink_bits_len,
	io_sink_bits_size,
	io_sink_bits_burst,
	io_sink_bits_lock,
	io_sink_bits_cache,
	io_sink_bits_prot,
	io_sink_bits_qos,
	io_sink_bits_region,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	input clock;
	input reset;
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [2:0] io_sources_0_bits_id;
	input [63:0] io_sources_0_bits_addr;
	input [7:0] io_sources_0_bits_len;
	input [2:0] io_sources_0_bits_size;
	input [1:0] io_sources_0_bits_burst;
	input io_sources_0_bits_lock;
	input [3:0] io_sources_0_bits_cache;
	input [2:0] io_sources_0_bits_prot;
	input [3:0] io_sources_0_bits_qos;
	input [3:0] io_sources_0_bits_region;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [2:0] io_sources_1_bits_id;
	input [63:0] io_sources_1_bits_addr;
	input [7:0] io_sources_1_bits_len;
	input [2:0] io_sources_1_bits_size;
	input [1:0] io_sources_1_bits_burst;
	input io_sources_1_bits_lock;
	input [3:0] io_sources_1_bits_cache;
	input [2:0] io_sources_1_bits_prot;
	input [3:0] io_sources_1_bits_qos;
	input [3:0] io_sources_1_bits_region;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [2:0] io_sources_2_bits_id;
	input [63:0] io_sources_2_bits_addr;
	input [7:0] io_sources_2_bits_len;
	input [2:0] io_sources_2_bits_size;
	input [1:0] io_sources_2_bits_burst;
	input io_sources_2_bits_lock;
	input [3:0] io_sources_2_bits_cache;
	input [2:0] io_sources_2_bits_prot;
	input [3:0] io_sources_2_bits_qos;
	input [3:0] io_sources_2_bits_region;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [2:0] io_sources_3_bits_id;
	input [63:0] io_sources_3_bits_addr;
	input [7:0] io_sources_3_bits_len;
	input [2:0] io_sources_3_bits_size;
	input [1:0] io_sources_3_bits_burst;
	input io_sources_3_bits_lock;
	input [3:0] io_sources_3_bits_cache;
	input [2:0] io_sources_3_bits_prot;
	input [3:0] io_sources_3_bits_qos;
	input [3:0] io_sources_3_bits_region;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [2:0] io_sink_bits_id;
	output wire [63:0] io_sink_bits_addr;
	output wire [7:0] io_sink_bits_len;
	output wire [2:0] io_sink_bits_size;
	output wire [1:0] io_sink_bits_burst;
	output wire io_sink_bits_lock;
	output wire [3:0] io_sink_bits_cache;
	output wire [2:0] io_sink_bits_prot;
	output wire [3:0] io_sink_bits_qos;
	output wire [3:0] io_sink_bits_region;
	input io_select_ready;
	output wire io_select_valid;
	output wire [1:0] io_select_bits;
	wire sourceReady;
	reg [1:0] chooser_lastChoice;
	wire _chooser_rrChoice_T_4 = (chooser_lastChoice == 2'h0) & io_sources_1_valid;
	wire [1:0] _chooser_rrChoice_T_9 = {1'h1, ~(~chooser_lastChoice[1] & io_sources_2_valid)};
	wire [1:0] chooser_rrChoice = (&chooser_lastChoice ? 2'h0 : (_chooser_rrChoice_T_4 ? 2'h1 : _chooser_rrChoice_T_9));
	wire [1:0] chooser_priorityChoice = (io_sources_0_valid ? 2'h0 : (io_sources_1_valid ? 2'h1 : {1'h1, ~io_sources_2_valid}));
	wire [3:0] _GEN = {io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [1:0] io_select_bits_0 = (_GEN[chooser_rrChoice] ? chooser_rrChoice : chooser_priorityChoice);
	wire [11:0] _GEN_0 = {io_sources_3_bits_id, io_sources_2_bits_id, io_sources_1_bits_id, io_sources_0_bits_id};
	wire [255:0] _GEN_1 = {io_sources_3_bits_addr, io_sources_2_bits_addr, io_sources_1_bits_addr, io_sources_0_bits_addr};
	wire [31:0] _GEN_2 = {io_sources_3_bits_len, io_sources_2_bits_len, io_sources_1_bits_len, io_sources_0_bits_len};
	wire [11:0] _GEN_3 = {io_sources_3_bits_size, io_sources_2_bits_size, io_sources_1_bits_size, io_sources_0_bits_size};
	wire [7:0] _GEN_4 = {io_sources_3_bits_burst, io_sources_2_bits_burst, io_sources_1_bits_burst, io_sources_0_bits_burst};
	wire [3:0] _GEN_5 = {io_sources_3_bits_lock, io_sources_2_bits_lock, io_sources_1_bits_lock, io_sources_0_bits_lock};
	wire [15:0] _GEN_6 = {io_sources_3_bits_cache, io_sources_2_bits_cache, io_sources_1_bits_cache, io_sources_0_bits_cache};
	wire [11:0] _GEN_7 = {io_sources_3_bits_prot, io_sources_2_bits_prot, io_sources_1_bits_prot, io_sources_0_bits_prot};
	wire [15:0] _GEN_8 = {io_sources_3_bits_qos, io_sources_2_bits_qos, io_sources_1_bits_qos, io_sources_0_bits_qos};
	wire [15:0] _GEN_9 = {io_sources_3_bits_region, io_sources_2_bits_region, io_sources_1_bits_region, io_sources_0_bits_region};
	reg sinkSent;
	reg selectSent;
	assign sourceReady = (sinkSent | io_sink_ready) & (selectSent | io_select_ready);
	always @(posedge clock)
		if (reset) begin
			chooser_lastChoice <= 2'h0;
			sinkSent <= 1'h0;
			selectSent <= 1'h0;
		end
		else begin
			if (_GEN[io_select_bits_0] & sourceReady) begin
				if (_GEN[chooser_rrChoice]) begin
					if (&chooser_lastChoice)
						chooser_lastChoice <= 2'h0;
					else if (_chooser_rrChoice_T_4)
						chooser_lastChoice <= 2'h1;
					else
						chooser_lastChoice <= _chooser_rrChoice_T_9;
				end
				else
					chooser_lastChoice <= chooser_priorityChoice;
			end
			sinkSent <= ((io_sink_ready | sinkSent) & _GEN[io_select_bits_0]) & ~sourceReady;
			selectSent <= ((io_select_ready | selectSent) & _GEN[io_select_bits_0]) & ~sourceReady;
		end
	assign io_sources_0_ready = sourceReady & (io_select_bits_0 == 2'h0);
	assign io_sources_1_ready = sourceReady & (io_select_bits_0 == 2'h1);
	assign io_sources_2_ready = sourceReady & (io_select_bits_0 == 2'h2);
	assign io_sources_3_ready = sourceReady & (&io_select_bits_0);
	assign io_sink_valid = _GEN[io_select_bits_0] & ~sinkSent;
	assign io_sink_bits_id = _GEN_0[io_select_bits_0 * 3+:3];
	assign io_sink_bits_addr = _GEN_1[io_select_bits_0 * 64+:64];
	assign io_sink_bits_len = _GEN_2[io_select_bits_0 * 8+:8];
	assign io_sink_bits_size = _GEN_3[io_select_bits_0 * 3+:3];
	assign io_sink_bits_burst = _GEN_4[io_select_bits_0 * 2+:2];
	assign io_sink_bits_lock = _GEN_5[io_select_bits_0];
	assign io_sink_bits_cache = _GEN_6[io_select_bits_0 * 4+:4];
	assign io_sink_bits_prot = _GEN_7[io_select_bits_0 * 3+:3];
	assign io_sink_bits_qos = _GEN_8[io_select_bits_0 * 4+:4];
	assign io_sink_bits_region = _GEN_9[io_select_bits_0 * 4+:4];
	assign io_select_valid = _GEN[io_select_bits_0] & ~selectSent;
	assign io_select_bits = io_select_bits_0;
endmodule
module elasticDemux_7 (
	io_source_ready,
	io_source_valid,
	io_source_bits_id,
	io_source_bits_data,
	io_source_bits_resp,
	io_source_bits_last,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_id,
	io_sinks_0_bits_data,
	io_sinks_0_bits_resp,
	io_sinks_0_bits_last,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_id,
	io_sinks_1_bits_data,
	io_sinks_1_bits_resp,
	io_sinks_1_bits_last,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_2_bits_id,
	io_sinks_2_bits_data,
	io_sinks_2_bits_resp,
	io_sinks_2_bits_last,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_3_bits_id,
	io_sinks_3_bits_data,
	io_sinks_3_bits_resp,
	io_sinks_3_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [2:0] io_source_bits_id;
	input [63:0] io_source_bits_data;
	input [1:0] io_source_bits_resp;
	input io_source_bits_last;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [2:0] io_sinks_0_bits_id;
	output wire [63:0] io_sinks_0_bits_data;
	output wire [1:0] io_sinks_0_bits_resp;
	output wire io_sinks_0_bits_last;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [2:0] io_sinks_1_bits_id;
	output wire [63:0] io_sinks_1_bits_data;
	output wire [1:0] io_sinks_1_bits_resp;
	output wire io_sinks_1_bits_last;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	output wire [2:0] io_sinks_2_bits_id;
	output wire [63:0] io_sinks_2_bits_data;
	output wire [1:0] io_sinks_2_bits_resp;
	output wire io_sinks_2_bits_last;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire [2:0] io_sinks_3_bits_id;
	output wire [63:0] io_sinks_3_bits_data;
	output wire [1:0] io_sinks_3_bits_resp;
	output wire io_sinks_3_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input [1:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [3:0] _GEN = {io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 2'h0);
	assign io_sinks_0_bits_id = io_source_bits_id;
	assign io_sinks_0_bits_data = io_source_bits_data;
	assign io_sinks_0_bits_resp = io_source_bits_resp;
	assign io_sinks_0_bits_last = io_source_bits_last;
	assign io_sinks_1_valid = valid & (io_select_bits == 2'h1);
	assign io_sinks_1_bits_id = io_source_bits_id;
	assign io_sinks_1_bits_data = io_source_bits_data;
	assign io_sinks_1_bits_resp = io_source_bits_resp;
	assign io_sinks_1_bits_last = io_source_bits_last;
	assign io_sinks_2_valid = valid & (io_select_bits == 2'h2);
	assign io_sinks_2_bits_id = io_source_bits_id;
	assign io_sinks_2_bits_data = io_source_bits_data;
	assign io_sinks_2_bits_resp = io_source_bits_resp;
	assign io_sinks_2_bits_last = io_source_bits_last;
	assign io_sinks_3_valid = valid & (&io_select_bits);
	assign io_sinks_3_bits_id = io_source_bits_id;
	assign io_sinks_3_bits_data = io_source_bits_data;
	assign io_sinks_3_bits_resp = io_source_bits_resp;
	assign io_sinks_3_bits_last = io_source_bits_last;
	assign io_select_ready = fire;
endmodule
module ram_32x2 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [4:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [1:0] R0_data;
	input [4:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [1:0] W0_data;
	reg [1:0] Memory [0:31];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 2'bxx);
endmodule
module Queue32_UInt2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits;
	wire io_enq_ready_0;
	wire [1:0] _ram_ext_R0_data;
	reg [4:0] enq_ptr_value;
	reg [4:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire io_deq_valid_0 = io_enq_valid | ~empty;
	wire do_deq = (~empty & io_deq_ready) & io_deq_valid_0;
	wire do_enq = (~(empty & io_deq_ready) & io_enq_ready_0) & io_enq_valid;
	assign io_enq_ready_0 = io_deq_ready | ~(ptr_match & maybe_full);
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 5'h00;
			deq_ptr_value <= 5'h00;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 5'h01;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 5'h01;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_32x2 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = io_enq_ready_0;
	assign io_deq_valid = io_deq_valid_0;
	assign io_deq_bits = (empty ? io_enq_bits : _ram_ext_R0_data);
endmodule
module elasticMux_4 (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_data,
	io_sources_0_bits_strb,
	io_sources_0_bits_last,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_data,
	io_sources_1_bits_strb,
	io_sources_1_bits_last,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_data,
	io_sources_2_bits_strb,
	io_sources_2_bits_last,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_data,
	io_sources_3_bits_strb,
	io_sources_3_bits_last,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_data,
	io_sink_bits_strb,
	io_sink_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [63:0] io_sources_0_bits_data;
	input [7:0] io_sources_0_bits_strb;
	input io_sources_0_bits_last;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [63:0] io_sources_1_bits_data;
	input [7:0] io_sources_1_bits_strb;
	input io_sources_1_bits_last;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [63:0] io_sources_2_bits_data;
	input [7:0] io_sources_2_bits_strb;
	input io_sources_2_bits_last;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [63:0] io_sources_3_bits_data;
	input [7:0] io_sources_3_bits_strb;
	input io_sources_3_bits_last;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [63:0] io_sink_bits_data;
	output wire [7:0] io_sink_bits_strb;
	output wire io_sink_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input [1:0] io_select_bits;
	wire [3:0] _GEN = {io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [255:0] _GEN_0 = {io_sources_3_bits_data, io_sources_2_bits_data, io_sources_1_bits_data, io_sources_0_bits_data};
	wire [31:0] _GEN_1 = {io_sources_3_bits_strb, io_sources_2_bits_strb, io_sources_1_bits_strb, io_sources_0_bits_strb};
	wire [3:0] _GEN_2 = {io_sources_3_bits_last, io_sources_2_bits_last, io_sources_1_bits_last, io_sources_0_bits_last};
	wire valid = io_select_valid & _GEN[io_select_bits];
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & (io_select_bits == 2'h0);
	assign io_sources_1_ready = fire & (io_select_bits == 2'h1);
	assign io_sources_2_ready = fire & (io_select_bits == 2'h2);
	assign io_sources_3_ready = fire & (&io_select_bits);
	assign io_sink_valid = valid;
	assign io_sink_bits_data = _GEN_0[io_select_bits * 64+:64];
	assign io_sink_bits_strb = _GEN_1[io_select_bits * 8+:8];
	assign io_sink_bits_last = _GEN_2[io_select_bits];
	assign io_select_ready = fire & _GEN_2[io_select_bits];
endmodule
module elasticDemux_8 (
	io_source_ready,
	io_source_valid,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire io_select_ready;
	input io_select_valid;
	input [1:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [3:0] _GEN = {io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 2'h0);
	assign io_sinks_1_valid = valid & (io_select_bits == 2'h1);
	assign io_sinks_2_valid = valid & (io_select_bits == 2'h2);
	assign io_sinks_3_valid = valid & (&io_select_bits);
	assign io_select_ready = fire;
endmodule
module axi4FullMux_2 (
	clock,
	reset,
	s_axi_0_ar_ready,
	s_axi_0_ar_valid,
	s_axi_0_ar_bits_addr,
	s_axi_0_r_ready,
	s_axi_0_r_valid,
	s_axi_0_r_bits_data,
	s_axi_1_ar_ready,
	s_axi_1_ar_valid,
	s_axi_1_ar_bits_addr,
	s_axi_1_r_ready,
	s_axi_1_r_valid,
	s_axi_1_r_bits_data,
	s_axi_2_ar_ready,
	s_axi_2_ar_valid,
	s_axi_2_ar_bits_addr,
	s_axi_2_r_ready,
	s_axi_2_r_valid,
	s_axi_2_r_bits_data,
	s_axi_3_ar_ready,
	s_axi_3_ar_valid,
	s_axi_3_ar_bits_addr,
	s_axi_3_r_ready,
	s_axi_3_r_valid,
	s_axi_3_r_bits_data,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_id,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_id,
	m_axi_r_bits_data,
	m_axi_r_bits_resp,
	m_axi_r_bits_last,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_id,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_strb,
	m_axi_w_bits_last,
	m_axi_b_ready,
	m_axi_b_valid,
	m_axi_b_bits_id,
	m_axi_b_bits_resp
);
	input clock;
	input reset;
	output wire s_axi_0_ar_ready;
	input s_axi_0_ar_valid;
	input [63:0] s_axi_0_ar_bits_addr;
	input s_axi_0_r_ready;
	output wire s_axi_0_r_valid;
	output wire [63:0] s_axi_0_r_bits_data;
	output wire s_axi_1_ar_ready;
	input s_axi_1_ar_valid;
	input [63:0] s_axi_1_ar_bits_addr;
	input s_axi_1_r_ready;
	output wire s_axi_1_r_valid;
	output wire [63:0] s_axi_1_r_bits_data;
	output wire s_axi_2_ar_ready;
	input s_axi_2_ar_valid;
	input [63:0] s_axi_2_ar_bits_addr;
	input s_axi_2_r_ready;
	output wire s_axi_2_r_valid;
	output wire [63:0] s_axi_2_r_bits_data;
	output wire s_axi_3_ar_ready;
	input s_axi_3_ar_valid;
	input [63:0] s_axi_3_ar_bits_addr;
	input s_axi_3_r_ready;
	output wire s_axi_3_r_valid;
	output wire [63:0] s_axi_3_r_bits_data;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [2:0] m_axi_ar_bits_id;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [2:0] m_axi_r_bits_id;
	input [63:0] m_axi_r_bits_data;
	input [1:0] m_axi_r_bits_resp;
	input m_axi_r_bits_last;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [2:0] m_axi_aw_bits_id;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [63:0] m_axi_w_bits_data;
	output wire [7:0] m_axi_w_bits_strb;
	output wire m_axi_w_bits_last;
	output wire m_axi_b_ready;
	input m_axi_b_valid;
	input [2:0] m_axi_b_bits_id;
	input [1:0] m_axi_b_bits_resp;
	wire _write_demux_io_source_ready;
	wire _write_demux_io_sinks_0_valid;
	wire _write_demux_io_sinks_1_valid;
	wire _write_demux_io_sinks_2_valid;
	wire _write_demux_io_sinks_3_valid;
	wire _write_demux_io_select_ready;
	wire _write_mux_io_sources_0_ready;
	wire _write_mux_io_sources_1_ready;
	wire _write_mux_io_sources_2_ready;
	wire _write_mux_io_sources_3_ready;
	wire _write_mux_io_sink_valid;
	wire [63:0] _write_mux_io_sink_bits_data;
	wire [7:0] _write_mux_io_sink_bits_strb;
	wire _write_mux_io_sink_bits_last;
	wire _write_mux_io_select_ready;
	wire _write_arbiter_io_sources_0_ready;
	wire _write_arbiter_io_sources_1_ready;
	wire _write_arbiter_io_sources_2_ready;
	wire _write_arbiter_io_sources_3_ready;
	wire _write_arbiter_io_sink_valid;
	wire [2:0] _write_arbiter_io_sink_bits_id;
	wire [63:0] _write_arbiter_io_sink_bits_addr;
	wire [7:0] _write_arbiter_io_sink_bits_len;
	wire [2:0] _write_arbiter_io_sink_bits_size;
	wire [1:0] _write_arbiter_io_sink_bits_burst;
	wire _write_arbiter_io_sink_bits_lock;
	wire [3:0] _write_arbiter_io_sink_bits_cache;
	wire [2:0] _write_arbiter_io_sink_bits_prot;
	wire [3:0] _write_arbiter_io_sink_bits_qos;
	wire [3:0] _write_arbiter_io_sink_bits_region;
	wire _write_arbiter_io_select_valid;
	wire [1:0] _write_arbiter_io_select_bits;
	wire _write_portQueue_io_enq_ready;
	wire _write_portQueue_io_deq_valid;
	wire [1:0] _write_portQueue_io_deq_bits;
	wire _read_demux_io_source_ready;
	wire _read_demux_io_sinks_0_valid;
	wire [2:0] _read_demux_io_sinks_0_bits_id;
	wire [63:0] _read_demux_io_sinks_0_bits_data;
	wire [1:0] _read_demux_io_sinks_0_bits_resp;
	wire _read_demux_io_sinks_0_bits_last;
	wire _read_demux_io_sinks_1_valid;
	wire [2:0] _read_demux_io_sinks_1_bits_id;
	wire [63:0] _read_demux_io_sinks_1_bits_data;
	wire [1:0] _read_demux_io_sinks_1_bits_resp;
	wire _read_demux_io_sinks_1_bits_last;
	wire _read_demux_io_sinks_2_valid;
	wire [2:0] _read_demux_io_sinks_2_bits_id;
	wire [63:0] _read_demux_io_sinks_2_bits_data;
	wire [1:0] _read_demux_io_sinks_2_bits_resp;
	wire _read_demux_io_sinks_2_bits_last;
	wire _read_demux_io_sinks_3_valid;
	wire [2:0] _read_demux_io_sinks_3_bits_id;
	wire [63:0] _read_demux_io_sinks_3_bits_data;
	wire [1:0] _read_demux_io_sinks_3_bits_resp;
	wire _read_demux_io_sinks_3_bits_last;
	wire _read_demux_io_select_ready;
	wire _read_arbiter_io_sources_0_ready;
	wire _read_arbiter_io_sources_1_ready;
	wire _read_arbiter_io_sources_2_ready;
	wire _read_arbiter_io_sources_3_ready;
	wire _read_arbiter_io_sink_valid;
	wire [2:0] _read_arbiter_io_sink_bits_id;
	wire [63:0] _read_arbiter_io_sink_bits_addr;
	wire [7:0] _read_arbiter_io_sink_bits_len;
	wire [2:0] _read_arbiter_io_sink_bits_size;
	wire [1:0] _read_arbiter_io_sink_bits_burst;
	wire _read_arbiter_io_sink_bits_lock;
	wire [3:0] _read_arbiter_io_sink_bits_cache;
	wire [2:0] _read_arbiter_io_sink_bits_prot;
	wire [3:0] _read_arbiter_io_sink_bits_qos;
	wire [3:0] _read_arbiter_io_sink_bits_region;
	wire _m_axi__sinkBuffer_1_io_deq_valid;
	wire [2:0] _m_axi__sinkBuffer_1_io_deq_bits_id;
	wire _m_axi__sourceBuffer_2_io_enq_ready;
	wire _m_axi__sourceBuffer_1_io_enq_ready;
	wire _m_axi__sinkBuffer_io_deq_valid;
	wire [2:0] _m_axi__sinkBuffer_io_deq_bits_id;
	wire [63:0] _m_axi__sinkBuffer_io_deq_bits_data;
	wire [1:0] _m_axi__sinkBuffer_io_deq_bits_resp;
	wire _m_axi__sinkBuffer_io_deq_bits_last;
	wire _m_axi__sourceBuffer_io_enq_ready;
	wire _s_axi__buffered_sinkBuffer_7_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_11_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_11_io_deq_bits_data;
	wire [7:0] _s_axi__buffered_sourceBuffer_11_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_11_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_10_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_10_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_10_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_6_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_9_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_9_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_9_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_5_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_8_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_8_io_deq_bits_data;
	wire [7:0] _s_axi__buffered_sourceBuffer_8_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_8_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_7_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_7_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_7_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_4_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_6_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_6_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_6_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_3_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_data;
	wire [7:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_2_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_1_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_io_deq_valid;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_id;
	wire [63:0] _s_axi__buffered_sourceBuffer_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_region;
	reg read_eagerFork_regs_0;
	reg read_eagerFork_regs_1;
	wire read_eagerFork_m_axi__r_ready_qual1_0 = _read_demux_io_source_ready | read_eagerFork_regs_0;
	wire read_eagerFork_m_axi__r_ready_qual1_1 = _read_demux_io_select_ready | read_eagerFork_regs_1;
	wire m_axi__r_ready = read_eagerFork_m_axi__r_ready_qual1_0 & read_eagerFork_m_axi__r_ready_qual1_1;
	reg write_eagerFork_regs_0;
	reg write_eagerFork_regs_1;
	wire write_eagerFork_m_axi__b_ready_qual1_0 = _write_demux_io_source_ready | write_eagerFork_regs_0;
	wire write_eagerFork_m_axi__b_ready_qual1_1 = _write_demux_io_select_ready | write_eagerFork_regs_1;
	wire m_axi__b_ready = write_eagerFork_m_axi__b_ready_qual1_0 & write_eagerFork_m_axi__b_ready_qual1_1;
	always @(posedge clock)
		if (reset) begin
			read_eagerFork_regs_0 <= 1'h0;
			read_eagerFork_regs_1 <= 1'h0;
			write_eagerFork_regs_0 <= 1'h0;
			write_eagerFork_regs_1 <= 1'h0;
		end
		else begin
			read_eagerFork_regs_0 <= (read_eagerFork_m_axi__r_ready_qual1_0 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			read_eagerFork_regs_1 <= (read_eagerFork_m_axi__r_ready_qual1_1 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			write_eagerFork_regs_0 <= (write_eagerFork_m_axi__b_ready_qual1_0 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
			write_eagerFork_regs_1 <= (write_eagerFork_m_axi__b_ready_qual1_1 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
		end
	Queue2_ReadAddressChannel_6 s_axi__buffered_sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_ar_ready),
		.io_enq_valid(s_axi_0_ar_valid),
		.io_enq_bits_addr(s_axi_0_ar_bits_addr),
		.io_deq_ready(_read_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_11 s_axi__buffered_sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_0_valid),
		.io_enq_bits_id(_read_demux_io_sinks_0_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_deq_ready(s_axi_0_r_ready),
		.io_deq_valid(s_axi_0_r_valid),
		.io_deq_bits_data(s_axi_0_r_bits_data)
	);
	Queue2_WriteAddressChannel_6 s_axi__buffered_sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_deq_ready(_write_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_1_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_11 s_axi__buffered_sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(64'h0000000000000000),
		.io_enq_bits_strb(8'h00),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_11 s_axi__buffered_sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_0_valid)
	);
	Queue2_ReadAddressChannel_6 s_axi__buffered_sourceBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_ar_ready),
		.io_enq_valid(s_axi_1_ar_valid),
		.io_enq_bits_addr(s_axi_1_ar_bits_addr),
		.io_deq_ready(_read_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_3_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_11 s_axi__buffered_sinkBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_1_valid),
		.io_enq_bits_id(_read_demux_io_sinks_1_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_deq_ready(s_axi_1_r_ready),
		.io_deq_valid(s_axi_1_r_valid),
		.io_deq_bits_data(s_axi_1_r_bits_data)
	);
	Queue2_WriteAddressChannel_6 s_axi__buffered_sourceBuffer_4(
		.clock(clock),
		.reset(reset),
		.io_deq_ready(_write_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_4_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_11 s_axi__buffered_sourceBuffer_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(64'h0000000000000000),
		.io_enq_bits_strb(8'h00),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_11 s_axi__buffered_sinkBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_1_valid)
	);
	Queue2_ReadAddressChannel_6 s_axi__buffered_sourceBuffer_6(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_2_ar_ready),
		.io_enq_valid(s_axi_2_ar_valid),
		.io_enq_bits_addr(s_axi_2_ar_bits_addr),
		.io_deq_ready(_read_arbiter_io_sources_2_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_6_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_6_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_6_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_6_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_6_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_6_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_6_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_6_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_6_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_6_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_6_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_11 s_axi__buffered_sinkBuffer_4(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_4_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_2_valid),
		.io_enq_bits_id(_read_demux_io_sinks_2_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_2_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_2_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_2_bits_last),
		.io_deq_ready(s_axi_2_r_ready),
		.io_deq_valid(s_axi_2_r_valid),
		.io_deq_bits_data(s_axi_2_r_bits_data)
	);
	Queue2_WriteAddressChannel_6 s_axi__buffered_sourceBuffer_7(
		.clock(clock),
		.reset(reset),
		.io_deq_ready(_write_arbiter_io_sources_2_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_7_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_7_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_7_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_7_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_7_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_7_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_7_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_7_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_7_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_7_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_7_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_11 s_axi__buffered_sourceBuffer_8(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(64'h0000000000000000),
		.io_enq_bits_strb(8'h00),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_2_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_8_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_8_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_8_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_8_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_11 s_axi__buffered_sinkBuffer_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_5_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_2_valid)
	);
	Queue2_ReadAddressChannel_6 s_axi__buffered_sourceBuffer_9(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_3_ar_ready),
		.io_enq_valid(s_axi_3_ar_valid),
		.io_enq_bits_addr(s_axi_3_ar_bits_addr),
		.io_deq_ready(_read_arbiter_io_sources_3_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_9_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_9_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_9_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_9_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_9_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_9_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_9_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_9_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_9_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_9_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_9_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_11 s_axi__buffered_sinkBuffer_6(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_6_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_3_valid),
		.io_enq_bits_id(_read_demux_io_sinks_3_bits_id[0]),
		.io_enq_bits_data(_read_demux_io_sinks_3_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_3_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_3_bits_last),
		.io_deq_ready(s_axi_3_r_ready),
		.io_deq_valid(s_axi_3_r_valid),
		.io_deq_bits_data(s_axi_3_r_bits_data)
	);
	Queue2_WriteAddressChannel_6 s_axi__buffered_sourceBuffer_10(
		.clock(clock),
		.reset(reset),
		.io_deq_ready(_write_arbiter_io_sources_3_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_10_io_deq_valid),
		.io_deq_bits_id(_s_axi__buffered_sourceBuffer_10_io_deq_bits_id),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_10_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_10_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_10_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_10_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_10_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_10_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_10_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_10_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_10_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_11 s_axi__buffered_sourceBuffer_11(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(64'h0000000000000000),
		.io_enq_bits_strb(8'h00),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_3_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_11_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_11_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_11_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_11_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_11 s_axi__buffered_sinkBuffer_7(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_7_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_3_valid)
	);
	Queue2_ReadAddressChannel_10 m_axi__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_enq_valid(_read_arbiter_io_sink_valid),
		.io_enq_bits_id(_read_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_read_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_read_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_read_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_id(m_axi_ar_bits_id),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	Queue2_ReadDataChannel_15 m_axi__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_r_ready),
		.io_enq_valid(m_axi_r_valid),
		.io_enq_bits_id(m_axi_r_bits_id),
		.io_enq_bits_data(m_axi_r_bits_data),
		.io_enq_bits_resp(m_axi_r_bits_resp),
		.io_enq_bits_last(m_axi_r_bits_last),
		.io_deq_ready(m_axi__r_ready),
		.io_deq_valid(_m_axi__sinkBuffer_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_deq_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_deq_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_deq_bits_last(_m_axi__sinkBuffer_io_deq_bits_last)
	);
	Queue2_WriteAddressChannel_10 m_axi__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_sink_valid),
		.io_enq_bits_id(_write_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_write_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_write_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_write_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_id(m_axi_aw_bits_id),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_WriteDataChannel_11 m_axi__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_enq_valid(_write_mux_io_sink_valid),
		.io_enq_bits_data(_write_mux_io_sink_bits_data),
		.io_enq_bits_strb(_write_mux_io_sink_bits_strb),
		.io_enq_bits_last(_write_mux_io_sink_bits_last),
		.io_deq_ready(m_axi_w_ready),
		.io_deq_valid(m_axi_w_valid),
		.io_deq_bits_data(m_axi_w_bits_data),
		.io_deq_bits_strb(m_axi_w_bits_strb),
		.io_deq_bits_last(m_axi_w_bits_last)
	);
	Queue2_WriteResponseChannel_15 m_axi__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_b_ready),
		.io_enq_valid(m_axi_b_valid),
		.io_enq_bits_id(m_axi_b_bits_id),
		.io_enq_bits_resp(m_axi_b_bits_resp),
		.io_deq_ready(m_axi__b_ready),
		.io_deq_valid(_m_axi__sinkBuffer_1_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_1_io_deq_bits_id)
	);
	elasticArbiter_4 read_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_read_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_sources_0_bits_id({2'h0, _s_axi__buffered_sourceBuffer_io_deq_bits_id}),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region),
		.io_sources_1_ready(_read_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_sources_1_bits_id({2'h1, _s_axi__buffered_sourceBuffer_3_io_deq_bits_id}),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region),
		.io_sources_2_ready(_read_arbiter_io_sources_2_ready),
		.io_sources_2_valid(_s_axi__buffered_sourceBuffer_6_io_deq_valid),
		.io_sources_2_bits_id({2'h2, _s_axi__buffered_sourceBuffer_6_io_deq_bits_id}),
		.io_sources_2_bits_addr(_s_axi__buffered_sourceBuffer_6_io_deq_bits_addr),
		.io_sources_2_bits_len(_s_axi__buffered_sourceBuffer_6_io_deq_bits_len),
		.io_sources_2_bits_size(_s_axi__buffered_sourceBuffer_6_io_deq_bits_size),
		.io_sources_2_bits_burst(_s_axi__buffered_sourceBuffer_6_io_deq_bits_burst),
		.io_sources_2_bits_lock(_s_axi__buffered_sourceBuffer_6_io_deq_bits_lock),
		.io_sources_2_bits_cache(_s_axi__buffered_sourceBuffer_6_io_deq_bits_cache),
		.io_sources_2_bits_prot(_s_axi__buffered_sourceBuffer_6_io_deq_bits_prot),
		.io_sources_2_bits_qos(_s_axi__buffered_sourceBuffer_6_io_deq_bits_qos),
		.io_sources_2_bits_region(_s_axi__buffered_sourceBuffer_6_io_deq_bits_region),
		.io_sources_3_ready(_read_arbiter_io_sources_3_ready),
		.io_sources_3_valid(_s_axi__buffered_sourceBuffer_9_io_deq_valid),
		.io_sources_3_bits_id({2'h3, _s_axi__buffered_sourceBuffer_9_io_deq_bits_id}),
		.io_sources_3_bits_addr(_s_axi__buffered_sourceBuffer_9_io_deq_bits_addr),
		.io_sources_3_bits_len(_s_axi__buffered_sourceBuffer_9_io_deq_bits_len),
		.io_sources_3_bits_size(_s_axi__buffered_sourceBuffer_9_io_deq_bits_size),
		.io_sources_3_bits_burst(_s_axi__buffered_sourceBuffer_9_io_deq_bits_burst),
		.io_sources_3_bits_lock(_s_axi__buffered_sourceBuffer_9_io_deq_bits_lock),
		.io_sources_3_bits_cache(_s_axi__buffered_sourceBuffer_9_io_deq_bits_cache),
		.io_sources_3_bits_prot(_s_axi__buffered_sourceBuffer_9_io_deq_bits_prot),
		.io_sources_3_bits_qos(_s_axi__buffered_sourceBuffer_9_io_deq_bits_qos),
		.io_sources_3_bits_region(_s_axi__buffered_sourceBuffer_9_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_sink_valid(_read_arbiter_io_sink_valid),
		.io_sink_bits_id(_read_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_read_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_read_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_read_arbiter_io_sink_bits_region),
		.io_select_ready(1'h1),
		.io_select_valid(),
		.io_select_bits()
	);
	elasticDemux_7 read_demux(
		.io_source_ready(_read_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_0),
		.io_source_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_source_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_source_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_source_bits_last(_m_axi__sinkBuffer_io_deq_bits_last),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_sinks_0_valid(_read_demux_io_sinks_0_valid),
		.io_sinks_0_bits_id(_read_demux_io_sinks_0_bits_id),
		.io_sinks_0_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_sinks_0_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_sinks_0_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_sinks_1_valid(_read_demux_io_sinks_1_valid),
		.io_sinks_1_bits_id(_read_demux_io_sinks_1_bits_id),
		.io_sinks_1_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_sinks_1_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_sinks_1_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_sinks_2_ready(_s_axi__buffered_sinkBuffer_4_io_enq_ready),
		.io_sinks_2_valid(_read_demux_io_sinks_2_valid),
		.io_sinks_2_bits_id(_read_demux_io_sinks_2_bits_id),
		.io_sinks_2_bits_data(_read_demux_io_sinks_2_bits_data),
		.io_sinks_2_bits_resp(_read_demux_io_sinks_2_bits_resp),
		.io_sinks_2_bits_last(_read_demux_io_sinks_2_bits_last),
		.io_sinks_3_ready(_s_axi__buffered_sinkBuffer_6_io_enq_ready),
		.io_sinks_3_valid(_read_demux_io_sinks_3_valid),
		.io_sinks_3_bits_id(_read_demux_io_sinks_3_bits_id),
		.io_sinks_3_bits_data(_read_demux_io_sinks_3_bits_data),
		.io_sinks_3_bits_resp(_read_demux_io_sinks_3_bits_resp),
		.io_sinks_3_bits_last(_read_demux_io_sinks_3_bits_last),
		.io_select_ready(_read_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_io_deq_bits_id[2:1])
	);
	Queue32_UInt2 write_portQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueue_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_select_valid),
		.io_enq_bits(_write_arbiter_io_select_bits),
		.io_deq_ready(_write_mux_io_select_ready),
		.io_deq_valid(_write_portQueue_io_deq_valid),
		.io_deq_bits(_write_portQueue_io_deq_bits)
	);
	elasticArbiter_4 write_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_write_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_sources_0_bits_id({2'h0, _s_axi__buffered_sourceBuffer_1_io_deq_bits_id}),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region),
		.io_sources_1_ready(_write_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_sources_1_bits_id({2'h1, _s_axi__buffered_sourceBuffer_4_io_deq_bits_id}),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region),
		.io_sources_2_ready(_write_arbiter_io_sources_2_ready),
		.io_sources_2_valid(_s_axi__buffered_sourceBuffer_7_io_deq_valid),
		.io_sources_2_bits_id({2'h2, _s_axi__buffered_sourceBuffer_7_io_deq_bits_id}),
		.io_sources_2_bits_addr(_s_axi__buffered_sourceBuffer_7_io_deq_bits_addr),
		.io_sources_2_bits_len(_s_axi__buffered_sourceBuffer_7_io_deq_bits_len),
		.io_sources_2_bits_size(_s_axi__buffered_sourceBuffer_7_io_deq_bits_size),
		.io_sources_2_bits_burst(_s_axi__buffered_sourceBuffer_7_io_deq_bits_burst),
		.io_sources_2_bits_lock(_s_axi__buffered_sourceBuffer_7_io_deq_bits_lock),
		.io_sources_2_bits_cache(_s_axi__buffered_sourceBuffer_7_io_deq_bits_cache),
		.io_sources_2_bits_prot(_s_axi__buffered_sourceBuffer_7_io_deq_bits_prot),
		.io_sources_2_bits_qos(_s_axi__buffered_sourceBuffer_7_io_deq_bits_qos),
		.io_sources_2_bits_region(_s_axi__buffered_sourceBuffer_7_io_deq_bits_region),
		.io_sources_3_ready(_write_arbiter_io_sources_3_ready),
		.io_sources_3_valid(_s_axi__buffered_sourceBuffer_10_io_deq_valid),
		.io_sources_3_bits_id({2'h3, _s_axi__buffered_sourceBuffer_10_io_deq_bits_id}),
		.io_sources_3_bits_addr(_s_axi__buffered_sourceBuffer_10_io_deq_bits_addr),
		.io_sources_3_bits_len(_s_axi__buffered_sourceBuffer_10_io_deq_bits_len),
		.io_sources_3_bits_size(_s_axi__buffered_sourceBuffer_10_io_deq_bits_size),
		.io_sources_3_bits_burst(_s_axi__buffered_sourceBuffer_10_io_deq_bits_burst),
		.io_sources_3_bits_lock(_s_axi__buffered_sourceBuffer_10_io_deq_bits_lock),
		.io_sources_3_bits_cache(_s_axi__buffered_sourceBuffer_10_io_deq_bits_cache),
		.io_sources_3_bits_prot(_s_axi__buffered_sourceBuffer_10_io_deq_bits_prot),
		.io_sources_3_bits_qos(_s_axi__buffered_sourceBuffer_10_io_deq_bits_qos),
		.io_sources_3_bits_region(_s_axi__buffered_sourceBuffer_10_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_sink_valid(_write_arbiter_io_sink_valid),
		.io_sink_bits_id(_write_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_write_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_write_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_write_arbiter_io_sink_bits_region),
		.io_select_ready(_write_portQueue_io_enq_ready),
		.io_select_valid(_write_arbiter_io_select_valid),
		.io_select_bits(_write_arbiter_io_select_bits)
	);
	elasticMux_4 write_mux(
		.io_sources_0_ready(_write_mux_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_sources_0_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_sources_0_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_sources_0_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last),
		.io_sources_1_ready(_write_mux_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_sources_1_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_sources_1_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_sources_1_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last),
		.io_sources_2_ready(_write_mux_io_sources_2_ready),
		.io_sources_2_valid(_s_axi__buffered_sourceBuffer_8_io_deq_valid),
		.io_sources_2_bits_data(_s_axi__buffered_sourceBuffer_8_io_deq_bits_data),
		.io_sources_2_bits_strb(_s_axi__buffered_sourceBuffer_8_io_deq_bits_strb),
		.io_sources_2_bits_last(_s_axi__buffered_sourceBuffer_8_io_deq_bits_last),
		.io_sources_3_ready(_write_mux_io_sources_3_ready),
		.io_sources_3_valid(_s_axi__buffered_sourceBuffer_11_io_deq_valid),
		.io_sources_3_bits_data(_s_axi__buffered_sourceBuffer_11_io_deq_bits_data),
		.io_sources_3_bits_strb(_s_axi__buffered_sourceBuffer_11_io_deq_bits_strb),
		.io_sources_3_bits_last(_s_axi__buffered_sourceBuffer_11_io_deq_bits_last),
		.io_sink_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_sink_valid(_write_mux_io_sink_valid),
		.io_sink_bits_data(_write_mux_io_sink_bits_data),
		.io_sink_bits_strb(_write_mux_io_sink_bits_strb),
		.io_sink_bits_last(_write_mux_io_sink_bits_last),
		.io_select_ready(_write_mux_io_select_ready),
		.io_select_valid(_write_portQueue_io_deq_valid),
		.io_select_bits(_write_portQueue_io_deq_bits)
	);
	elasticDemux_8 write_demux(
		.io_source_ready(_write_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_0),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_sinks_0_valid(_write_demux_io_sinks_0_valid),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_sinks_1_valid(_write_demux_io_sinks_1_valid),
		.io_sinks_2_ready(_s_axi__buffered_sinkBuffer_5_io_enq_ready),
		.io_sinks_2_valid(_write_demux_io_sinks_2_valid),
		.io_sinks_3_ready(_s_axi__buffered_sinkBuffer_7_io_enq_ready),
		.io_sinks_3_valid(_write_demux_io_sinks_3_valid),
		.io_select_ready(_write_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_1_io_deq_bits_id[2:1])
	);
endmodule
module AxisDataWidthConverter_192 (
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [63:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [63:0] io_dataOut_TDATA;
	assign io_dataIn_TREADY = io_dataOut_TREADY;
	assign io_dataOut_TVALID = io_dataIn_TVALID;
	assign io_dataOut_TDATA = io_dataIn_TDATA;
endmodule
module Allocator (
	clock,
	reset,
	io_export_closureOut_0_TREADY,
	io_export_closureOut_0_TVALID,
	io_export_closureOut_0_TDATA,
	io_export_closureOut_1_TREADY,
	io_export_closureOut_1_TVALID,
	io_export_closureOut_1_TDATA,
	io_export_closureOut_2_TREADY,
	io_export_closureOut_2_TVALID,
	io_export_closureOut_2_TDATA,
	io_export_closureOut_3_TREADY,
	io_export_closureOut_3_TVALID,
	io_export_closureOut_3_TDATA,
	io_export_closureOut_4_TREADY,
	io_export_closureOut_4_TVALID,
	io_export_closureOut_4_TDATA,
	io_export_closureOut_5_TREADY,
	io_export_closureOut_5_TVALID,
	io_export_closureOut_5_TDATA,
	io_export_closureOut_6_TREADY,
	io_export_closureOut_6_TVALID,
	io_export_closureOut_6_TDATA,
	io_export_closureOut_7_TREADY,
	io_export_closureOut_7_TVALID,
	io_export_closureOut_7_TDATA,
	io_export_closureOut_8_TREADY,
	io_export_closureOut_8_TVALID,
	io_export_closureOut_8_TDATA,
	io_export_closureOut_9_TREADY,
	io_export_closureOut_9_TVALID,
	io_export_closureOut_9_TDATA,
	io_export_closureOut_10_TREADY,
	io_export_closureOut_10_TVALID,
	io_export_closureOut_10_TDATA,
	io_export_closureOut_11_TREADY,
	io_export_closureOut_11_TVALID,
	io_export_closureOut_11_TDATA,
	io_export_closureOut_12_TREADY,
	io_export_closureOut_12_TVALID,
	io_export_closureOut_12_TDATA,
	io_export_closureOut_13_TREADY,
	io_export_closureOut_13_TVALID,
	io_export_closureOut_13_TDATA,
	io_export_closureOut_14_TREADY,
	io_export_closureOut_14_TVALID,
	io_export_closureOut_14_TDATA,
	io_export_closureOut_15_TREADY,
	io_export_closureOut_15_TVALID,
	io_export_closureOut_15_TDATA,
	io_export_closureOut_16_TREADY,
	io_export_closureOut_16_TVALID,
	io_export_closureOut_16_TDATA,
	io_export_closureOut_17_TREADY,
	io_export_closureOut_17_TVALID,
	io_export_closureOut_17_TDATA,
	io_export_closureOut_18_TREADY,
	io_export_closureOut_18_TVALID,
	io_export_closureOut_18_TDATA,
	io_export_closureOut_19_TREADY,
	io_export_closureOut_19_TVALID,
	io_export_closureOut_19_TDATA,
	io_export_closureOut_20_TREADY,
	io_export_closureOut_20_TVALID,
	io_export_closureOut_20_TDATA,
	io_export_closureOut_21_TREADY,
	io_export_closureOut_21_TVALID,
	io_export_closureOut_21_TDATA,
	io_export_closureOut_22_TREADY,
	io_export_closureOut_22_TVALID,
	io_export_closureOut_22_TDATA,
	io_export_closureOut_23_TREADY,
	io_export_closureOut_23_TVALID,
	io_export_closureOut_23_TDATA,
	io_export_closureOut_24_TREADY,
	io_export_closureOut_24_TVALID,
	io_export_closureOut_24_TDATA,
	io_export_closureOut_25_TREADY,
	io_export_closureOut_25_TVALID,
	io_export_closureOut_25_TDATA,
	io_export_closureOut_26_TREADY,
	io_export_closureOut_26_TVALID,
	io_export_closureOut_26_TDATA,
	io_export_closureOut_27_TREADY,
	io_export_closureOut_27_TVALID,
	io_export_closureOut_27_TDATA,
	io_export_closureOut_28_TREADY,
	io_export_closureOut_28_TVALID,
	io_export_closureOut_28_TDATA,
	io_export_closureOut_29_TREADY,
	io_export_closureOut_29_TVALID,
	io_export_closureOut_29_TDATA,
	io_export_closureOut_30_TREADY,
	io_export_closureOut_30_TVALID,
	io_export_closureOut_30_TDATA,
	io_export_closureOut_31_TREADY,
	io_export_closureOut_31_TVALID,
	io_export_closureOut_31_TDATA,
	io_export_closureOut_32_TREADY,
	io_export_closureOut_32_TVALID,
	io_export_closureOut_32_TDATA,
	io_export_closureOut_33_TREADY,
	io_export_closureOut_33_TVALID,
	io_export_closureOut_33_TDATA,
	io_export_closureOut_34_TREADY,
	io_export_closureOut_34_TVALID,
	io_export_closureOut_34_TDATA,
	io_export_closureOut_35_TREADY,
	io_export_closureOut_35_TVALID,
	io_export_closureOut_35_TDATA,
	io_export_closureOut_36_TREADY,
	io_export_closureOut_36_TVALID,
	io_export_closureOut_36_TDATA,
	io_export_closureOut_37_TREADY,
	io_export_closureOut_37_TVALID,
	io_export_closureOut_37_TDATA,
	io_export_closureOut_38_TREADY,
	io_export_closureOut_38_TVALID,
	io_export_closureOut_38_TDATA,
	io_export_closureOut_39_TREADY,
	io_export_closureOut_39_TVALID,
	io_export_closureOut_39_TDATA,
	io_export_closureOut_40_TREADY,
	io_export_closureOut_40_TVALID,
	io_export_closureOut_40_TDATA,
	io_export_closureOut_41_TREADY,
	io_export_closureOut_41_TVALID,
	io_export_closureOut_41_TDATA,
	io_export_closureOut_42_TREADY,
	io_export_closureOut_42_TVALID,
	io_export_closureOut_42_TDATA,
	io_export_closureOut_43_TREADY,
	io_export_closureOut_43_TVALID,
	io_export_closureOut_43_TDATA,
	io_export_closureOut_44_TREADY,
	io_export_closureOut_44_TVALID,
	io_export_closureOut_44_TDATA,
	io_export_closureOut_45_TREADY,
	io_export_closureOut_45_TVALID,
	io_export_closureOut_45_TDATA,
	io_export_closureOut_46_TREADY,
	io_export_closureOut_46_TVALID,
	io_export_closureOut_46_TDATA,
	io_export_closureOut_47_TREADY,
	io_export_closureOut_47_TVALID,
	io_export_closureOut_47_TDATA,
	io_export_closureOut_48_TREADY,
	io_export_closureOut_48_TVALID,
	io_export_closureOut_48_TDATA,
	io_export_closureOut_49_TREADY,
	io_export_closureOut_49_TVALID,
	io_export_closureOut_49_TDATA,
	io_export_closureOut_50_TREADY,
	io_export_closureOut_50_TVALID,
	io_export_closureOut_50_TDATA,
	io_export_closureOut_51_TREADY,
	io_export_closureOut_51_TVALID,
	io_export_closureOut_51_TDATA,
	io_export_closureOut_52_TREADY,
	io_export_closureOut_52_TVALID,
	io_export_closureOut_52_TDATA,
	io_export_closureOut_53_TREADY,
	io_export_closureOut_53_TVALID,
	io_export_closureOut_53_TDATA,
	io_export_closureOut_54_TREADY,
	io_export_closureOut_54_TVALID,
	io_export_closureOut_54_TDATA,
	io_export_closureOut_55_TREADY,
	io_export_closureOut_55_TVALID,
	io_export_closureOut_55_TDATA,
	io_export_closureOut_56_TREADY,
	io_export_closureOut_56_TVALID,
	io_export_closureOut_56_TDATA,
	io_export_closureOut_57_TREADY,
	io_export_closureOut_57_TVALID,
	io_export_closureOut_57_TDATA,
	io_export_closureOut_58_TREADY,
	io_export_closureOut_58_TVALID,
	io_export_closureOut_58_TDATA,
	io_export_closureOut_59_TREADY,
	io_export_closureOut_59_TVALID,
	io_export_closureOut_59_TDATA,
	io_export_closureOut_60_TREADY,
	io_export_closureOut_60_TVALID,
	io_export_closureOut_60_TDATA,
	io_export_closureOut_61_TREADY,
	io_export_closureOut_61_TVALID,
	io_export_closureOut_61_TDATA,
	io_export_closureOut_62_TREADY,
	io_export_closureOut_62_TVALID,
	io_export_closureOut_62_TDATA,
	io_export_closureOut_63_TREADY,
	io_export_closureOut_63_TVALID,
	io_export_closureOut_63_TDATA,
	io_internal_vcas_axi_full_0_ar_ready,
	io_internal_vcas_axi_full_0_ar_valid,
	io_internal_vcas_axi_full_0_ar_bits_id,
	io_internal_vcas_axi_full_0_ar_bits_addr,
	io_internal_vcas_axi_full_0_ar_bits_len,
	io_internal_vcas_axi_full_0_ar_bits_size,
	io_internal_vcas_axi_full_0_ar_bits_burst,
	io_internal_vcas_axi_full_0_ar_bits_lock,
	io_internal_vcas_axi_full_0_ar_bits_cache,
	io_internal_vcas_axi_full_0_ar_bits_prot,
	io_internal_vcas_axi_full_0_ar_bits_qos,
	io_internal_vcas_axi_full_0_ar_bits_region,
	io_internal_vcas_axi_full_0_r_ready,
	io_internal_vcas_axi_full_0_r_valid,
	io_internal_vcas_axi_full_0_r_bits_id,
	io_internal_vcas_axi_full_0_r_bits_data,
	io_internal_vcas_axi_full_0_r_bits_resp,
	io_internal_vcas_axi_full_0_r_bits_last,
	io_internal_vcas_axi_full_0_aw_ready,
	io_internal_vcas_axi_full_0_aw_valid,
	io_internal_vcas_axi_full_0_aw_bits_id,
	io_internal_vcas_axi_full_0_aw_bits_addr,
	io_internal_vcas_axi_full_0_aw_bits_len,
	io_internal_vcas_axi_full_0_aw_bits_size,
	io_internal_vcas_axi_full_0_aw_bits_burst,
	io_internal_vcas_axi_full_0_aw_bits_lock,
	io_internal_vcas_axi_full_0_aw_bits_cache,
	io_internal_vcas_axi_full_0_aw_bits_prot,
	io_internal_vcas_axi_full_0_aw_bits_qos,
	io_internal_vcas_axi_full_0_aw_bits_region,
	io_internal_vcas_axi_full_0_w_ready,
	io_internal_vcas_axi_full_0_w_valid,
	io_internal_vcas_axi_full_0_w_bits_data,
	io_internal_vcas_axi_full_0_w_bits_strb,
	io_internal_vcas_axi_full_0_w_bits_last,
	io_internal_vcas_axi_full_0_b_ready,
	io_internal_vcas_axi_full_0_b_valid,
	io_internal_vcas_axi_full_0_b_bits_id,
	io_internal_vcas_axi_full_0_b_bits_resp,
	io_internal_axi_mgmt_vcas_0_ar_ready,
	io_internal_axi_mgmt_vcas_0_ar_valid,
	io_internal_axi_mgmt_vcas_0_ar_bits_addr,
	io_internal_axi_mgmt_vcas_0_ar_bits_prot,
	io_internal_axi_mgmt_vcas_0_r_ready,
	io_internal_axi_mgmt_vcas_0_r_valid,
	io_internal_axi_mgmt_vcas_0_r_bits_data,
	io_internal_axi_mgmt_vcas_0_r_bits_resp,
	io_internal_axi_mgmt_vcas_0_aw_ready,
	io_internal_axi_mgmt_vcas_0_aw_valid,
	io_internal_axi_mgmt_vcas_0_aw_bits_addr,
	io_internal_axi_mgmt_vcas_0_aw_bits_prot,
	io_internal_axi_mgmt_vcas_0_w_ready,
	io_internal_axi_mgmt_vcas_0_w_valid,
	io_internal_axi_mgmt_vcas_0_w_bits_data,
	io_internal_axi_mgmt_vcas_0_w_bits_strb,
	io_internal_axi_mgmt_vcas_0_b_ready,
	io_internal_axi_mgmt_vcas_0_b_valid,
	io_internal_axi_mgmt_vcas_0_b_bits_resp,
	io_internal_axi_mgmt_vcas_1_ar_ready,
	io_internal_axi_mgmt_vcas_1_ar_valid,
	io_internal_axi_mgmt_vcas_1_ar_bits_addr,
	io_internal_axi_mgmt_vcas_1_ar_bits_prot,
	io_internal_axi_mgmt_vcas_1_r_ready,
	io_internal_axi_mgmt_vcas_1_r_valid,
	io_internal_axi_mgmt_vcas_1_r_bits_data,
	io_internal_axi_mgmt_vcas_1_r_bits_resp,
	io_internal_axi_mgmt_vcas_1_aw_ready,
	io_internal_axi_mgmt_vcas_1_aw_valid,
	io_internal_axi_mgmt_vcas_1_aw_bits_addr,
	io_internal_axi_mgmt_vcas_1_aw_bits_prot,
	io_internal_axi_mgmt_vcas_1_w_ready,
	io_internal_axi_mgmt_vcas_1_w_valid,
	io_internal_axi_mgmt_vcas_1_w_bits_data,
	io_internal_axi_mgmt_vcas_1_w_bits_strb,
	io_internal_axi_mgmt_vcas_1_b_ready,
	io_internal_axi_mgmt_vcas_1_b_valid,
	io_internal_axi_mgmt_vcas_1_b_bits_resp,
	io_internal_axi_mgmt_vcas_2_ar_ready,
	io_internal_axi_mgmt_vcas_2_ar_valid,
	io_internal_axi_mgmt_vcas_2_ar_bits_addr,
	io_internal_axi_mgmt_vcas_2_ar_bits_prot,
	io_internal_axi_mgmt_vcas_2_r_ready,
	io_internal_axi_mgmt_vcas_2_r_valid,
	io_internal_axi_mgmt_vcas_2_r_bits_data,
	io_internal_axi_mgmt_vcas_2_r_bits_resp,
	io_internal_axi_mgmt_vcas_2_aw_ready,
	io_internal_axi_mgmt_vcas_2_aw_valid,
	io_internal_axi_mgmt_vcas_2_aw_bits_addr,
	io_internal_axi_mgmt_vcas_2_aw_bits_prot,
	io_internal_axi_mgmt_vcas_2_w_ready,
	io_internal_axi_mgmt_vcas_2_w_valid,
	io_internal_axi_mgmt_vcas_2_w_bits_data,
	io_internal_axi_mgmt_vcas_2_w_bits_strb,
	io_internal_axi_mgmt_vcas_2_b_ready,
	io_internal_axi_mgmt_vcas_2_b_valid,
	io_internal_axi_mgmt_vcas_2_b_bits_resp,
	io_internal_axi_mgmt_vcas_3_ar_ready,
	io_internal_axi_mgmt_vcas_3_ar_valid,
	io_internal_axi_mgmt_vcas_3_ar_bits_addr,
	io_internal_axi_mgmt_vcas_3_ar_bits_prot,
	io_internal_axi_mgmt_vcas_3_r_ready,
	io_internal_axi_mgmt_vcas_3_r_valid,
	io_internal_axi_mgmt_vcas_3_r_bits_data,
	io_internal_axi_mgmt_vcas_3_r_bits_resp,
	io_internal_axi_mgmt_vcas_3_aw_ready,
	io_internal_axi_mgmt_vcas_3_aw_valid,
	io_internal_axi_mgmt_vcas_3_aw_bits_addr,
	io_internal_axi_mgmt_vcas_3_aw_bits_prot,
	io_internal_axi_mgmt_vcas_3_w_ready,
	io_internal_axi_mgmt_vcas_3_w_valid,
	io_internal_axi_mgmt_vcas_3_w_bits_data,
	io_internal_axi_mgmt_vcas_3_w_bits_strb,
	io_internal_axi_mgmt_vcas_3_b_ready,
	io_internal_axi_mgmt_vcas_3_b_valid,
	io_internal_axi_mgmt_vcas_3_b_bits_resp
);
	input clock;
	input reset;
	input io_export_closureOut_0_TREADY;
	output wire io_export_closureOut_0_TVALID;
	output wire [63:0] io_export_closureOut_0_TDATA;
	input io_export_closureOut_1_TREADY;
	output wire io_export_closureOut_1_TVALID;
	output wire [63:0] io_export_closureOut_1_TDATA;
	input io_export_closureOut_2_TREADY;
	output wire io_export_closureOut_2_TVALID;
	output wire [63:0] io_export_closureOut_2_TDATA;
	input io_export_closureOut_3_TREADY;
	output wire io_export_closureOut_3_TVALID;
	output wire [63:0] io_export_closureOut_3_TDATA;
	input io_export_closureOut_4_TREADY;
	output wire io_export_closureOut_4_TVALID;
	output wire [63:0] io_export_closureOut_4_TDATA;
	input io_export_closureOut_5_TREADY;
	output wire io_export_closureOut_5_TVALID;
	output wire [63:0] io_export_closureOut_5_TDATA;
	input io_export_closureOut_6_TREADY;
	output wire io_export_closureOut_6_TVALID;
	output wire [63:0] io_export_closureOut_6_TDATA;
	input io_export_closureOut_7_TREADY;
	output wire io_export_closureOut_7_TVALID;
	output wire [63:0] io_export_closureOut_7_TDATA;
	input io_export_closureOut_8_TREADY;
	output wire io_export_closureOut_8_TVALID;
	output wire [63:0] io_export_closureOut_8_TDATA;
	input io_export_closureOut_9_TREADY;
	output wire io_export_closureOut_9_TVALID;
	output wire [63:0] io_export_closureOut_9_TDATA;
	input io_export_closureOut_10_TREADY;
	output wire io_export_closureOut_10_TVALID;
	output wire [63:0] io_export_closureOut_10_TDATA;
	input io_export_closureOut_11_TREADY;
	output wire io_export_closureOut_11_TVALID;
	output wire [63:0] io_export_closureOut_11_TDATA;
	input io_export_closureOut_12_TREADY;
	output wire io_export_closureOut_12_TVALID;
	output wire [63:0] io_export_closureOut_12_TDATA;
	input io_export_closureOut_13_TREADY;
	output wire io_export_closureOut_13_TVALID;
	output wire [63:0] io_export_closureOut_13_TDATA;
	input io_export_closureOut_14_TREADY;
	output wire io_export_closureOut_14_TVALID;
	output wire [63:0] io_export_closureOut_14_TDATA;
	input io_export_closureOut_15_TREADY;
	output wire io_export_closureOut_15_TVALID;
	output wire [63:0] io_export_closureOut_15_TDATA;
	input io_export_closureOut_16_TREADY;
	output wire io_export_closureOut_16_TVALID;
	output wire [63:0] io_export_closureOut_16_TDATA;
	input io_export_closureOut_17_TREADY;
	output wire io_export_closureOut_17_TVALID;
	output wire [63:0] io_export_closureOut_17_TDATA;
	input io_export_closureOut_18_TREADY;
	output wire io_export_closureOut_18_TVALID;
	output wire [63:0] io_export_closureOut_18_TDATA;
	input io_export_closureOut_19_TREADY;
	output wire io_export_closureOut_19_TVALID;
	output wire [63:0] io_export_closureOut_19_TDATA;
	input io_export_closureOut_20_TREADY;
	output wire io_export_closureOut_20_TVALID;
	output wire [63:0] io_export_closureOut_20_TDATA;
	input io_export_closureOut_21_TREADY;
	output wire io_export_closureOut_21_TVALID;
	output wire [63:0] io_export_closureOut_21_TDATA;
	input io_export_closureOut_22_TREADY;
	output wire io_export_closureOut_22_TVALID;
	output wire [63:0] io_export_closureOut_22_TDATA;
	input io_export_closureOut_23_TREADY;
	output wire io_export_closureOut_23_TVALID;
	output wire [63:0] io_export_closureOut_23_TDATA;
	input io_export_closureOut_24_TREADY;
	output wire io_export_closureOut_24_TVALID;
	output wire [63:0] io_export_closureOut_24_TDATA;
	input io_export_closureOut_25_TREADY;
	output wire io_export_closureOut_25_TVALID;
	output wire [63:0] io_export_closureOut_25_TDATA;
	input io_export_closureOut_26_TREADY;
	output wire io_export_closureOut_26_TVALID;
	output wire [63:0] io_export_closureOut_26_TDATA;
	input io_export_closureOut_27_TREADY;
	output wire io_export_closureOut_27_TVALID;
	output wire [63:0] io_export_closureOut_27_TDATA;
	input io_export_closureOut_28_TREADY;
	output wire io_export_closureOut_28_TVALID;
	output wire [63:0] io_export_closureOut_28_TDATA;
	input io_export_closureOut_29_TREADY;
	output wire io_export_closureOut_29_TVALID;
	output wire [63:0] io_export_closureOut_29_TDATA;
	input io_export_closureOut_30_TREADY;
	output wire io_export_closureOut_30_TVALID;
	output wire [63:0] io_export_closureOut_30_TDATA;
	input io_export_closureOut_31_TREADY;
	output wire io_export_closureOut_31_TVALID;
	output wire [63:0] io_export_closureOut_31_TDATA;
	input io_export_closureOut_32_TREADY;
	output wire io_export_closureOut_32_TVALID;
	output wire [63:0] io_export_closureOut_32_TDATA;
	input io_export_closureOut_33_TREADY;
	output wire io_export_closureOut_33_TVALID;
	output wire [63:0] io_export_closureOut_33_TDATA;
	input io_export_closureOut_34_TREADY;
	output wire io_export_closureOut_34_TVALID;
	output wire [63:0] io_export_closureOut_34_TDATA;
	input io_export_closureOut_35_TREADY;
	output wire io_export_closureOut_35_TVALID;
	output wire [63:0] io_export_closureOut_35_TDATA;
	input io_export_closureOut_36_TREADY;
	output wire io_export_closureOut_36_TVALID;
	output wire [63:0] io_export_closureOut_36_TDATA;
	input io_export_closureOut_37_TREADY;
	output wire io_export_closureOut_37_TVALID;
	output wire [63:0] io_export_closureOut_37_TDATA;
	input io_export_closureOut_38_TREADY;
	output wire io_export_closureOut_38_TVALID;
	output wire [63:0] io_export_closureOut_38_TDATA;
	input io_export_closureOut_39_TREADY;
	output wire io_export_closureOut_39_TVALID;
	output wire [63:0] io_export_closureOut_39_TDATA;
	input io_export_closureOut_40_TREADY;
	output wire io_export_closureOut_40_TVALID;
	output wire [63:0] io_export_closureOut_40_TDATA;
	input io_export_closureOut_41_TREADY;
	output wire io_export_closureOut_41_TVALID;
	output wire [63:0] io_export_closureOut_41_TDATA;
	input io_export_closureOut_42_TREADY;
	output wire io_export_closureOut_42_TVALID;
	output wire [63:0] io_export_closureOut_42_TDATA;
	input io_export_closureOut_43_TREADY;
	output wire io_export_closureOut_43_TVALID;
	output wire [63:0] io_export_closureOut_43_TDATA;
	input io_export_closureOut_44_TREADY;
	output wire io_export_closureOut_44_TVALID;
	output wire [63:0] io_export_closureOut_44_TDATA;
	input io_export_closureOut_45_TREADY;
	output wire io_export_closureOut_45_TVALID;
	output wire [63:0] io_export_closureOut_45_TDATA;
	input io_export_closureOut_46_TREADY;
	output wire io_export_closureOut_46_TVALID;
	output wire [63:0] io_export_closureOut_46_TDATA;
	input io_export_closureOut_47_TREADY;
	output wire io_export_closureOut_47_TVALID;
	output wire [63:0] io_export_closureOut_47_TDATA;
	input io_export_closureOut_48_TREADY;
	output wire io_export_closureOut_48_TVALID;
	output wire [63:0] io_export_closureOut_48_TDATA;
	input io_export_closureOut_49_TREADY;
	output wire io_export_closureOut_49_TVALID;
	output wire [63:0] io_export_closureOut_49_TDATA;
	input io_export_closureOut_50_TREADY;
	output wire io_export_closureOut_50_TVALID;
	output wire [63:0] io_export_closureOut_50_TDATA;
	input io_export_closureOut_51_TREADY;
	output wire io_export_closureOut_51_TVALID;
	output wire [63:0] io_export_closureOut_51_TDATA;
	input io_export_closureOut_52_TREADY;
	output wire io_export_closureOut_52_TVALID;
	output wire [63:0] io_export_closureOut_52_TDATA;
	input io_export_closureOut_53_TREADY;
	output wire io_export_closureOut_53_TVALID;
	output wire [63:0] io_export_closureOut_53_TDATA;
	input io_export_closureOut_54_TREADY;
	output wire io_export_closureOut_54_TVALID;
	output wire [63:0] io_export_closureOut_54_TDATA;
	input io_export_closureOut_55_TREADY;
	output wire io_export_closureOut_55_TVALID;
	output wire [63:0] io_export_closureOut_55_TDATA;
	input io_export_closureOut_56_TREADY;
	output wire io_export_closureOut_56_TVALID;
	output wire [63:0] io_export_closureOut_56_TDATA;
	input io_export_closureOut_57_TREADY;
	output wire io_export_closureOut_57_TVALID;
	output wire [63:0] io_export_closureOut_57_TDATA;
	input io_export_closureOut_58_TREADY;
	output wire io_export_closureOut_58_TVALID;
	output wire [63:0] io_export_closureOut_58_TDATA;
	input io_export_closureOut_59_TREADY;
	output wire io_export_closureOut_59_TVALID;
	output wire [63:0] io_export_closureOut_59_TDATA;
	input io_export_closureOut_60_TREADY;
	output wire io_export_closureOut_60_TVALID;
	output wire [63:0] io_export_closureOut_60_TDATA;
	input io_export_closureOut_61_TREADY;
	output wire io_export_closureOut_61_TVALID;
	output wire [63:0] io_export_closureOut_61_TDATA;
	input io_export_closureOut_62_TREADY;
	output wire io_export_closureOut_62_TVALID;
	output wire [63:0] io_export_closureOut_62_TDATA;
	input io_export_closureOut_63_TREADY;
	output wire io_export_closureOut_63_TVALID;
	output wire [63:0] io_export_closureOut_63_TDATA;
	input io_internal_vcas_axi_full_0_ar_ready;
	output wire io_internal_vcas_axi_full_0_ar_valid;
	output wire [6:0] io_internal_vcas_axi_full_0_ar_bits_id;
	output wire [63:0] io_internal_vcas_axi_full_0_ar_bits_addr;
	output wire [7:0] io_internal_vcas_axi_full_0_ar_bits_len;
	output wire [2:0] io_internal_vcas_axi_full_0_ar_bits_size;
	output wire [1:0] io_internal_vcas_axi_full_0_ar_bits_burst;
	output wire io_internal_vcas_axi_full_0_ar_bits_lock;
	output wire [3:0] io_internal_vcas_axi_full_0_ar_bits_cache;
	output wire [2:0] io_internal_vcas_axi_full_0_ar_bits_prot;
	output wire [3:0] io_internal_vcas_axi_full_0_ar_bits_qos;
	output wire [3:0] io_internal_vcas_axi_full_0_ar_bits_region;
	output wire io_internal_vcas_axi_full_0_r_ready;
	input io_internal_vcas_axi_full_0_r_valid;
	input [6:0] io_internal_vcas_axi_full_0_r_bits_id;
	input [63:0] io_internal_vcas_axi_full_0_r_bits_data;
	input [1:0] io_internal_vcas_axi_full_0_r_bits_resp;
	input io_internal_vcas_axi_full_0_r_bits_last;
	input io_internal_vcas_axi_full_0_aw_ready;
	output wire io_internal_vcas_axi_full_0_aw_valid;
	output wire [6:0] io_internal_vcas_axi_full_0_aw_bits_id;
	output wire [63:0] io_internal_vcas_axi_full_0_aw_bits_addr;
	output wire [7:0] io_internal_vcas_axi_full_0_aw_bits_len;
	output wire [2:0] io_internal_vcas_axi_full_0_aw_bits_size;
	output wire [1:0] io_internal_vcas_axi_full_0_aw_bits_burst;
	output wire io_internal_vcas_axi_full_0_aw_bits_lock;
	output wire [3:0] io_internal_vcas_axi_full_0_aw_bits_cache;
	output wire [2:0] io_internal_vcas_axi_full_0_aw_bits_prot;
	output wire [3:0] io_internal_vcas_axi_full_0_aw_bits_qos;
	output wire [3:0] io_internal_vcas_axi_full_0_aw_bits_region;
	input io_internal_vcas_axi_full_0_w_ready;
	output wire io_internal_vcas_axi_full_0_w_valid;
	output wire [63:0] io_internal_vcas_axi_full_0_w_bits_data;
	output wire [7:0] io_internal_vcas_axi_full_0_w_bits_strb;
	output wire io_internal_vcas_axi_full_0_w_bits_last;
	output wire io_internal_vcas_axi_full_0_b_ready;
	input io_internal_vcas_axi_full_0_b_valid;
	input [6:0] io_internal_vcas_axi_full_0_b_bits_id;
	input [1:0] io_internal_vcas_axi_full_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_0_ar_ready;
	input io_internal_axi_mgmt_vcas_0_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_0_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_0_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_0_r_ready;
	output wire io_internal_axi_mgmt_vcas_0_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_0_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_0_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_0_aw_ready;
	input io_internal_axi_mgmt_vcas_0_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_0_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_0_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_0_w_ready;
	input io_internal_axi_mgmt_vcas_0_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_0_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_0_w_bits_strb;
	input io_internal_axi_mgmt_vcas_0_b_ready;
	output wire io_internal_axi_mgmt_vcas_0_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_1_ar_ready;
	input io_internal_axi_mgmt_vcas_1_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_1_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_1_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_1_r_ready;
	output wire io_internal_axi_mgmt_vcas_1_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_1_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_1_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_1_aw_ready;
	input io_internal_axi_mgmt_vcas_1_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_1_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_1_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_1_w_ready;
	input io_internal_axi_mgmt_vcas_1_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_1_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_1_w_bits_strb;
	input io_internal_axi_mgmt_vcas_1_b_ready;
	output wire io_internal_axi_mgmt_vcas_1_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_1_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_2_ar_ready;
	input io_internal_axi_mgmt_vcas_2_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_2_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_2_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_2_r_ready;
	output wire io_internal_axi_mgmt_vcas_2_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_2_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_2_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_2_aw_ready;
	input io_internal_axi_mgmt_vcas_2_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_2_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_2_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_2_w_ready;
	input io_internal_axi_mgmt_vcas_2_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_2_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_2_w_bits_strb;
	input io_internal_axi_mgmt_vcas_2_b_ready;
	output wire io_internal_axi_mgmt_vcas_2_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_2_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_3_ar_ready;
	input io_internal_axi_mgmt_vcas_3_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_3_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_3_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_3_r_ready;
	output wire io_internal_axi_mgmt_vcas_3_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_3_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_3_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_3_aw_ready;
	input io_internal_axi_mgmt_vcas_3_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_3_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_3_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_3_w_ready;
	input io_internal_axi_mgmt_vcas_3_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_3_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_3_w_bits_strb;
	input io_internal_axi_mgmt_vcas_3_b_ready;
	output wire io_internal_axi_mgmt_vcas_3_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_3_b_bits_resp;
	wire _axis_stream_converters_out_63_io_dataIn_TREADY;
	wire _axis_stream_converters_out_62_io_dataIn_TREADY;
	wire _axis_stream_converters_out_61_io_dataIn_TREADY;
	wire _axis_stream_converters_out_60_io_dataIn_TREADY;
	wire _axis_stream_converters_out_59_io_dataIn_TREADY;
	wire _axis_stream_converters_out_58_io_dataIn_TREADY;
	wire _axis_stream_converters_out_57_io_dataIn_TREADY;
	wire _axis_stream_converters_out_56_io_dataIn_TREADY;
	wire _axis_stream_converters_out_55_io_dataIn_TREADY;
	wire _axis_stream_converters_out_54_io_dataIn_TREADY;
	wire _axis_stream_converters_out_53_io_dataIn_TREADY;
	wire _axis_stream_converters_out_52_io_dataIn_TREADY;
	wire _axis_stream_converters_out_51_io_dataIn_TREADY;
	wire _axis_stream_converters_out_50_io_dataIn_TREADY;
	wire _axis_stream_converters_out_49_io_dataIn_TREADY;
	wire _axis_stream_converters_out_48_io_dataIn_TREADY;
	wire _axis_stream_converters_out_47_io_dataIn_TREADY;
	wire _axis_stream_converters_out_46_io_dataIn_TREADY;
	wire _axis_stream_converters_out_45_io_dataIn_TREADY;
	wire _axis_stream_converters_out_44_io_dataIn_TREADY;
	wire _axis_stream_converters_out_43_io_dataIn_TREADY;
	wire _axis_stream_converters_out_42_io_dataIn_TREADY;
	wire _axis_stream_converters_out_41_io_dataIn_TREADY;
	wire _axis_stream_converters_out_40_io_dataIn_TREADY;
	wire _axis_stream_converters_out_39_io_dataIn_TREADY;
	wire _axis_stream_converters_out_38_io_dataIn_TREADY;
	wire _axis_stream_converters_out_37_io_dataIn_TREADY;
	wire _axis_stream_converters_out_36_io_dataIn_TREADY;
	wire _axis_stream_converters_out_35_io_dataIn_TREADY;
	wire _axis_stream_converters_out_34_io_dataIn_TREADY;
	wire _axis_stream_converters_out_33_io_dataIn_TREADY;
	wire _axis_stream_converters_out_32_io_dataIn_TREADY;
	wire _axis_stream_converters_out_31_io_dataIn_TREADY;
	wire _axis_stream_converters_out_30_io_dataIn_TREADY;
	wire _axis_stream_converters_out_29_io_dataIn_TREADY;
	wire _axis_stream_converters_out_28_io_dataIn_TREADY;
	wire _axis_stream_converters_out_27_io_dataIn_TREADY;
	wire _axis_stream_converters_out_26_io_dataIn_TREADY;
	wire _axis_stream_converters_out_25_io_dataIn_TREADY;
	wire _axis_stream_converters_out_24_io_dataIn_TREADY;
	wire _axis_stream_converters_out_23_io_dataIn_TREADY;
	wire _axis_stream_converters_out_22_io_dataIn_TREADY;
	wire _axis_stream_converters_out_21_io_dataIn_TREADY;
	wire _axis_stream_converters_out_20_io_dataIn_TREADY;
	wire _axis_stream_converters_out_19_io_dataIn_TREADY;
	wire _axis_stream_converters_out_18_io_dataIn_TREADY;
	wire _axis_stream_converters_out_17_io_dataIn_TREADY;
	wire _axis_stream_converters_out_16_io_dataIn_TREADY;
	wire _axis_stream_converters_out_15_io_dataIn_TREADY;
	wire _axis_stream_converters_out_14_io_dataIn_TREADY;
	wire _axis_stream_converters_out_13_io_dataIn_TREADY;
	wire _axis_stream_converters_out_12_io_dataIn_TREADY;
	wire _axis_stream_converters_out_11_io_dataIn_TREADY;
	wire _axis_stream_converters_out_10_io_dataIn_TREADY;
	wire _axis_stream_converters_out_9_io_dataIn_TREADY;
	wire _axis_stream_converters_out_8_io_dataIn_TREADY;
	wire _axis_stream_converters_out_7_io_dataIn_TREADY;
	wire _axis_stream_converters_out_6_io_dataIn_TREADY;
	wire _axis_stream_converters_out_5_io_dataIn_TREADY;
	wire _axis_stream_converters_out_4_io_dataIn_TREADY;
	wire _axis_stream_converters_out_3_io_dataIn_TREADY;
	wire _axis_stream_converters_out_2_io_dataIn_TREADY;
	wire _axis_stream_converters_out_1_io_dataIn_TREADY;
	wire _axis_stream_converters_out_0_io_dataIn_TREADY;
	wire _mux_s_axi_0_ar_ready;
	wire _mux_s_axi_0_r_valid;
	wire [63:0] _mux_s_axi_0_r_bits_data;
	wire _mux_s_axi_1_ar_ready;
	wire _mux_s_axi_1_r_valid;
	wire [63:0] _mux_s_axi_1_r_bits_data;
	wire _mux_s_axi_2_ar_ready;
	wire _mux_s_axi_2_r_valid;
	wire [63:0] _mux_s_axi_2_r_bits_data;
	wire _mux_s_axi_3_ar_ready;
	wire _mux_s_axi_3_r_valid;
	wire [63:0] _mux_s_axi_3_r_bits_data;
	wire [2:0] _mux_m_axi_ar_bits_id;
	wire [2:0] _mux_m_axi_aw_bits_id;
	wire _vcasRvmRO_3_io_read_address_ready;
	wire _vcasRvmRO_3_io_read_data_valid;
	wire [63:0] _vcasRvmRO_3_io_read_data_bits;
	wire _vcasRvmRO_3_axi_ar_valid;
	wire [63:0] _vcasRvmRO_3_axi_ar_bits_addr;
	wire _vcasRvmRO_3_axi_r_ready;
	wire _vcasRvmRO_2_io_read_address_ready;
	wire _vcasRvmRO_2_io_read_data_valid;
	wire [63:0] _vcasRvmRO_2_io_read_data_bits;
	wire _vcasRvmRO_2_axi_ar_valid;
	wire [63:0] _vcasRvmRO_2_axi_ar_bits_addr;
	wire _vcasRvmRO_2_axi_r_ready;
	wire _vcasRvmRO_1_io_read_address_ready;
	wire _vcasRvmRO_1_io_read_data_valid;
	wire [63:0] _vcasRvmRO_1_io_read_data_bits;
	wire _vcasRvmRO_1_axi_ar_valid;
	wire [63:0] _vcasRvmRO_1_axi_ar_bits_addr;
	wire _vcasRvmRO_1_axi_r_ready;
	wire _vcasRvmRO_0_io_read_address_ready;
	wire _vcasRvmRO_0_io_read_data_valid;
	wire [63:0] _vcasRvmRO_0_io_read_data_bits;
	wire _vcasRvmRO_0_axi_ar_valid;
	wire [63:0] _vcasRvmRO_0_axi_ar_bits_addr;
	wire _vcasRvmRO_0_axi_r_ready;
	wire _vcas_3_io_dataOut_valid;
	wire [63:0] _vcas_3_io_dataOut_bits;
	wire _vcas_3_io_read_address_valid;
	wire [63:0] _vcas_3_io_read_address_bits;
	wire _vcas_3_io_read_data_ready;
	wire _vcas_2_io_dataOut_valid;
	wire [63:0] _vcas_2_io_dataOut_bits;
	wire _vcas_2_io_read_address_valid;
	wire [63:0] _vcas_2_io_read_address_bits;
	wire _vcas_2_io_read_data_ready;
	wire _vcas_1_io_dataOut_valid;
	wire [63:0] _vcas_1_io_dataOut_bits;
	wire _vcas_1_io_read_address_valid;
	wire [63:0] _vcas_1_io_read_address_bits;
	wire _vcas_1_io_read_data_ready;
	wire _vcas_0_io_dataOut_valid;
	wire [63:0] _vcas_0_io_dataOut_bits;
	wire _vcas_0_io_read_address_valid;
	wire [63:0] _vcas_0_io_read_address_bits;
	wire _vcas_0_io_read_data_ready;
	wire _continuationNetwork_io_connVCAS_0_ready;
	wire _continuationNetwork_io_connVCAS_1_ready;
	wire _continuationNetwork_io_connVCAS_2_ready;
	wire _continuationNetwork_io_connVCAS_3_ready;
	wire _continuationNetwork_io_connPE_0_valid;
	wire [63:0] _continuationNetwork_io_connPE_0_bits;
	wire _continuationNetwork_io_connPE_1_valid;
	wire [63:0] _continuationNetwork_io_connPE_1_bits;
	wire _continuationNetwork_io_connPE_2_valid;
	wire [63:0] _continuationNetwork_io_connPE_2_bits;
	wire _continuationNetwork_io_connPE_3_valid;
	wire [63:0] _continuationNetwork_io_connPE_3_bits;
	wire _continuationNetwork_io_connPE_4_valid;
	wire [63:0] _continuationNetwork_io_connPE_4_bits;
	wire _continuationNetwork_io_connPE_5_valid;
	wire [63:0] _continuationNetwork_io_connPE_5_bits;
	wire _continuationNetwork_io_connPE_6_valid;
	wire [63:0] _continuationNetwork_io_connPE_6_bits;
	wire _continuationNetwork_io_connPE_7_valid;
	wire [63:0] _continuationNetwork_io_connPE_7_bits;
	wire _continuationNetwork_io_connPE_8_valid;
	wire [63:0] _continuationNetwork_io_connPE_8_bits;
	wire _continuationNetwork_io_connPE_9_valid;
	wire [63:0] _continuationNetwork_io_connPE_9_bits;
	wire _continuationNetwork_io_connPE_10_valid;
	wire [63:0] _continuationNetwork_io_connPE_10_bits;
	wire _continuationNetwork_io_connPE_11_valid;
	wire [63:0] _continuationNetwork_io_connPE_11_bits;
	wire _continuationNetwork_io_connPE_12_valid;
	wire [63:0] _continuationNetwork_io_connPE_12_bits;
	wire _continuationNetwork_io_connPE_13_valid;
	wire [63:0] _continuationNetwork_io_connPE_13_bits;
	wire _continuationNetwork_io_connPE_14_valid;
	wire [63:0] _continuationNetwork_io_connPE_14_bits;
	wire _continuationNetwork_io_connPE_15_valid;
	wire [63:0] _continuationNetwork_io_connPE_15_bits;
	wire _continuationNetwork_io_connPE_16_valid;
	wire [63:0] _continuationNetwork_io_connPE_16_bits;
	wire _continuationNetwork_io_connPE_17_valid;
	wire [63:0] _continuationNetwork_io_connPE_17_bits;
	wire _continuationNetwork_io_connPE_18_valid;
	wire [63:0] _continuationNetwork_io_connPE_18_bits;
	wire _continuationNetwork_io_connPE_19_valid;
	wire [63:0] _continuationNetwork_io_connPE_19_bits;
	wire _continuationNetwork_io_connPE_20_valid;
	wire [63:0] _continuationNetwork_io_connPE_20_bits;
	wire _continuationNetwork_io_connPE_21_valid;
	wire [63:0] _continuationNetwork_io_connPE_21_bits;
	wire _continuationNetwork_io_connPE_22_valid;
	wire [63:0] _continuationNetwork_io_connPE_22_bits;
	wire _continuationNetwork_io_connPE_23_valid;
	wire [63:0] _continuationNetwork_io_connPE_23_bits;
	wire _continuationNetwork_io_connPE_24_valid;
	wire [63:0] _continuationNetwork_io_connPE_24_bits;
	wire _continuationNetwork_io_connPE_25_valid;
	wire [63:0] _continuationNetwork_io_connPE_25_bits;
	wire _continuationNetwork_io_connPE_26_valid;
	wire [63:0] _continuationNetwork_io_connPE_26_bits;
	wire _continuationNetwork_io_connPE_27_valid;
	wire [63:0] _continuationNetwork_io_connPE_27_bits;
	wire _continuationNetwork_io_connPE_28_valid;
	wire [63:0] _continuationNetwork_io_connPE_28_bits;
	wire _continuationNetwork_io_connPE_29_valid;
	wire [63:0] _continuationNetwork_io_connPE_29_bits;
	wire _continuationNetwork_io_connPE_30_valid;
	wire [63:0] _continuationNetwork_io_connPE_30_bits;
	wire _continuationNetwork_io_connPE_31_valid;
	wire [63:0] _continuationNetwork_io_connPE_31_bits;
	wire _continuationNetwork_io_connPE_32_valid;
	wire [63:0] _continuationNetwork_io_connPE_32_bits;
	wire _continuationNetwork_io_connPE_33_valid;
	wire [63:0] _continuationNetwork_io_connPE_33_bits;
	wire _continuationNetwork_io_connPE_34_valid;
	wire [63:0] _continuationNetwork_io_connPE_34_bits;
	wire _continuationNetwork_io_connPE_35_valid;
	wire [63:0] _continuationNetwork_io_connPE_35_bits;
	wire _continuationNetwork_io_connPE_36_valid;
	wire [63:0] _continuationNetwork_io_connPE_36_bits;
	wire _continuationNetwork_io_connPE_37_valid;
	wire [63:0] _continuationNetwork_io_connPE_37_bits;
	wire _continuationNetwork_io_connPE_38_valid;
	wire [63:0] _continuationNetwork_io_connPE_38_bits;
	wire _continuationNetwork_io_connPE_39_valid;
	wire [63:0] _continuationNetwork_io_connPE_39_bits;
	wire _continuationNetwork_io_connPE_40_valid;
	wire [63:0] _continuationNetwork_io_connPE_40_bits;
	wire _continuationNetwork_io_connPE_41_valid;
	wire [63:0] _continuationNetwork_io_connPE_41_bits;
	wire _continuationNetwork_io_connPE_42_valid;
	wire [63:0] _continuationNetwork_io_connPE_42_bits;
	wire _continuationNetwork_io_connPE_43_valid;
	wire [63:0] _continuationNetwork_io_connPE_43_bits;
	wire _continuationNetwork_io_connPE_44_valid;
	wire [63:0] _continuationNetwork_io_connPE_44_bits;
	wire _continuationNetwork_io_connPE_45_valid;
	wire [63:0] _continuationNetwork_io_connPE_45_bits;
	wire _continuationNetwork_io_connPE_46_valid;
	wire [63:0] _continuationNetwork_io_connPE_46_bits;
	wire _continuationNetwork_io_connPE_47_valid;
	wire [63:0] _continuationNetwork_io_connPE_47_bits;
	wire _continuationNetwork_io_connPE_48_valid;
	wire [63:0] _continuationNetwork_io_connPE_48_bits;
	wire _continuationNetwork_io_connPE_49_valid;
	wire [63:0] _continuationNetwork_io_connPE_49_bits;
	wire _continuationNetwork_io_connPE_50_valid;
	wire [63:0] _continuationNetwork_io_connPE_50_bits;
	wire _continuationNetwork_io_connPE_51_valid;
	wire [63:0] _continuationNetwork_io_connPE_51_bits;
	wire _continuationNetwork_io_connPE_52_valid;
	wire [63:0] _continuationNetwork_io_connPE_52_bits;
	wire _continuationNetwork_io_connPE_53_valid;
	wire [63:0] _continuationNetwork_io_connPE_53_bits;
	wire _continuationNetwork_io_connPE_54_valid;
	wire [63:0] _continuationNetwork_io_connPE_54_bits;
	wire _continuationNetwork_io_connPE_55_valid;
	wire [63:0] _continuationNetwork_io_connPE_55_bits;
	wire _continuationNetwork_io_connPE_56_valid;
	wire [63:0] _continuationNetwork_io_connPE_56_bits;
	wire _continuationNetwork_io_connPE_57_valid;
	wire [63:0] _continuationNetwork_io_connPE_57_bits;
	wire _continuationNetwork_io_connPE_58_valid;
	wire [63:0] _continuationNetwork_io_connPE_58_bits;
	wire _continuationNetwork_io_connPE_59_valid;
	wire [63:0] _continuationNetwork_io_connPE_59_bits;
	wire _continuationNetwork_io_connPE_60_valid;
	wire [63:0] _continuationNetwork_io_connPE_60_bits;
	wire _continuationNetwork_io_connPE_61_valid;
	wire [63:0] _continuationNetwork_io_connPE_61_bits;
	wire _continuationNetwork_io_connPE_62_valid;
	wire [63:0] _continuationNetwork_io_connPE_62_bits;
	wire _continuationNetwork_io_connPE_63_valid;
	wire [63:0] _continuationNetwork_io_connPE_63_bits;
	AllocatorNetwork continuationNetwork(
		.clock(clock),
		.reset(reset),
		.io_connVCAS_0_ready(_continuationNetwork_io_connVCAS_0_ready),
		.io_connVCAS_0_valid(_vcas_0_io_dataOut_valid),
		.io_connVCAS_0_bits(_vcas_0_io_dataOut_bits),
		.io_connVCAS_1_ready(_continuationNetwork_io_connVCAS_1_ready),
		.io_connVCAS_1_valid(_vcas_1_io_dataOut_valid),
		.io_connVCAS_1_bits(_vcas_1_io_dataOut_bits),
		.io_connVCAS_2_ready(_continuationNetwork_io_connVCAS_2_ready),
		.io_connVCAS_2_valid(_vcas_2_io_dataOut_valid),
		.io_connVCAS_2_bits(_vcas_2_io_dataOut_bits),
		.io_connVCAS_3_ready(_continuationNetwork_io_connVCAS_3_ready),
		.io_connVCAS_3_valid(_vcas_3_io_dataOut_valid),
		.io_connVCAS_3_bits(_vcas_3_io_dataOut_bits),
		.io_connPE_0_ready(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_connPE_0_valid(_continuationNetwork_io_connPE_0_valid),
		.io_connPE_0_bits(_continuationNetwork_io_connPE_0_bits),
		.io_connPE_1_ready(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_connPE_1_valid(_continuationNetwork_io_connPE_1_valid),
		.io_connPE_1_bits(_continuationNetwork_io_connPE_1_bits),
		.io_connPE_2_ready(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_connPE_2_valid(_continuationNetwork_io_connPE_2_valid),
		.io_connPE_2_bits(_continuationNetwork_io_connPE_2_bits),
		.io_connPE_3_ready(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_connPE_3_valid(_continuationNetwork_io_connPE_3_valid),
		.io_connPE_3_bits(_continuationNetwork_io_connPE_3_bits),
		.io_connPE_4_ready(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_connPE_4_valid(_continuationNetwork_io_connPE_4_valid),
		.io_connPE_4_bits(_continuationNetwork_io_connPE_4_bits),
		.io_connPE_5_ready(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_connPE_5_valid(_continuationNetwork_io_connPE_5_valid),
		.io_connPE_5_bits(_continuationNetwork_io_connPE_5_bits),
		.io_connPE_6_ready(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_connPE_6_valid(_continuationNetwork_io_connPE_6_valid),
		.io_connPE_6_bits(_continuationNetwork_io_connPE_6_bits),
		.io_connPE_7_ready(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_connPE_7_valid(_continuationNetwork_io_connPE_7_valid),
		.io_connPE_7_bits(_continuationNetwork_io_connPE_7_bits),
		.io_connPE_8_ready(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_connPE_8_valid(_continuationNetwork_io_connPE_8_valid),
		.io_connPE_8_bits(_continuationNetwork_io_connPE_8_bits),
		.io_connPE_9_ready(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_connPE_9_valid(_continuationNetwork_io_connPE_9_valid),
		.io_connPE_9_bits(_continuationNetwork_io_connPE_9_bits),
		.io_connPE_10_ready(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_connPE_10_valid(_continuationNetwork_io_connPE_10_valid),
		.io_connPE_10_bits(_continuationNetwork_io_connPE_10_bits),
		.io_connPE_11_ready(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_connPE_11_valid(_continuationNetwork_io_connPE_11_valid),
		.io_connPE_11_bits(_continuationNetwork_io_connPE_11_bits),
		.io_connPE_12_ready(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_connPE_12_valid(_continuationNetwork_io_connPE_12_valid),
		.io_connPE_12_bits(_continuationNetwork_io_connPE_12_bits),
		.io_connPE_13_ready(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_connPE_13_valid(_continuationNetwork_io_connPE_13_valid),
		.io_connPE_13_bits(_continuationNetwork_io_connPE_13_bits),
		.io_connPE_14_ready(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_connPE_14_valid(_continuationNetwork_io_connPE_14_valid),
		.io_connPE_14_bits(_continuationNetwork_io_connPE_14_bits),
		.io_connPE_15_ready(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_connPE_15_valid(_continuationNetwork_io_connPE_15_valid),
		.io_connPE_15_bits(_continuationNetwork_io_connPE_15_bits),
		.io_connPE_16_ready(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_connPE_16_valid(_continuationNetwork_io_connPE_16_valid),
		.io_connPE_16_bits(_continuationNetwork_io_connPE_16_bits),
		.io_connPE_17_ready(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_connPE_17_valid(_continuationNetwork_io_connPE_17_valid),
		.io_connPE_17_bits(_continuationNetwork_io_connPE_17_bits),
		.io_connPE_18_ready(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_connPE_18_valid(_continuationNetwork_io_connPE_18_valid),
		.io_connPE_18_bits(_continuationNetwork_io_connPE_18_bits),
		.io_connPE_19_ready(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_connPE_19_valid(_continuationNetwork_io_connPE_19_valid),
		.io_connPE_19_bits(_continuationNetwork_io_connPE_19_bits),
		.io_connPE_20_ready(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_connPE_20_valid(_continuationNetwork_io_connPE_20_valid),
		.io_connPE_20_bits(_continuationNetwork_io_connPE_20_bits),
		.io_connPE_21_ready(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_connPE_21_valid(_continuationNetwork_io_connPE_21_valid),
		.io_connPE_21_bits(_continuationNetwork_io_connPE_21_bits),
		.io_connPE_22_ready(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_connPE_22_valid(_continuationNetwork_io_connPE_22_valid),
		.io_connPE_22_bits(_continuationNetwork_io_connPE_22_bits),
		.io_connPE_23_ready(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_connPE_23_valid(_continuationNetwork_io_connPE_23_valid),
		.io_connPE_23_bits(_continuationNetwork_io_connPE_23_bits),
		.io_connPE_24_ready(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_connPE_24_valid(_continuationNetwork_io_connPE_24_valid),
		.io_connPE_24_bits(_continuationNetwork_io_connPE_24_bits),
		.io_connPE_25_ready(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_connPE_25_valid(_continuationNetwork_io_connPE_25_valid),
		.io_connPE_25_bits(_continuationNetwork_io_connPE_25_bits),
		.io_connPE_26_ready(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_connPE_26_valid(_continuationNetwork_io_connPE_26_valid),
		.io_connPE_26_bits(_continuationNetwork_io_connPE_26_bits),
		.io_connPE_27_ready(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_connPE_27_valid(_continuationNetwork_io_connPE_27_valid),
		.io_connPE_27_bits(_continuationNetwork_io_connPE_27_bits),
		.io_connPE_28_ready(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_connPE_28_valid(_continuationNetwork_io_connPE_28_valid),
		.io_connPE_28_bits(_continuationNetwork_io_connPE_28_bits),
		.io_connPE_29_ready(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_connPE_29_valid(_continuationNetwork_io_connPE_29_valid),
		.io_connPE_29_bits(_continuationNetwork_io_connPE_29_bits),
		.io_connPE_30_ready(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_connPE_30_valid(_continuationNetwork_io_connPE_30_valid),
		.io_connPE_30_bits(_continuationNetwork_io_connPE_30_bits),
		.io_connPE_31_ready(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_connPE_31_valid(_continuationNetwork_io_connPE_31_valid),
		.io_connPE_31_bits(_continuationNetwork_io_connPE_31_bits),
		.io_connPE_32_ready(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_connPE_32_valid(_continuationNetwork_io_connPE_32_valid),
		.io_connPE_32_bits(_continuationNetwork_io_connPE_32_bits),
		.io_connPE_33_ready(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_connPE_33_valid(_continuationNetwork_io_connPE_33_valid),
		.io_connPE_33_bits(_continuationNetwork_io_connPE_33_bits),
		.io_connPE_34_ready(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_connPE_34_valid(_continuationNetwork_io_connPE_34_valid),
		.io_connPE_34_bits(_continuationNetwork_io_connPE_34_bits),
		.io_connPE_35_ready(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_connPE_35_valid(_continuationNetwork_io_connPE_35_valid),
		.io_connPE_35_bits(_continuationNetwork_io_connPE_35_bits),
		.io_connPE_36_ready(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_connPE_36_valid(_continuationNetwork_io_connPE_36_valid),
		.io_connPE_36_bits(_continuationNetwork_io_connPE_36_bits),
		.io_connPE_37_ready(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_connPE_37_valid(_continuationNetwork_io_connPE_37_valid),
		.io_connPE_37_bits(_continuationNetwork_io_connPE_37_bits),
		.io_connPE_38_ready(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_connPE_38_valid(_continuationNetwork_io_connPE_38_valid),
		.io_connPE_38_bits(_continuationNetwork_io_connPE_38_bits),
		.io_connPE_39_ready(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_connPE_39_valid(_continuationNetwork_io_connPE_39_valid),
		.io_connPE_39_bits(_continuationNetwork_io_connPE_39_bits),
		.io_connPE_40_ready(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_connPE_40_valid(_continuationNetwork_io_connPE_40_valid),
		.io_connPE_40_bits(_continuationNetwork_io_connPE_40_bits),
		.io_connPE_41_ready(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_connPE_41_valid(_continuationNetwork_io_connPE_41_valid),
		.io_connPE_41_bits(_continuationNetwork_io_connPE_41_bits),
		.io_connPE_42_ready(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_connPE_42_valid(_continuationNetwork_io_connPE_42_valid),
		.io_connPE_42_bits(_continuationNetwork_io_connPE_42_bits),
		.io_connPE_43_ready(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_connPE_43_valid(_continuationNetwork_io_connPE_43_valid),
		.io_connPE_43_bits(_continuationNetwork_io_connPE_43_bits),
		.io_connPE_44_ready(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_connPE_44_valid(_continuationNetwork_io_connPE_44_valid),
		.io_connPE_44_bits(_continuationNetwork_io_connPE_44_bits),
		.io_connPE_45_ready(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_connPE_45_valid(_continuationNetwork_io_connPE_45_valid),
		.io_connPE_45_bits(_continuationNetwork_io_connPE_45_bits),
		.io_connPE_46_ready(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_connPE_46_valid(_continuationNetwork_io_connPE_46_valid),
		.io_connPE_46_bits(_continuationNetwork_io_connPE_46_bits),
		.io_connPE_47_ready(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_connPE_47_valid(_continuationNetwork_io_connPE_47_valid),
		.io_connPE_47_bits(_continuationNetwork_io_connPE_47_bits),
		.io_connPE_48_ready(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_connPE_48_valid(_continuationNetwork_io_connPE_48_valid),
		.io_connPE_48_bits(_continuationNetwork_io_connPE_48_bits),
		.io_connPE_49_ready(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_connPE_49_valid(_continuationNetwork_io_connPE_49_valid),
		.io_connPE_49_bits(_continuationNetwork_io_connPE_49_bits),
		.io_connPE_50_ready(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_connPE_50_valid(_continuationNetwork_io_connPE_50_valid),
		.io_connPE_50_bits(_continuationNetwork_io_connPE_50_bits),
		.io_connPE_51_ready(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_connPE_51_valid(_continuationNetwork_io_connPE_51_valid),
		.io_connPE_51_bits(_continuationNetwork_io_connPE_51_bits),
		.io_connPE_52_ready(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_connPE_52_valid(_continuationNetwork_io_connPE_52_valid),
		.io_connPE_52_bits(_continuationNetwork_io_connPE_52_bits),
		.io_connPE_53_ready(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_connPE_53_valid(_continuationNetwork_io_connPE_53_valid),
		.io_connPE_53_bits(_continuationNetwork_io_connPE_53_bits),
		.io_connPE_54_ready(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_connPE_54_valid(_continuationNetwork_io_connPE_54_valid),
		.io_connPE_54_bits(_continuationNetwork_io_connPE_54_bits),
		.io_connPE_55_ready(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_connPE_55_valid(_continuationNetwork_io_connPE_55_valid),
		.io_connPE_55_bits(_continuationNetwork_io_connPE_55_bits),
		.io_connPE_56_ready(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_connPE_56_valid(_continuationNetwork_io_connPE_56_valid),
		.io_connPE_56_bits(_continuationNetwork_io_connPE_56_bits),
		.io_connPE_57_ready(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_connPE_57_valid(_continuationNetwork_io_connPE_57_valid),
		.io_connPE_57_bits(_continuationNetwork_io_connPE_57_bits),
		.io_connPE_58_ready(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_connPE_58_valid(_continuationNetwork_io_connPE_58_valid),
		.io_connPE_58_bits(_continuationNetwork_io_connPE_58_bits),
		.io_connPE_59_ready(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_connPE_59_valid(_continuationNetwork_io_connPE_59_valid),
		.io_connPE_59_bits(_continuationNetwork_io_connPE_59_bits),
		.io_connPE_60_ready(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_connPE_60_valid(_continuationNetwork_io_connPE_60_valid),
		.io_connPE_60_bits(_continuationNetwork_io_connPE_60_bits),
		.io_connPE_61_ready(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_connPE_61_valid(_continuationNetwork_io_connPE_61_valid),
		.io_connPE_61_bits(_continuationNetwork_io_connPE_61_bits),
		.io_connPE_62_ready(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_connPE_62_valid(_continuationNetwork_io_connPE_62_valid),
		.io_connPE_62_bits(_continuationNetwork_io_connPE_62_bits),
		.io_connPE_63_ready(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_connPE_63_valid(_continuationNetwork_io_connPE_63_valid),
		.io_connPE_63_bits(_continuationNetwork_io_connPE_63_bits)
	);
	AllocatorServer vcas_0(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_0_ready),
		.io_dataOut_valid(_vcas_0_io_dataOut_valid),
		.io_dataOut_bits(_vcas_0_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_0_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_0_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_0_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_0_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_0_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_0_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_0_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_0_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_0_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_0_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_0_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_0_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_0_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_0_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_0_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_0_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_0_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_0_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_0_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_0_io_read_address_ready),
		.io_read_address_valid(_vcas_0_io_read_address_valid),
		.io_read_address_bits(_vcas_0_io_read_address_bits),
		.io_read_data_ready(_vcas_0_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_0_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_0_io_read_data_bits)
	);
	AllocatorServer vcas_1(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_1_ready),
		.io_dataOut_valid(_vcas_1_io_dataOut_valid),
		.io_dataOut_bits(_vcas_1_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_1_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_1_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_1_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_1_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_1_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_1_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_1_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_1_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_1_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_1_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_1_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_1_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_1_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_1_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_1_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_1_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_1_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_1_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_1_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_1_io_read_address_ready),
		.io_read_address_valid(_vcas_1_io_read_address_valid),
		.io_read_address_bits(_vcas_1_io_read_address_bits),
		.io_read_data_ready(_vcas_1_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_1_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_1_io_read_data_bits)
	);
	AllocatorServer vcas_2(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_2_ready),
		.io_dataOut_valid(_vcas_2_io_dataOut_valid),
		.io_dataOut_bits(_vcas_2_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_2_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_2_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_2_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_2_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_2_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_2_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_2_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_2_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_2_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_2_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_2_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_2_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_2_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_2_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_2_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_2_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_2_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_2_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_2_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_2_io_read_address_ready),
		.io_read_address_valid(_vcas_2_io_read_address_valid),
		.io_read_address_bits(_vcas_2_io_read_address_bits),
		.io_read_data_ready(_vcas_2_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_2_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_2_io_read_data_bits)
	);
	AllocatorServer vcas_3(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_3_ready),
		.io_dataOut_valid(_vcas_3_io_dataOut_valid),
		.io_dataOut_bits(_vcas_3_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_3_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_3_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_3_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_3_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_3_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_3_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_3_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_3_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_3_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_3_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_3_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_3_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_3_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_3_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_3_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_3_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_3_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_3_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_3_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_3_io_read_address_ready),
		.io_read_address_valid(_vcas_3_io_read_address_valid),
		.io_read_address_bits(_vcas_3_io_read_address_bits),
		.io_read_data_ready(_vcas_3_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_3_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_3_io_read_data_bits)
	);
	RVtoAXIBridge_4 vcasRvmRO_0(
		.io_read_address_ready(_vcasRvmRO_0_io_read_address_ready),
		.io_read_address_valid(_vcas_0_io_read_address_valid),
		.io_read_address_bits(_vcas_0_io_read_address_bits),
		.io_read_data_ready(_vcas_0_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_0_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_0_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_0_ar_ready),
		.axi_ar_valid(_vcasRvmRO_0_axi_ar_valid),
		.axi_ar_bits_addr(_vcasRvmRO_0_axi_ar_bits_addr),
		.axi_r_ready(_vcasRvmRO_0_axi_r_ready),
		.axi_r_valid(_mux_s_axi_0_r_valid),
		.axi_r_bits_data(_mux_s_axi_0_r_bits_data)
	);
	RVtoAXIBridge_4 vcasRvmRO_1(
		.io_read_address_ready(_vcasRvmRO_1_io_read_address_ready),
		.io_read_address_valid(_vcas_1_io_read_address_valid),
		.io_read_address_bits(_vcas_1_io_read_address_bits),
		.io_read_data_ready(_vcas_1_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_1_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_1_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_1_ar_ready),
		.axi_ar_valid(_vcasRvmRO_1_axi_ar_valid),
		.axi_ar_bits_addr(_vcasRvmRO_1_axi_ar_bits_addr),
		.axi_r_ready(_vcasRvmRO_1_axi_r_ready),
		.axi_r_valid(_mux_s_axi_1_r_valid),
		.axi_r_bits_data(_mux_s_axi_1_r_bits_data)
	);
	RVtoAXIBridge_4 vcasRvmRO_2(
		.io_read_address_ready(_vcasRvmRO_2_io_read_address_ready),
		.io_read_address_valid(_vcas_2_io_read_address_valid),
		.io_read_address_bits(_vcas_2_io_read_address_bits),
		.io_read_data_ready(_vcas_2_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_2_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_2_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_2_ar_ready),
		.axi_ar_valid(_vcasRvmRO_2_axi_ar_valid),
		.axi_ar_bits_addr(_vcasRvmRO_2_axi_ar_bits_addr),
		.axi_r_ready(_vcasRvmRO_2_axi_r_ready),
		.axi_r_valid(_mux_s_axi_2_r_valid),
		.axi_r_bits_data(_mux_s_axi_2_r_bits_data)
	);
	RVtoAXIBridge_4 vcasRvmRO_3(
		.io_read_address_ready(_vcasRvmRO_3_io_read_address_ready),
		.io_read_address_valid(_vcas_3_io_read_address_valid),
		.io_read_address_bits(_vcas_3_io_read_address_bits),
		.io_read_data_ready(_vcas_3_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_3_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_3_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_3_ar_ready),
		.axi_ar_valid(_vcasRvmRO_3_axi_ar_valid),
		.axi_ar_bits_addr(_vcasRvmRO_3_axi_ar_bits_addr),
		.axi_r_ready(_vcasRvmRO_3_axi_r_ready),
		.axi_r_valid(_mux_s_axi_3_r_valid),
		.axi_r_bits_data(_mux_s_axi_3_r_bits_data)
	);
	axi4FullMux_2 mux(
		.clock(clock),
		.reset(reset),
		.s_axi_0_ar_ready(_mux_s_axi_0_ar_ready),
		.s_axi_0_ar_valid(_vcasRvmRO_0_axi_ar_valid),
		.s_axi_0_ar_bits_addr(_vcasRvmRO_0_axi_ar_bits_addr),
		.s_axi_0_r_ready(_vcasRvmRO_0_axi_r_ready),
		.s_axi_0_r_valid(_mux_s_axi_0_r_valid),
		.s_axi_0_r_bits_data(_mux_s_axi_0_r_bits_data),
		.s_axi_1_ar_ready(_mux_s_axi_1_ar_ready),
		.s_axi_1_ar_valid(_vcasRvmRO_1_axi_ar_valid),
		.s_axi_1_ar_bits_addr(_vcasRvmRO_1_axi_ar_bits_addr),
		.s_axi_1_r_ready(_vcasRvmRO_1_axi_r_ready),
		.s_axi_1_r_valid(_mux_s_axi_1_r_valid),
		.s_axi_1_r_bits_data(_mux_s_axi_1_r_bits_data),
		.s_axi_2_ar_ready(_mux_s_axi_2_ar_ready),
		.s_axi_2_ar_valid(_vcasRvmRO_2_axi_ar_valid),
		.s_axi_2_ar_bits_addr(_vcasRvmRO_2_axi_ar_bits_addr),
		.s_axi_2_r_ready(_vcasRvmRO_2_axi_r_ready),
		.s_axi_2_r_valid(_mux_s_axi_2_r_valid),
		.s_axi_2_r_bits_data(_mux_s_axi_2_r_bits_data),
		.s_axi_3_ar_ready(_mux_s_axi_3_ar_ready),
		.s_axi_3_ar_valid(_vcasRvmRO_3_axi_ar_valid),
		.s_axi_3_ar_bits_addr(_vcasRvmRO_3_axi_ar_bits_addr),
		.s_axi_3_r_ready(_vcasRvmRO_3_axi_r_ready),
		.s_axi_3_r_valid(_mux_s_axi_3_r_valid),
		.s_axi_3_r_bits_data(_mux_s_axi_3_r_bits_data),
		.m_axi_ar_ready(io_internal_vcas_axi_full_0_ar_ready),
		.m_axi_ar_valid(io_internal_vcas_axi_full_0_ar_valid),
		.m_axi_ar_bits_id(_mux_m_axi_ar_bits_id),
		.m_axi_ar_bits_addr(io_internal_vcas_axi_full_0_ar_bits_addr),
		.m_axi_ar_bits_len(io_internal_vcas_axi_full_0_ar_bits_len),
		.m_axi_ar_bits_size(io_internal_vcas_axi_full_0_ar_bits_size),
		.m_axi_ar_bits_burst(io_internal_vcas_axi_full_0_ar_bits_burst),
		.m_axi_ar_bits_lock(io_internal_vcas_axi_full_0_ar_bits_lock),
		.m_axi_ar_bits_cache(io_internal_vcas_axi_full_0_ar_bits_cache),
		.m_axi_ar_bits_prot(io_internal_vcas_axi_full_0_ar_bits_prot),
		.m_axi_ar_bits_qos(io_internal_vcas_axi_full_0_ar_bits_qos),
		.m_axi_ar_bits_region(io_internal_vcas_axi_full_0_ar_bits_region),
		.m_axi_r_ready(io_internal_vcas_axi_full_0_r_ready),
		.m_axi_r_valid(io_internal_vcas_axi_full_0_r_valid),
		.m_axi_r_bits_id(io_internal_vcas_axi_full_0_r_bits_id[2:0]),
		.m_axi_r_bits_data(io_internal_vcas_axi_full_0_r_bits_data),
		.m_axi_r_bits_resp(io_internal_vcas_axi_full_0_r_bits_resp),
		.m_axi_r_bits_last(io_internal_vcas_axi_full_0_r_bits_last),
		.m_axi_aw_ready(io_internal_vcas_axi_full_0_aw_ready),
		.m_axi_aw_valid(io_internal_vcas_axi_full_0_aw_valid),
		.m_axi_aw_bits_id(_mux_m_axi_aw_bits_id),
		.m_axi_aw_bits_addr(io_internal_vcas_axi_full_0_aw_bits_addr),
		.m_axi_aw_bits_len(io_internal_vcas_axi_full_0_aw_bits_len),
		.m_axi_aw_bits_size(io_internal_vcas_axi_full_0_aw_bits_size),
		.m_axi_aw_bits_burst(io_internal_vcas_axi_full_0_aw_bits_burst),
		.m_axi_aw_bits_lock(io_internal_vcas_axi_full_0_aw_bits_lock),
		.m_axi_aw_bits_cache(io_internal_vcas_axi_full_0_aw_bits_cache),
		.m_axi_aw_bits_prot(io_internal_vcas_axi_full_0_aw_bits_prot),
		.m_axi_aw_bits_qos(io_internal_vcas_axi_full_0_aw_bits_qos),
		.m_axi_aw_bits_region(io_internal_vcas_axi_full_0_aw_bits_region),
		.m_axi_w_ready(io_internal_vcas_axi_full_0_w_ready),
		.m_axi_w_valid(io_internal_vcas_axi_full_0_w_valid),
		.m_axi_w_bits_data(io_internal_vcas_axi_full_0_w_bits_data),
		.m_axi_w_bits_strb(io_internal_vcas_axi_full_0_w_bits_strb),
		.m_axi_w_bits_last(io_internal_vcas_axi_full_0_w_bits_last),
		.m_axi_b_ready(io_internal_vcas_axi_full_0_b_ready),
		.m_axi_b_valid(io_internal_vcas_axi_full_0_b_valid),
		.m_axi_b_bits_id(io_internal_vcas_axi_full_0_b_bits_id[2:0]),
		.m_axi_b_bits_resp(io_internal_vcas_axi_full_0_b_bits_resp)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_0(
		.io_dataIn_TREADY(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_0_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_0_bits),
		.io_dataOut_TREADY(io_export_closureOut_0_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_0_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_0_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_1(
		.io_dataIn_TREADY(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_1_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_1_bits),
		.io_dataOut_TREADY(io_export_closureOut_1_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_1_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_1_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_2(
		.io_dataIn_TREADY(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_2_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_2_bits),
		.io_dataOut_TREADY(io_export_closureOut_2_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_2_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_2_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_3(
		.io_dataIn_TREADY(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_3_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_3_bits),
		.io_dataOut_TREADY(io_export_closureOut_3_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_3_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_3_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_4(
		.io_dataIn_TREADY(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_4_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_4_bits),
		.io_dataOut_TREADY(io_export_closureOut_4_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_4_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_4_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_5(
		.io_dataIn_TREADY(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_5_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_5_bits),
		.io_dataOut_TREADY(io_export_closureOut_5_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_5_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_5_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_6(
		.io_dataIn_TREADY(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_6_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_6_bits),
		.io_dataOut_TREADY(io_export_closureOut_6_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_6_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_6_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_7(
		.io_dataIn_TREADY(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_7_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_7_bits),
		.io_dataOut_TREADY(io_export_closureOut_7_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_7_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_7_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_8(
		.io_dataIn_TREADY(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_8_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_8_bits),
		.io_dataOut_TREADY(io_export_closureOut_8_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_8_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_8_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_9(
		.io_dataIn_TREADY(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_9_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_9_bits),
		.io_dataOut_TREADY(io_export_closureOut_9_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_9_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_9_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_10(
		.io_dataIn_TREADY(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_10_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_10_bits),
		.io_dataOut_TREADY(io_export_closureOut_10_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_10_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_10_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_11(
		.io_dataIn_TREADY(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_11_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_11_bits),
		.io_dataOut_TREADY(io_export_closureOut_11_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_11_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_11_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_12(
		.io_dataIn_TREADY(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_12_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_12_bits),
		.io_dataOut_TREADY(io_export_closureOut_12_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_12_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_12_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_13(
		.io_dataIn_TREADY(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_13_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_13_bits),
		.io_dataOut_TREADY(io_export_closureOut_13_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_13_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_13_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_14(
		.io_dataIn_TREADY(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_14_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_14_bits),
		.io_dataOut_TREADY(io_export_closureOut_14_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_14_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_14_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_15(
		.io_dataIn_TREADY(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_15_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_15_bits),
		.io_dataOut_TREADY(io_export_closureOut_15_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_15_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_15_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_16(
		.io_dataIn_TREADY(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_16_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_16_bits),
		.io_dataOut_TREADY(io_export_closureOut_16_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_16_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_16_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_17(
		.io_dataIn_TREADY(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_17_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_17_bits),
		.io_dataOut_TREADY(io_export_closureOut_17_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_17_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_17_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_18(
		.io_dataIn_TREADY(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_18_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_18_bits),
		.io_dataOut_TREADY(io_export_closureOut_18_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_18_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_18_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_19(
		.io_dataIn_TREADY(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_19_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_19_bits),
		.io_dataOut_TREADY(io_export_closureOut_19_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_19_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_19_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_20(
		.io_dataIn_TREADY(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_20_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_20_bits),
		.io_dataOut_TREADY(io_export_closureOut_20_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_20_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_20_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_21(
		.io_dataIn_TREADY(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_21_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_21_bits),
		.io_dataOut_TREADY(io_export_closureOut_21_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_21_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_21_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_22(
		.io_dataIn_TREADY(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_22_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_22_bits),
		.io_dataOut_TREADY(io_export_closureOut_22_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_22_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_22_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_23(
		.io_dataIn_TREADY(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_23_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_23_bits),
		.io_dataOut_TREADY(io_export_closureOut_23_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_23_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_23_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_24(
		.io_dataIn_TREADY(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_24_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_24_bits),
		.io_dataOut_TREADY(io_export_closureOut_24_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_24_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_24_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_25(
		.io_dataIn_TREADY(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_25_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_25_bits),
		.io_dataOut_TREADY(io_export_closureOut_25_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_25_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_25_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_26(
		.io_dataIn_TREADY(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_26_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_26_bits),
		.io_dataOut_TREADY(io_export_closureOut_26_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_26_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_26_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_27(
		.io_dataIn_TREADY(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_27_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_27_bits),
		.io_dataOut_TREADY(io_export_closureOut_27_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_27_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_27_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_28(
		.io_dataIn_TREADY(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_28_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_28_bits),
		.io_dataOut_TREADY(io_export_closureOut_28_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_28_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_28_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_29(
		.io_dataIn_TREADY(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_29_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_29_bits),
		.io_dataOut_TREADY(io_export_closureOut_29_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_29_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_29_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_30(
		.io_dataIn_TREADY(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_30_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_30_bits),
		.io_dataOut_TREADY(io_export_closureOut_30_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_30_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_30_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_31(
		.io_dataIn_TREADY(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_31_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_31_bits),
		.io_dataOut_TREADY(io_export_closureOut_31_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_31_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_31_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_32(
		.io_dataIn_TREADY(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_32_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_32_bits),
		.io_dataOut_TREADY(io_export_closureOut_32_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_32_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_32_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_33(
		.io_dataIn_TREADY(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_33_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_33_bits),
		.io_dataOut_TREADY(io_export_closureOut_33_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_33_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_33_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_34(
		.io_dataIn_TREADY(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_34_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_34_bits),
		.io_dataOut_TREADY(io_export_closureOut_34_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_34_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_34_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_35(
		.io_dataIn_TREADY(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_35_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_35_bits),
		.io_dataOut_TREADY(io_export_closureOut_35_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_35_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_35_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_36(
		.io_dataIn_TREADY(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_36_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_36_bits),
		.io_dataOut_TREADY(io_export_closureOut_36_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_36_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_36_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_37(
		.io_dataIn_TREADY(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_37_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_37_bits),
		.io_dataOut_TREADY(io_export_closureOut_37_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_37_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_37_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_38(
		.io_dataIn_TREADY(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_38_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_38_bits),
		.io_dataOut_TREADY(io_export_closureOut_38_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_38_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_38_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_39(
		.io_dataIn_TREADY(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_39_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_39_bits),
		.io_dataOut_TREADY(io_export_closureOut_39_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_39_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_39_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_40(
		.io_dataIn_TREADY(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_40_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_40_bits),
		.io_dataOut_TREADY(io_export_closureOut_40_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_40_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_40_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_41(
		.io_dataIn_TREADY(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_41_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_41_bits),
		.io_dataOut_TREADY(io_export_closureOut_41_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_41_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_41_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_42(
		.io_dataIn_TREADY(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_42_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_42_bits),
		.io_dataOut_TREADY(io_export_closureOut_42_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_42_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_42_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_43(
		.io_dataIn_TREADY(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_43_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_43_bits),
		.io_dataOut_TREADY(io_export_closureOut_43_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_43_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_43_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_44(
		.io_dataIn_TREADY(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_44_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_44_bits),
		.io_dataOut_TREADY(io_export_closureOut_44_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_44_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_44_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_45(
		.io_dataIn_TREADY(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_45_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_45_bits),
		.io_dataOut_TREADY(io_export_closureOut_45_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_45_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_45_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_46(
		.io_dataIn_TREADY(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_46_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_46_bits),
		.io_dataOut_TREADY(io_export_closureOut_46_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_46_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_46_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_47(
		.io_dataIn_TREADY(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_47_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_47_bits),
		.io_dataOut_TREADY(io_export_closureOut_47_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_47_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_47_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_48(
		.io_dataIn_TREADY(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_48_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_48_bits),
		.io_dataOut_TREADY(io_export_closureOut_48_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_48_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_48_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_49(
		.io_dataIn_TREADY(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_49_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_49_bits),
		.io_dataOut_TREADY(io_export_closureOut_49_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_49_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_49_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_50(
		.io_dataIn_TREADY(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_50_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_50_bits),
		.io_dataOut_TREADY(io_export_closureOut_50_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_50_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_50_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_51(
		.io_dataIn_TREADY(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_51_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_51_bits),
		.io_dataOut_TREADY(io_export_closureOut_51_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_51_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_51_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_52(
		.io_dataIn_TREADY(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_52_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_52_bits),
		.io_dataOut_TREADY(io_export_closureOut_52_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_52_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_52_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_53(
		.io_dataIn_TREADY(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_53_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_53_bits),
		.io_dataOut_TREADY(io_export_closureOut_53_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_53_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_53_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_54(
		.io_dataIn_TREADY(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_54_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_54_bits),
		.io_dataOut_TREADY(io_export_closureOut_54_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_54_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_54_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_55(
		.io_dataIn_TREADY(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_55_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_55_bits),
		.io_dataOut_TREADY(io_export_closureOut_55_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_55_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_55_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_56(
		.io_dataIn_TREADY(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_56_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_56_bits),
		.io_dataOut_TREADY(io_export_closureOut_56_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_56_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_56_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_57(
		.io_dataIn_TREADY(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_57_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_57_bits),
		.io_dataOut_TREADY(io_export_closureOut_57_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_57_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_57_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_58(
		.io_dataIn_TREADY(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_58_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_58_bits),
		.io_dataOut_TREADY(io_export_closureOut_58_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_58_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_58_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_59(
		.io_dataIn_TREADY(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_59_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_59_bits),
		.io_dataOut_TREADY(io_export_closureOut_59_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_59_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_59_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_60(
		.io_dataIn_TREADY(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_60_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_60_bits),
		.io_dataOut_TREADY(io_export_closureOut_60_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_60_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_60_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_61(
		.io_dataIn_TREADY(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_61_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_61_bits),
		.io_dataOut_TREADY(io_export_closureOut_61_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_61_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_61_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_62(
		.io_dataIn_TREADY(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_62_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_62_bits),
		.io_dataOut_TREADY(io_export_closureOut_62_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_62_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_62_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_out_63(
		.io_dataIn_TREADY(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_63_valid),
		.io_dataIn_TDATA(_continuationNetwork_io_connPE_63_bits),
		.io_dataOut_TREADY(io_export_closureOut_63_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_63_TVALID),
		.io_dataOut_TDATA(io_export_closureOut_63_TDATA)
	);
	assign io_internal_vcas_axi_full_0_ar_bits_id = {4'h0, _mux_m_axi_ar_bits_id};
	assign io_internal_vcas_axi_full_0_aw_bits_id = {4'h0, _mux_m_axi_aw_bits_id};
endmodule
module ArgumentNotifierNetworkUnit (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_peAddress_ready,
	io_peAddress_valid,
	io_peAddress_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	output wire io_peAddress_ready;
	input io_peAddress_valid;
	input [63:0] io_peAddress_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg stateReg;
	reg [63:0] addressReg;
	reg priorityReg;
	wire _GEN = io_addressIn_valid & io_peAddress_valid;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 1'h0;
			addressReg <= 64'h0000000000000000;
			priorityReg <= 1'h1;
		end
		else begin
			if (stateReg)
				stateReg <= stateReg & ~io_addressOut_ready;
			else begin
				stateReg <= (io_addressIn_valid | io_peAddress_valid) | stateReg;
				if (_GEN)
					addressReg <= (priorityReg ? io_peAddress_bits : io_addressIn_bits);
				else if (io_peAddress_valid)
					addressReg <= io_peAddress_bits;
				else if (io_addressIn_valid)
					addressReg <= io_addressIn_bits;
			end
			priorityReg <= (~stateReg & _GEN) ^ priorityReg;
		end
	assign io_addressIn_ready = ~stateReg & (_GEN ? ~priorityReg : ~io_peAddress_valid & io_addressIn_valid);
	assign io_peAddress_ready = ~stateReg & (_GEN ? priorityReg : io_peAddress_valid);
	assign io_addressOut_valid = stateReg;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h0 ? 2'h2 : 2'h1);
			end
			else if (_GEN_0 | ~(_GEN_1 & io_vasAddressOut_ready))
				;
			else
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_1 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h1 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_2 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h2 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_3 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h3 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_4 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h4 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_5 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h5 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_6 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h6 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_7 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h7 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_8 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h8 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_9 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'h9 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_10 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'ha ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_11 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'hb ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_12 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'hc ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_13 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'hd ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_14 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[8:5] == 4'he ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_15 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (&io_addressIn_bits[8:5] ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ram_32x64 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [4:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [63:0] R0_data;
	input [4:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [63:0] W0_data;
	reg [63:0] Memory [0:31];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue32_UInt (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits;
	reg [4:0] enq_ptr_value;
	reg [4:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 5'h00;
			deq_ptr_value <= 5'h00;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 5'h01;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 5'h01;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_32x64 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module AllocatorBuffer_64 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	Queue32_UInt q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_addressIn_ready),
		.io_enq_valid(io_addressIn_valid),
		.io_enq_bits(io_addressIn_bits),
		.io_deq_ready(io_addressOut_ready),
		.io_deq_valid(io_addressOut_valid),
		.io_deq_bits(io_addressOut_bits)
	);
endmodule
module ArgumentNotifierNetwork (
	clock,
	reset,
	io_connVAS_0_ready,
	io_connVAS_0_valid,
	io_connVAS_0_bits,
	io_connVAS_1_ready,
	io_connVAS_1_valid,
	io_connVAS_1_bits,
	io_connVAS_2_ready,
	io_connVAS_2_valid,
	io_connVAS_2_bits,
	io_connVAS_3_ready,
	io_connVAS_3_valid,
	io_connVAS_3_bits,
	io_connVAS_4_ready,
	io_connVAS_4_valid,
	io_connVAS_4_bits,
	io_connVAS_5_ready,
	io_connVAS_5_valid,
	io_connVAS_5_bits,
	io_connVAS_6_ready,
	io_connVAS_6_valid,
	io_connVAS_6_bits,
	io_connVAS_7_ready,
	io_connVAS_7_valid,
	io_connVAS_7_bits,
	io_connVAS_8_ready,
	io_connVAS_8_valid,
	io_connVAS_8_bits,
	io_connVAS_9_ready,
	io_connVAS_9_valid,
	io_connVAS_9_bits,
	io_connVAS_10_ready,
	io_connVAS_10_valid,
	io_connVAS_10_bits,
	io_connVAS_11_ready,
	io_connVAS_11_valid,
	io_connVAS_11_bits,
	io_connVAS_12_ready,
	io_connVAS_12_valid,
	io_connVAS_12_bits,
	io_connVAS_13_ready,
	io_connVAS_13_valid,
	io_connVAS_13_bits,
	io_connVAS_14_ready,
	io_connVAS_14_valid,
	io_connVAS_14_bits,
	io_connVAS_15_ready,
	io_connVAS_15_valid,
	io_connVAS_15_bits,
	io_connPE_0_ready,
	io_connPE_0_valid,
	io_connPE_0_bits,
	io_connPE_1_ready,
	io_connPE_1_valid,
	io_connPE_1_bits,
	io_connPE_2_ready,
	io_connPE_2_valid,
	io_connPE_2_bits,
	io_connPE_3_ready,
	io_connPE_3_valid,
	io_connPE_3_bits,
	io_connPE_4_ready,
	io_connPE_4_valid,
	io_connPE_4_bits,
	io_connPE_5_ready,
	io_connPE_5_valid,
	io_connPE_5_bits,
	io_connPE_6_ready,
	io_connPE_6_valid,
	io_connPE_6_bits,
	io_connPE_7_ready,
	io_connPE_7_valid,
	io_connPE_7_bits,
	io_connPE_8_ready,
	io_connPE_8_valid,
	io_connPE_8_bits,
	io_connPE_9_ready,
	io_connPE_9_valid,
	io_connPE_9_bits,
	io_connPE_10_ready,
	io_connPE_10_valid,
	io_connPE_10_bits,
	io_connPE_11_ready,
	io_connPE_11_valid,
	io_connPE_11_bits,
	io_connPE_12_ready,
	io_connPE_12_valid,
	io_connPE_12_bits,
	io_connPE_13_ready,
	io_connPE_13_valid,
	io_connPE_13_bits,
	io_connPE_14_ready,
	io_connPE_14_valid,
	io_connPE_14_bits,
	io_connPE_15_ready,
	io_connPE_15_valid,
	io_connPE_15_bits,
	io_connPE_16_ready,
	io_connPE_16_valid,
	io_connPE_16_bits,
	io_connPE_17_ready,
	io_connPE_17_valid,
	io_connPE_17_bits,
	io_connPE_18_ready,
	io_connPE_18_valid,
	io_connPE_18_bits,
	io_connPE_19_ready,
	io_connPE_19_valid,
	io_connPE_19_bits,
	io_connPE_20_ready,
	io_connPE_20_valid,
	io_connPE_20_bits,
	io_connPE_21_ready,
	io_connPE_21_valid,
	io_connPE_21_bits,
	io_connPE_22_ready,
	io_connPE_22_valid,
	io_connPE_22_bits,
	io_connPE_23_ready,
	io_connPE_23_valid,
	io_connPE_23_bits,
	io_connPE_24_ready,
	io_connPE_24_valid,
	io_connPE_24_bits,
	io_connPE_25_ready,
	io_connPE_25_valid,
	io_connPE_25_bits,
	io_connPE_26_ready,
	io_connPE_26_valid,
	io_connPE_26_bits,
	io_connPE_27_ready,
	io_connPE_27_valid,
	io_connPE_27_bits,
	io_connPE_28_ready,
	io_connPE_28_valid,
	io_connPE_28_bits,
	io_connPE_29_ready,
	io_connPE_29_valid,
	io_connPE_29_bits,
	io_connPE_30_ready,
	io_connPE_30_valid,
	io_connPE_30_bits,
	io_connPE_31_ready,
	io_connPE_31_valid,
	io_connPE_31_bits,
	io_connPE_32_ready,
	io_connPE_32_valid,
	io_connPE_32_bits,
	io_connPE_33_ready,
	io_connPE_33_valid,
	io_connPE_33_bits,
	io_connPE_34_ready,
	io_connPE_34_valid,
	io_connPE_34_bits,
	io_connPE_35_ready,
	io_connPE_35_valid,
	io_connPE_35_bits,
	io_connPE_36_ready,
	io_connPE_36_valid,
	io_connPE_36_bits,
	io_connPE_37_ready,
	io_connPE_37_valid,
	io_connPE_37_bits,
	io_connPE_38_ready,
	io_connPE_38_valid,
	io_connPE_38_bits,
	io_connPE_39_ready,
	io_connPE_39_valid,
	io_connPE_39_bits,
	io_connPE_40_ready,
	io_connPE_40_valid,
	io_connPE_40_bits,
	io_connPE_41_ready,
	io_connPE_41_valid,
	io_connPE_41_bits,
	io_connPE_42_ready,
	io_connPE_42_valid,
	io_connPE_42_bits,
	io_connPE_43_ready,
	io_connPE_43_valid,
	io_connPE_43_bits,
	io_connPE_44_ready,
	io_connPE_44_valid,
	io_connPE_44_bits,
	io_connPE_45_ready,
	io_connPE_45_valid,
	io_connPE_45_bits,
	io_connPE_46_ready,
	io_connPE_46_valid,
	io_connPE_46_bits,
	io_connPE_47_ready,
	io_connPE_47_valid,
	io_connPE_47_bits,
	io_connPE_48_ready,
	io_connPE_48_valid,
	io_connPE_48_bits,
	io_connPE_49_ready,
	io_connPE_49_valid,
	io_connPE_49_bits,
	io_connPE_50_ready,
	io_connPE_50_valid,
	io_connPE_50_bits,
	io_connPE_51_ready,
	io_connPE_51_valid,
	io_connPE_51_bits,
	io_connPE_52_ready,
	io_connPE_52_valid,
	io_connPE_52_bits,
	io_connPE_53_ready,
	io_connPE_53_valid,
	io_connPE_53_bits,
	io_connPE_54_ready,
	io_connPE_54_valid,
	io_connPE_54_bits,
	io_connPE_55_ready,
	io_connPE_55_valid,
	io_connPE_55_bits,
	io_connPE_56_ready,
	io_connPE_56_valid,
	io_connPE_56_bits,
	io_connPE_57_ready,
	io_connPE_57_valid,
	io_connPE_57_bits,
	io_connPE_58_ready,
	io_connPE_58_valid,
	io_connPE_58_bits,
	io_connPE_59_ready,
	io_connPE_59_valid,
	io_connPE_59_bits,
	io_connPE_60_ready,
	io_connPE_60_valid,
	io_connPE_60_bits,
	io_connPE_61_ready,
	io_connPE_61_valid,
	io_connPE_61_bits,
	io_connPE_62_ready,
	io_connPE_62_valid,
	io_connPE_62_bits,
	io_connPE_63_ready,
	io_connPE_63_valid,
	io_connPE_63_bits,
	io_connPE_64_ready,
	io_connPE_64_valid,
	io_connPE_64_bits,
	io_connPE_65_ready,
	io_connPE_65_valid,
	io_connPE_65_bits,
	io_connPE_66_ready,
	io_connPE_66_valid,
	io_connPE_66_bits,
	io_connPE_67_ready,
	io_connPE_67_valid,
	io_connPE_67_bits,
	io_connPE_68_ready,
	io_connPE_68_valid,
	io_connPE_68_bits,
	io_connPE_69_ready,
	io_connPE_69_valid,
	io_connPE_69_bits,
	io_connPE_70_ready,
	io_connPE_70_valid,
	io_connPE_70_bits,
	io_connPE_71_ready,
	io_connPE_71_valid,
	io_connPE_71_bits,
	io_connPE_72_ready,
	io_connPE_72_valid,
	io_connPE_72_bits,
	io_connPE_73_ready,
	io_connPE_73_valid,
	io_connPE_73_bits,
	io_connPE_74_ready,
	io_connPE_74_valid,
	io_connPE_74_bits,
	io_connPE_75_ready,
	io_connPE_75_valid,
	io_connPE_75_bits,
	io_connPE_76_ready,
	io_connPE_76_valid,
	io_connPE_76_bits,
	io_connPE_77_ready,
	io_connPE_77_valid,
	io_connPE_77_bits,
	io_connPE_78_ready,
	io_connPE_78_valid,
	io_connPE_78_bits,
	io_connPE_79_ready,
	io_connPE_79_valid,
	io_connPE_79_bits,
	io_connPE_80_ready,
	io_connPE_80_valid,
	io_connPE_80_bits,
	io_connPE_81_ready,
	io_connPE_81_valid,
	io_connPE_81_bits,
	io_connPE_82_ready,
	io_connPE_82_valid,
	io_connPE_82_bits,
	io_connPE_83_ready,
	io_connPE_83_valid,
	io_connPE_83_bits,
	io_connPE_84_ready,
	io_connPE_84_valid,
	io_connPE_84_bits,
	io_connPE_85_ready,
	io_connPE_85_valid,
	io_connPE_85_bits,
	io_connPE_86_ready,
	io_connPE_86_valid,
	io_connPE_86_bits,
	io_connPE_87_ready,
	io_connPE_87_valid,
	io_connPE_87_bits,
	io_connPE_88_ready,
	io_connPE_88_valid,
	io_connPE_88_bits,
	io_connPE_89_ready,
	io_connPE_89_valid,
	io_connPE_89_bits,
	io_connPE_90_ready,
	io_connPE_90_valid,
	io_connPE_90_bits,
	io_connPE_91_ready,
	io_connPE_91_valid,
	io_connPE_91_bits,
	io_connPE_92_ready,
	io_connPE_92_valid,
	io_connPE_92_bits,
	io_connPE_93_ready,
	io_connPE_93_valid,
	io_connPE_93_bits,
	io_connPE_94_ready,
	io_connPE_94_valid,
	io_connPE_94_bits,
	io_connPE_95_ready,
	io_connPE_95_valid,
	io_connPE_95_bits,
	io_connPE_96_ready,
	io_connPE_96_valid,
	io_connPE_96_bits,
	io_connPE_97_ready,
	io_connPE_97_valid,
	io_connPE_97_bits,
	io_connPE_98_ready,
	io_connPE_98_valid,
	io_connPE_98_bits,
	io_connPE_99_ready,
	io_connPE_99_valid,
	io_connPE_99_bits,
	io_connPE_100_ready,
	io_connPE_100_valid,
	io_connPE_100_bits,
	io_connPE_101_ready,
	io_connPE_101_valid,
	io_connPE_101_bits,
	io_connPE_102_ready,
	io_connPE_102_valid,
	io_connPE_102_bits,
	io_connPE_103_ready,
	io_connPE_103_valid,
	io_connPE_103_bits,
	io_connPE_104_ready,
	io_connPE_104_valid,
	io_connPE_104_bits,
	io_connPE_105_ready,
	io_connPE_105_valid,
	io_connPE_105_bits,
	io_connPE_106_ready,
	io_connPE_106_valid,
	io_connPE_106_bits,
	io_connPE_107_ready,
	io_connPE_107_valid,
	io_connPE_107_bits,
	io_connPE_108_ready,
	io_connPE_108_valid,
	io_connPE_108_bits,
	io_connPE_109_ready,
	io_connPE_109_valid,
	io_connPE_109_bits,
	io_connPE_110_ready,
	io_connPE_110_valid,
	io_connPE_110_bits,
	io_connPE_111_ready,
	io_connPE_111_valid,
	io_connPE_111_bits,
	io_connPE_112_ready,
	io_connPE_112_valid,
	io_connPE_112_bits,
	io_connPE_113_ready,
	io_connPE_113_valid,
	io_connPE_113_bits,
	io_connPE_114_ready,
	io_connPE_114_valid,
	io_connPE_114_bits,
	io_connPE_115_ready,
	io_connPE_115_valid,
	io_connPE_115_bits,
	io_connPE_116_ready,
	io_connPE_116_valid,
	io_connPE_116_bits,
	io_connPE_117_ready,
	io_connPE_117_valid,
	io_connPE_117_bits,
	io_connPE_118_ready,
	io_connPE_118_valid,
	io_connPE_118_bits,
	io_connPE_119_ready,
	io_connPE_119_valid,
	io_connPE_119_bits,
	io_connPE_120_ready,
	io_connPE_120_valid,
	io_connPE_120_bits,
	io_connPE_121_ready,
	io_connPE_121_valid,
	io_connPE_121_bits,
	io_connPE_122_ready,
	io_connPE_122_valid,
	io_connPE_122_bits,
	io_connPE_123_ready,
	io_connPE_123_valid,
	io_connPE_123_bits,
	io_connPE_124_ready,
	io_connPE_124_valid,
	io_connPE_124_bits,
	io_connPE_125_ready,
	io_connPE_125_valid,
	io_connPE_125_bits,
	io_connPE_126_ready,
	io_connPE_126_valid,
	io_connPE_126_bits,
	io_connPE_127_ready,
	io_connPE_127_valid,
	io_connPE_127_bits
);
	input clock;
	input reset;
	input io_connVAS_0_ready;
	output wire io_connVAS_0_valid;
	output wire [63:0] io_connVAS_0_bits;
	input io_connVAS_1_ready;
	output wire io_connVAS_1_valid;
	output wire [63:0] io_connVAS_1_bits;
	input io_connVAS_2_ready;
	output wire io_connVAS_2_valid;
	output wire [63:0] io_connVAS_2_bits;
	input io_connVAS_3_ready;
	output wire io_connVAS_3_valid;
	output wire [63:0] io_connVAS_3_bits;
	input io_connVAS_4_ready;
	output wire io_connVAS_4_valid;
	output wire [63:0] io_connVAS_4_bits;
	input io_connVAS_5_ready;
	output wire io_connVAS_5_valid;
	output wire [63:0] io_connVAS_5_bits;
	input io_connVAS_6_ready;
	output wire io_connVAS_6_valid;
	output wire [63:0] io_connVAS_6_bits;
	input io_connVAS_7_ready;
	output wire io_connVAS_7_valid;
	output wire [63:0] io_connVAS_7_bits;
	input io_connVAS_8_ready;
	output wire io_connVAS_8_valid;
	output wire [63:0] io_connVAS_8_bits;
	input io_connVAS_9_ready;
	output wire io_connVAS_9_valid;
	output wire [63:0] io_connVAS_9_bits;
	input io_connVAS_10_ready;
	output wire io_connVAS_10_valid;
	output wire [63:0] io_connVAS_10_bits;
	input io_connVAS_11_ready;
	output wire io_connVAS_11_valid;
	output wire [63:0] io_connVAS_11_bits;
	input io_connVAS_12_ready;
	output wire io_connVAS_12_valid;
	output wire [63:0] io_connVAS_12_bits;
	input io_connVAS_13_ready;
	output wire io_connVAS_13_valid;
	output wire [63:0] io_connVAS_13_bits;
	input io_connVAS_14_ready;
	output wire io_connVAS_14_valid;
	output wire [63:0] io_connVAS_14_bits;
	input io_connVAS_15_ready;
	output wire io_connVAS_15_valid;
	output wire [63:0] io_connVAS_15_bits;
	output wire io_connPE_0_ready;
	input io_connPE_0_valid;
	input [63:0] io_connPE_0_bits;
	output wire io_connPE_1_ready;
	input io_connPE_1_valid;
	input [63:0] io_connPE_1_bits;
	output wire io_connPE_2_ready;
	input io_connPE_2_valid;
	input [63:0] io_connPE_2_bits;
	output wire io_connPE_3_ready;
	input io_connPE_3_valid;
	input [63:0] io_connPE_3_bits;
	output wire io_connPE_4_ready;
	input io_connPE_4_valid;
	input [63:0] io_connPE_4_bits;
	output wire io_connPE_5_ready;
	input io_connPE_5_valid;
	input [63:0] io_connPE_5_bits;
	output wire io_connPE_6_ready;
	input io_connPE_6_valid;
	input [63:0] io_connPE_6_bits;
	output wire io_connPE_7_ready;
	input io_connPE_7_valid;
	input [63:0] io_connPE_7_bits;
	output wire io_connPE_8_ready;
	input io_connPE_8_valid;
	input [63:0] io_connPE_8_bits;
	output wire io_connPE_9_ready;
	input io_connPE_9_valid;
	input [63:0] io_connPE_9_bits;
	output wire io_connPE_10_ready;
	input io_connPE_10_valid;
	input [63:0] io_connPE_10_bits;
	output wire io_connPE_11_ready;
	input io_connPE_11_valid;
	input [63:0] io_connPE_11_bits;
	output wire io_connPE_12_ready;
	input io_connPE_12_valid;
	input [63:0] io_connPE_12_bits;
	output wire io_connPE_13_ready;
	input io_connPE_13_valid;
	input [63:0] io_connPE_13_bits;
	output wire io_connPE_14_ready;
	input io_connPE_14_valid;
	input [63:0] io_connPE_14_bits;
	output wire io_connPE_15_ready;
	input io_connPE_15_valid;
	input [63:0] io_connPE_15_bits;
	output wire io_connPE_16_ready;
	input io_connPE_16_valid;
	input [63:0] io_connPE_16_bits;
	output wire io_connPE_17_ready;
	input io_connPE_17_valid;
	input [63:0] io_connPE_17_bits;
	output wire io_connPE_18_ready;
	input io_connPE_18_valid;
	input [63:0] io_connPE_18_bits;
	output wire io_connPE_19_ready;
	input io_connPE_19_valid;
	input [63:0] io_connPE_19_bits;
	output wire io_connPE_20_ready;
	input io_connPE_20_valid;
	input [63:0] io_connPE_20_bits;
	output wire io_connPE_21_ready;
	input io_connPE_21_valid;
	input [63:0] io_connPE_21_bits;
	output wire io_connPE_22_ready;
	input io_connPE_22_valid;
	input [63:0] io_connPE_22_bits;
	output wire io_connPE_23_ready;
	input io_connPE_23_valid;
	input [63:0] io_connPE_23_bits;
	output wire io_connPE_24_ready;
	input io_connPE_24_valid;
	input [63:0] io_connPE_24_bits;
	output wire io_connPE_25_ready;
	input io_connPE_25_valid;
	input [63:0] io_connPE_25_bits;
	output wire io_connPE_26_ready;
	input io_connPE_26_valid;
	input [63:0] io_connPE_26_bits;
	output wire io_connPE_27_ready;
	input io_connPE_27_valid;
	input [63:0] io_connPE_27_bits;
	output wire io_connPE_28_ready;
	input io_connPE_28_valid;
	input [63:0] io_connPE_28_bits;
	output wire io_connPE_29_ready;
	input io_connPE_29_valid;
	input [63:0] io_connPE_29_bits;
	output wire io_connPE_30_ready;
	input io_connPE_30_valid;
	input [63:0] io_connPE_30_bits;
	output wire io_connPE_31_ready;
	input io_connPE_31_valid;
	input [63:0] io_connPE_31_bits;
	output wire io_connPE_32_ready;
	input io_connPE_32_valid;
	input [63:0] io_connPE_32_bits;
	output wire io_connPE_33_ready;
	input io_connPE_33_valid;
	input [63:0] io_connPE_33_bits;
	output wire io_connPE_34_ready;
	input io_connPE_34_valid;
	input [63:0] io_connPE_34_bits;
	output wire io_connPE_35_ready;
	input io_connPE_35_valid;
	input [63:0] io_connPE_35_bits;
	output wire io_connPE_36_ready;
	input io_connPE_36_valid;
	input [63:0] io_connPE_36_bits;
	output wire io_connPE_37_ready;
	input io_connPE_37_valid;
	input [63:0] io_connPE_37_bits;
	output wire io_connPE_38_ready;
	input io_connPE_38_valid;
	input [63:0] io_connPE_38_bits;
	output wire io_connPE_39_ready;
	input io_connPE_39_valid;
	input [63:0] io_connPE_39_bits;
	output wire io_connPE_40_ready;
	input io_connPE_40_valid;
	input [63:0] io_connPE_40_bits;
	output wire io_connPE_41_ready;
	input io_connPE_41_valid;
	input [63:0] io_connPE_41_bits;
	output wire io_connPE_42_ready;
	input io_connPE_42_valid;
	input [63:0] io_connPE_42_bits;
	output wire io_connPE_43_ready;
	input io_connPE_43_valid;
	input [63:0] io_connPE_43_bits;
	output wire io_connPE_44_ready;
	input io_connPE_44_valid;
	input [63:0] io_connPE_44_bits;
	output wire io_connPE_45_ready;
	input io_connPE_45_valid;
	input [63:0] io_connPE_45_bits;
	output wire io_connPE_46_ready;
	input io_connPE_46_valid;
	input [63:0] io_connPE_46_bits;
	output wire io_connPE_47_ready;
	input io_connPE_47_valid;
	input [63:0] io_connPE_47_bits;
	output wire io_connPE_48_ready;
	input io_connPE_48_valid;
	input [63:0] io_connPE_48_bits;
	output wire io_connPE_49_ready;
	input io_connPE_49_valid;
	input [63:0] io_connPE_49_bits;
	output wire io_connPE_50_ready;
	input io_connPE_50_valid;
	input [63:0] io_connPE_50_bits;
	output wire io_connPE_51_ready;
	input io_connPE_51_valid;
	input [63:0] io_connPE_51_bits;
	output wire io_connPE_52_ready;
	input io_connPE_52_valid;
	input [63:0] io_connPE_52_bits;
	output wire io_connPE_53_ready;
	input io_connPE_53_valid;
	input [63:0] io_connPE_53_bits;
	output wire io_connPE_54_ready;
	input io_connPE_54_valid;
	input [63:0] io_connPE_54_bits;
	output wire io_connPE_55_ready;
	input io_connPE_55_valid;
	input [63:0] io_connPE_55_bits;
	output wire io_connPE_56_ready;
	input io_connPE_56_valid;
	input [63:0] io_connPE_56_bits;
	output wire io_connPE_57_ready;
	input io_connPE_57_valid;
	input [63:0] io_connPE_57_bits;
	output wire io_connPE_58_ready;
	input io_connPE_58_valid;
	input [63:0] io_connPE_58_bits;
	output wire io_connPE_59_ready;
	input io_connPE_59_valid;
	input [63:0] io_connPE_59_bits;
	output wire io_connPE_60_ready;
	input io_connPE_60_valid;
	input [63:0] io_connPE_60_bits;
	output wire io_connPE_61_ready;
	input io_connPE_61_valid;
	input [63:0] io_connPE_61_bits;
	output wire io_connPE_62_ready;
	input io_connPE_62_valid;
	input [63:0] io_connPE_62_bits;
	output wire io_connPE_63_ready;
	input io_connPE_63_valid;
	input [63:0] io_connPE_63_bits;
	output wire io_connPE_64_ready;
	input io_connPE_64_valid;
	input [63:0] io_connPE_64_bits;
	output wire io_connPE_65_ready;
	input io_connPE_65_valid;
	input [63:0] io_connPE_65_bits;
	output wire io_connPE_66_ready;
	input io_connPE_66_valid;
	input [63:0] io_connPE_66_bits;
	output wire io_connPE_67_ready;
	input io_connPE_67_valid;
	input [63:0] io_connPE_67_bits;
	output wire io_connPE_68_ready;
	input io_connPE_68_valid;
	input [63:0] io_connPE_68_bits;
	output wire io_connPE_69_ready;
	input io_connPE_69_valid;
	input [63:0] io_connPE_69_bits;
	output wire io_connPE_70_ready;
	input io_connPE_70_valid;
	input [63:0] io_connPE_70_bits;
	output wire io_connPE_71_ready;
	input io_connPE_71_valid;
	input [63:0] io_connPE_71_bits;
	output wire io_connPE_72_ready;
	input io_connPE_72_valid;
	input [63:0] io_connPE_72_bits;
	output wire io_connPE_73_ready;
	input io_connPE_73_valid;
	input [63:0] io_connPE_73_bits;
	output wire io_connPE_74_ready;
	input io_connPE_74_valid;
	input [63:0] io_connPE_74_bits;
	output wire io_connPE_75_ready;
	input io_connPE_75_valid;
	input [63:0] io_connPE_75_bits;
	output wire io_connPE_76_ready;
	input io_connPE_76_valid;
	input [63:0] io_connPE_76_bits;
	output wire io_connPE_77_ready;
	input io_connPE_77_valid;
	input [63:0] io_connPE_77_bits;
	output wire io_connPE_78_ready;
	input io_connPE_78_valid;
	input [63:0] io_connPE_78_bits;
	output wire io_connPE_79_ready;
	input io_connPE_79_valid;
	input [63:0] io_connPE_79_bits;
	output wire io_connPE_80_ready;
	input io_connPE_80_valid;
	input [63:0] io_connPE_80_bits;
	output wire io_connPE_81_ready;
	input io_connPE_81_valid;
	input [63:0] io_connPE_81_bits;
	output wire io_connPE_82_ready;
	input io_connPE_82_valid;
	input [63:0] io_connPE_82_bits;
	output wire io_connPE_83_ready;
	input io_connPE_83_valid;
	input [63:0] io_connPE_83_bits;
	output wire io_connPE_84_ready;
	input io_connPE_84_valid;
	input [63:0] io_connPE_84_bits;
	output wire io_connPE_85_ready;
	input io_connPE_85_valid;
	input [63:0] io_connPE_85_bits;
	output wire io_connPE_86_ready;
	input io_connPE_86_valid;
	input [63:0] io_connPE_86_bits;
	output wire io_connPE_87_ready;
	input io_connPE_87_valid;
	input [63:0] io_connPE_87_bits;
	output wire io_connPE_88_ready;
	input io_connPE_88_valid;
	input [63:0] io_connPE_88_bits;
	output wire io_connPE_89_ready;
	input io_connPE_89_valid;
	input [63:0] io_connPE_89_bits;
	output wire io_connPE_90_ready;
	input io_connPE_90_valid;
	input [63:0] io_connPE_90_bits;
	output wire io_connPE_91_ready;
	input io_connPE_91_valid;
	input [63:0] io_connPE_91_bits;
	output wire io_connPE_92_ready;
	input io_connPE_92_valid;
	input [63:0] io_connPE_92_bits;
	output wire io_connPE_93_ready;
	input io_connPE_93_valid;
	input [63:0] io_connPE_93_bits;
	output wire io_connPE_94_ready;
	input io_connPE_94_valid;
	input [63:0] io_connPE_94_bits;
	output wire io_connPE_95_ready;
	input io_connPE_95_valid;
	input [63:0] io_connPE_95_bits;
	output wire io_connPE_96_ready;
	input io_connPE_96_valid;
	input [63:0] io_connPE_96_bits;
	output wire io_connPE_97_ready;
	input io_connPE_97_valid;
	input [63:0] io_connPE_97_bits;
	output wire io_connPE_98_ready;
	input io_connPE_98_valid;
	input [63:0] io_connPE_98_bits;
	output wire io_connPE_99_ready;
	input io_connPE_99_valid;
	input [63:0] io_connPE_99_bits;
	output wire io_connPE_100_ready;
	input io_connPE_100_valid;
	input [63:0] io_connPE_100_bits;
	output wire io_connPE_101_ready;
	input io_connPE_101_valid;
	input [63:0] io_connPE_101_bits;
	output wire io_connPE_102_ready;
	input io_connPE_102_valid;
	input [63:0] io_connPE_102_bits;
	output wire io_connPE_103_ready;
	input io_connPE_103_valid;
	input [63:0] io_connPE_103_bits;
	output wire io_connPE_104_ready;
	input io_connPE_104_valid;
	input [63:0] io_connPE_104_bits;
	output wire io_connPE_105_ready;
	input io_connPE_105_valid;
	input [63:0] io_connPE_105_bits;
	output wire io_connPE_106_ready;
	input io_connPE_106_valid;
	input [63:0] io_connPE_106_bits;
	output wire io_connPE_107_ready;
	input io_connPE_107_valid;
	input [63:0] io_connPE_107_bits;
	output wire io_connPE_108_ready;
	input io_connPE_108_valid;
	input [63:0] io_connPE_108_bits;
	output wire io_connPE_109_ready;
	input io_connPE_109_valid;
	input [63:0] io_connPE_109_bits;
	output wire io_connPE_110_ready;
	input io_connPE_110_valid;
	input [63:0] io_connPE_110_bits;
	output wire io_connPE_111_ready;
	input io_connPE_111_valid;
	input [63:0] io_connPE_111_bits;
	output wire io_connPE_112_ready;
	input io_connPE_112_valid;
	input [63:0] io_connPE_112_bits;
	output wire io_connPE_113_ready;
	input io_connPE_113_valid;
	input [63:0] io_connPE_113_bits;
	output wire io_connPE_114_ready;
	input io_connPE_114_valid;
	input [63:0] io_connPE_114_bits;
	output wire io_connPE_115_ready;
	input io_connPE_115_valid;
	input [63:0] io_connPE_115_bits;
	output wire io_connPE_116_ready;
	input io_connPE_116_valid;
	input [63:0] io_connPE_116_bits;
	output wire io_connPE_117_ready;
	input io_connPE_117_valid;
	input [63:0] io_connPE_117_bits;
	output wire io_connPE_118_ready;
	input io_connPE_118_valid;
	input [63:0] io_connPE_118_bits;
	output wire io_connPE_119_ready;
	input io_connPE_119_valid;
	input [63:0] io_connPE_119_bits;
	output wire io_connPE_120_ready;
	input io_connPE_120_valid;
	input [63:0] io_connPE_120_bits;
	output wire io_connPE_121_ready;
	input io_connPE_121_valid;
	input [63:0] io_connPE_121_bits;
	output wire io_connPE_122_ready;
	input io_connPE_122_valid;
	input [63:0] io_connPE_122_bits;
	output wire io_connPE_123_ready;
	input io_connPE_123_valid;
	input [63:0] io_connPE_123_bits;
	output wire io_connPE_124_ready;
	input io_connPE_124_valid;
	input [63:0] io_connPE_124_bits;
	output wire io_connPE_125_ready;
	input io_connPE_125_valid;
	input [63:0] io_connPE_125_bits;
	output wire io_connPE_126_ready;
	input io_connPE_126_valid;
	input [63:0] io_connPE_126_bits;
	output wire io_connPE_127_ready;
	input io_connPE_127_valid;
	input [63:0] io_connPE_127_bits;
	wire _queues_127_io_addressOut_valid;
	wire [63:0] _queues_127_io_addressOut_bits;
	wire _queues_126_io_addressOut_valid;
	wire [63:0] _queues_126_io_addressOut_bits;
	wire _queues_125_io_addressOut_valid;
	wire [63:0] _queues_125_io_addressOut_bits;
	wire _queues_124_io_addressOut_valid;
	wire [63:0] _queues_124_io_addressOut_bits;
	wire _queues_123_io_addressOut_valid;
	wire [63:0] _queues_123_io_addressOut_bits;
	wire _queues_122_io_addressOut_valid;
	wire [63:0] _queues_122_io_addressOut_bits;
	wire _queues_121_io_addressOut_valid;
	wire [63:0] _queues_121_io_addressOut_bits;
	wire _queues_120_io_addressOut_valid;
	wire [63:0] _queues_120_io_addressOut_bits;
	wire _queues_119_io_addressOut_valid;
	wire [63:0] _queues_119_io_addressOut_bits;
	wire _queues_118_io_addressOut_valid;
	wire [63:0] _queues_118_io_addressOut_bits;
	wire _queues_117_io_addressOut_valid;
	wire [63:0] _queues_117_io_addressOut_bits;
	wire _queues_116_io_addressOut_valid;
	wire [63:0] _queues_116_io_addressOut_bits;
	wire _queues_115_io_addressOut_valid;
	wire [63:0] _queues_115_io_addressOut_bits;
	wire _queues_114_io_addressOut_valid;
	wire [63:0] _queues_114_io_addressOut_bits;
	wire _queues_113_io_addressOut_valid;
	wire [63:0] _queues_113_io_addressOut_bits;
	wire _queues_112_io_addressOut_valid;
	wire [63:0] _queues_112_io_addressOut_bits;
	wire _queues_111_io_addressOut_valid;
	wire [63:0] _queues_111_io_addressOut_bits;
	wire _queues_110_io_addressOut_valid;
	wire [63:0] _queues_110_io_addressOut_bits;
	wire _queues_109_io_addressOut_valid;
	wire [63:0] _queues_109_io_addressOut_bits;
	wire _queues_108_io_addressOut_valid;
	wire [63:0] _queues_108_io_addressOut_bits;
	wire _queues_107_io_addressOut_valid;
	wire [63:0] _queues_107_io_addressOut_bits;
	wire _queues_106_io_addressOut_valid;
	wire [63:0] _queues_106_io_addressOut_bits;
	wire _queues_105_io_addressOut_valid;
	wire [63:0] _queues_105_io_addressOut_bits;
	wire _queues_104_io_addressOut_valid;
	wire [63:0] _queues_104_io_addressOut_bits;
	wire _queues_103_io_addressOut_valid;
	wire [63:0] _queues_103_io_addressOut_bits;
	wire _queues_102_io_addressOut_valid;
	wire [63:0] _queues_102_io_addressOut_bits;
	wire _queues_101_io_addressOut_valid;
	wire [63:0] _queues_101_io_addressOut_bits;
	wire _queues_100_io_addressOut_valid;
	wire [63:0] _queues_100_io_addressOut_bits;
	wire _queues_99_io_addressOut_valid;
	wire [63:0] _queues_99_io_addressOut_bits;
	wire _queues_98_io_addressOut_valid;
	wire [63:0] _queues_98_io_addressOut_bits;
	wire _queues_97_io_addressOut_valid;
	wire [63:0] _queues_97_io_addressOut_bits;
	wire _queues_96_io_addressOut_valid;
	wire [63:0] _queues_96_io_addressOut_bits;
	wire _queues_95_io_addressOut_valid;
	wire [63:0] _queues_95_io_addressOut_bits;
	wire _queues_94_io_addressOut_valid;
	wire [63:0] _queues_94_io_addressOut_bits;
	wire _queues_93_io_addressOut_valid;
	wire [63:0] _queues_93_io_addressOut_bits;
	wire _queues_92_io_addressOut_valid;
	wire [63:0] _queues_92_io_addressOut_bits;
	wire _queues_91_io_addressOut_valid;
	wire [63:0] _queues_91_io_addressOut_bits;
	wire _queues_90_io_addressOut_valid;
	wire [63:0] _queues_90_io_addressOut_bits;
	wire _queues_89_io_addressOut_valid;
	wire [63:0] _queues_89_io_addressOut_bits;
	wire _queues_88_io_addressOut_valid;
	wire [63:0] _queues_88_io_addressOut_bits;
	wire _queues_87_io_addressOut_valid;
	wire [63:0] _queues_87_io_addressOut_bits;
	wire _queues_86_io_addressOut_valid;
	wire [63:0] _queues_86_io_addressOut_bits;
	wire _queues_85_io_addressOut_valid;
	wire [63:0] _queues_85_io_addressOut_bits;
	wire _queues_84_io_addressOut_valid;
	wire [63:0] _queues_84_io_addressOut_bits;
	wire _queues_83_io_addressOut_valid;
	wire [63:0] _queues_83_io_addressOut_bits;
	wire _queues_82_io_addressOut_valid;
	wire [63:0] _queues_82_io_addressOut_bits;
	wire _queues_81_io_addressOut_valid;
	wire [63:0] _queues_81_io_addressOut_bits;
	wire _queues_80_io_addressOut_valid;
	wire [63:0] _queues_80_io_addressOut_bits;
	wire _queues_79_io_addressOut_valid;
	wire [63:0] _queues_79_io_addressOut_bits;
	wire _queues_78_io_addressOut_valid;
	wire [63:0] _queues_78_io_addressOut_bits;
	wire _queues_77_io_addressOut_valid;
	wire [63:0] _queues_77_io_addressOut_bits;
	wire _queues_76_io_addressOut_valid;
	wire [63:0] _queues_76_io_addressOut_bits;
	wire _queues_75_io_addressOut_valid;
	wire [63:0] _queues_75_io_addressOut_bits;
	wire _queues_74_io_addressOut_valid;
	wire [63:0] _queues_74_io_addressOut_bits;
	wire _queues_73_io_addressOut_valid;
	wire [63:0] _queues_73_io_addressOut_bits;
	wire _queues_72_io_addressOut_valid;
	wire [63:0] _queues_72_io_addressOut_bits;
	wire _queues_71_io_addressOut_valid;
	wire [63:0] _queues_71_io_addressOut_bits;
	wire _queues_70_io_addressOut_valid;
	wire [63:0] _queues_70_io_addressOut_bits;
	wire _queues_69_io_addressOut_valid;
	wire [63:0] _queues_69_io_addressOut_bits;
	wire _queues_68_io_addressOut_valid;
	wire [63:0] _queues_68_io_addressOut_bits;
	wire _queues_67_io_addressOut_valid;
	wire [63:0] _queues_67_io_addressOut_bits;
	wire _queues_66_io_addressOut_valid;
	wire [63:0] _queues_66_io_addressOut_bits;
	wire _queues_65_io_addressOut_valid;
	wire [63:0] _queues_65_io_addressOut_bits;
	wire _queues_64_io_addressOut_valid;
	wire [63:0] _queues_64_io_addressOut_bits;
	wire _queues_63_io_addressOut_valid;
	wire [63:0] _queues_63_io_addressOut_bits;
	wire _queues_62_io_addressOut_valid;
	wire [63:0] _queues_62_io_addressOut_bits;
	wire _queues_61_io_addressOut_valid;
	wire [63:0] _queues_61_io_addressOut_bits;
	wire _queues_60_io_addressOut_valid;
	wire [63:0] _queues_60_io_addressOut_bits;
	wire _queues_59_io_addressOut_valid;
	wire [63:0] _queues_59_io_addressOut_bits;
	wire _queues_58_io_addressOut_valid;
	wire [63:0] _queues_58_io_addressOut_bits;
	wire _queues_57_io_addressOut_valid;
	wire [63:0] _queues_57_io_addressOut_bits;
	wire _queues_56_io_addressOut_valid;
	wire [63:0] _queues_56_io_addressOut_bits;
	wire _queues_55_io_addressOut_valid;
	wire [63:0] _queues_55_io_addressOut_bits;
	wire _queues_54_io_addressOut_valid;
	wire [63:0] _queues_54_io_addressOut_bits;
	wire _queues_53_io_addressOut_valid;
	wire [63:0] _queues_53_io_addressOut_bits;
	wire _queues_52_io_addressOut_valid;
	wire [63:0] _queues_52_io_addressOut_bits;
	wire _queues_51_io_addressOut_valid;
	wire [63:0] _queues_51_io_addressOut_bits;
	wire _queues_50_io_addressOut_valid;
	wire [63:0] _queues_50_io_addressOut_bits;
	wire _queues_49_io_addressOut_valid;
	wire [63:0] _queues_49_io_addressOut_bits;
	wire _queues_48_io_addressOut_valid;
	wire [63:0] _queues_48_io_addressOut_bits;
	wire _queues_47_io_addressOut_valid;
	wire [63:0] _queues_47_io_addressOut_bits;
	wire _queues_46_io_addressOut_valid;
	wire [63:0] _queues_46_io_addressOut_bits;
	wire _queues_45_io_addressOut_valid;
	wire [63:0] _queues_45_io_addressOut_bits;
	wire _queues_44_io_addressOut_valid;
	wire [63:0] _queues_44_io_addressOut_bits;
	wire _queues_43_io_addressOut_valid;
	wire [63:0] _queues_43_io_addressOut_bits;
	wire _queues_42_io_addressOut_valid;
	wire [63:0] _queues_42_io_addressOut_bits;
	wire _queues_41_io_addressOut_valid;
	wire [63:0] _queues_41_io_addressOut_bits;
	wire _queues_40_io_addressOut_valid;
	wire [63:0] _queues_40_io_addressOut_bits;
	wire _queues_39_io_addressOut_valid;
	wire [63:0] _queues_39_io_addressOut_bits;
	wire _queues_38_io_addressOut_valid;
	wire [63:0] _queues_38_io_addressOut_bits;
	wire _queues_37_io_addressOut_valid;
	wire [63:0] _queues_37_io_addressOut_bits;
	wire _queues_36_io_addressOut_valid;
	wire [63:0] _queues_36_io_addressOut_bits;
	wire _queues_35_io_addressOut_valid;
	wire [63:0] _queues_35_io_addressOut_bits;
	wire _queues_34_io_addressOut_valid;
	wire [63:0] _queues_34_io_addressOut_bits;
	wire _queues_33_io_addressOut_valid;
	wire [63:0] _queues_33_io_addressOut_bits;
	wire _queues_32_io_addressOut_valid;
	wire [63:0] _queues_32_io_addressOut_bits;
	wire _queues_31_io_addressOut_valid;
	wire [63:0] _queues_31_io_addressOut_bits;
	wire _queues_30_io_addressOut_valid;
	wire [63:0] _queues_30_io_addressOut_bits;
	wire _queues_29_io_addressOut_valid;
	wire [63:0] _queues_29_io_addressOut_bits;
	wire _queues_28_io_addressOut_valid;
	wire [63:0] _queues_28_io_addressOut_bits;
	wire _queues_27_io_addressOut_valid;
	wire [63:0] _queues_27_io_addressOut_bits;
	wire _queues_26_io_addressOut_valid;
	wire [63:0] _queues_26_io_addressOut_bits;
	wire _queues_25_io_addressOut_valid;
	wire [63:0] _queues_25_io_addressOut_bits;
	wire _queues_24_io_addressOut_valid;
	wire [63:0] _queues_24_io_addressOut_bits;
	wire _queues_23_io_addressOut_valid;
	wire [63:0] _queues_23_io_addressOut_bits;
	wire _queues_22_io_addressOut_valid;
	wire [63:0] _queues_22_io_addressOut_bits;
	wire _queues_21_io_addressOut_valid;
	wire [63:0] _queues_21_io_addressOut_bits;
	wire _queues_20_io_addressOut_valid;
	wire [63:0] _queues_20_io_addressOut_bits;
	wire _queues_19_io_addressOut_valid;
	wire [63:0] _queues_19_io_addressOut_bits;
	wire _queues_18_io_addressOut_valid;
	wire [63:0] _queues_18_io_addressOut_bits;
	wire _queues_17_io_addressOut_valid;
	wire [63:0] _queues_17_io_addressOut_bits;
	wire _queues_16_io_addressOut_valid;
	wire [63:0] _queues_16_io_addressOut_bits;
	wire _queues_15_io_addressOut_valid;
	wire [63:0] _queues_15_io_addressOut_bits;
	wire _queues_14_io_addressOut_valid;
	wire [63:0] _queues_14_io_addressOut_bits;
	wire _queues_13_io_addressOut_valid;
	wire [63:0] _queues_13_io_addressOut_bits;
	wire _queues_12_io_addressOut_valid;
	wire [63:0] _queues_12_io_addressOut_bits;
	wire _queues_11_io_addressOut_valid;
	wire [63:0] _queues_11_io_addressOut_bits;
	wire _queues_10_io_addressOut_valid;
	wire [63:0] _queues_10_io_addressOut_bits;
	wire _queues_9_io_addressOut_valid;
	wire [63:0] _queues_9_io_addressOut_bits;
	wire _queues_8_io_addressOut_valid;
	wire [63:0] _queues_8_io_addressOut_bits;
	wire _queues_7_io_addressOut_valid;
	wire [63:0] _queues_7_io_addressOut_bits;
	wire _queues_6_io_addressOut_valid;
	wire [63:0] _queues_6_io_addressOut_bits;
	wire _queues_5_io_addressOut_valid;
	wire [63:0] _queues_5_io_addressOut_bits;
	wire _queues_4_io_addressOut_valid;
	wire [63:0] _queues_4_io_addressOut_bits;
	wire _queues_3_io_addressOut_valid;
	wire [63:0] _queues_3_io_addressOut_bits;
	wire _queues_2_io_addressOut_valid;
	wire [63:0] _queues_2_io_addressOut_bits;
	wire _queues_1_io_addressOut_valid;
	wire [63:0] _queues_1_io_addressOut_bits;
	wire _queues_0_io_addressOut_valid;
	wire [63:0] _queues_0_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_15_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_15_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_15_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_14_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_14_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_14_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_13_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_13_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_13_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_12_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_12_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_12_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_11_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_11_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_11_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_10_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_10_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_10_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_9_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_9_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_9_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_8_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_8_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_8_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_7_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_7_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_7_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_6_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_6_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_6_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_5_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_5_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_5_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_4_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_4_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_4_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_3_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_3_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_3_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_2_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_2_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_2_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_1_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_1_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_1_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_io_addressIn_ready;
	wire _networkUnits_127_io_peAddress_ready;
	wire _networkUnits_127_io_addressOut_valid;
	wire [63:0] _networkUnits_127_io_addressOut_bits;
	wire _networkUnits_126_io_addressIn_ready;
	wire _networkUnits_126_io_peAddress_ready;
	wire _networkUnits_126_io_addressOut_valid;
	wire [63:0] _networkUnits_126_io_addressOut_bits;
	wire _networkUnits_125_io_addressIn_ready;
	wire _networkUnits_125_io_peAddress_ready;
	wire _networkUnits_125_io_addressOut_valid;
	wire [63:0] _networkUnits_125_io_addressOut_bits;
	wire _networkUnits_124_io_addressIn_ready;
	wire _networkUnits_124_io_peAddress_ready;
	wire _networkUnits_124_io_addressOut_valid;
	wire [63:0] _networkUnits_124_io_addressOut_bits;
	wire _networkUnits_123_io_addressIn_ready;
	wire _networkUnits_123_io_peAddress_ready;
	wire _networkUnits_123_io_addressOut_valid;
	wire [63:0] _networkUnits_123_io_addressOut_bits;
	wire _networkUnits_122_io_addressIn_ready;
	wire _networkUnits_122_io_peAddress_ready;
	wire _networkUnits_122_io_addressOut_valid;
	wire [63:0] _networkUnits_122_io_addressOut_bits;
	wire _networkUnits_121_io_addressIn_ready;
	wire _networkUnits_121_io_peAddress_ready;
	wire _networkUnits_121_io_addressOut_valid;
	wire [63:0] _networkUnits_121_io_addressOut_bits;
	wire _networkUnits_120_io_addressIn_ready;
	wire _networkUnits_120_io_peAddress_ready;
	wire _networkUnits_120_io_addressOut_valid;
	wire [63:0] _networkUnits_120_io_addressOut_bits;
	wire _networkUnits_119_io_addressIn_ready;
	wire _networkUnits_119_io_peAddress_ready;
	wire _networkUnits_119_io_addressOut_valid;
	wire [63:0] _networkUnits_119_io_addressOut_bits;
	wire _networkUnits_118_io_addressIn_ready;
	wire _networkUnits_118_io_peAddress_ready;
	wire _networkUnits_118_io_addressOut_valid;
	wire [63:0] _networkUnits_118_io_addressOut_bits;
	wire _networkUnits_117_io_addressIn_ready;
	wire _networkUnits_117_io_peAddress_ready;
	wire _networkUnits_117_io_addressOut_valid;
	wire [63:0] _networkUnits_117_io_addressOut_bits;
	wire _networkUnits_116_io_addressIn_ready;
	wire _networkUnits_116_io_peAddress_ready;
	wire _networkUnits_116_io_addressOut_valid;
	wire [63:0] _networkUnits_116_io_addressOut_bits;
	wire _networkUnits_115_io_addressIn_ready;
	wire _networkUnits_115_io_peAddress_ready;
	wire _networkUnits_115_io_addressOut_valid;
	wire [63:0] _networkUnits_115_io_addressOut_bits;
	wire _networkUnits_114_io_addressIn_ready;
	wire _networkUnits_114_io_peAddress_ready;
	wire _networkUnits_114_io_addressOut_valid;
	wire [63:0] _networkUnits_114_io_addressOut_bits;
	wire _networkUnits_113_io_addressIn_ready;
	wire _networkUnits_113_io_peAddress_ready;
	wire _networkUnits_113_io_addressOut_valid;
	wire [63:0] _networkUnits_113_io_addressOut_bits;
	wire _networkUnits_112_io_addressIn_ready;
	wire _networkUnits_112_io_peAddress_ready;
	wire _networkUnits_112_io_addressOut_valid;
	wire [63:0] _networkUnits_112_io_addressOut_bits;
	wire _networkUnits_111_io_addressIn_ready;
	wire _networkUnits_111_io_peAddress_ready;
	wire _networkUnits_111_io_addressOut_valid;
	wire [63:0] _networkUnits_111_io_addressOut_bits;
	wire _networkUnits_110_io_addressIn_ready;
	wire _networkUnits_110_io_peAddress_ready;
	wire _networkUnits_110_io_addressOut_valid;
	wire [63:0] _networkUnits_110_io_addressOut_bits;
	wire _networkUnits_109_io_addressIn_ready;
	wire _networkUnits_109_io_peAddress_ready;
	wire _networkUnits_109_io_addressOut_valid;
	wire [63:0] _networkUnits_109_io_addressOut_bits;
	wire _networkUnits_108_io_addressIn_ready;
	wire _networkUnits_108_io_peAddress_ready;
	wire _networkUnits_108_io_addressOut_valid;
	wire [63:0] _networkUnits_108_io_addressOut_bits;
	wire _networkUnits_107_io_addressIn_ready;
	wire _networkUnits_107_io_peAddress_ready;
	wire _networkUnits_107_io_addressOut_valid;
	wire [63:0] _networkUnits_107_io_addressOut_bits;
	wire _networkUnits_106_io_addressIn_ready;
	wire _networkUnits_106_io_peAddress_ready;
	wire _networkUnits_106_io_addressOut_valid;
	wire [63:0] _networkUnits_106_io_addressOut_bits;
	wire _networkUnits_105_io_addressIn_ready;
	wire _networkUnits_105_io_peAddress_ready;
	wire _networkUnits_105_io_addressOut_valid;
	wire [63:0] _networkUnits_105_io_addressOut_bits;
	wire _networkUnits_104_io_addressIn_ready;
	wire _networkUnits_104_io_peAddress_ready;
	wire _networkUnits_104_io_addressOut_valid;
	wire [63:0] _networkUnits_104_io_addressOut_bits;
	wire _networkUnits_103_io_addressIn_ready;
	wire _networkUnits_103_io_peAddress_ready;
	wire _networkUnits_103_io_addressOut_valid;
	wire [63:0] _networkUnits_103_io_addressOut_bits;
	wire _networkUnits_102_io_addressIn_ready;
	wire _networkUnits_102_io_peAddress_ready;
	wire _networkUnits_102_io_addressOut_valid;
	wire [63:0] _networkUnits_102_io_addressOut_bits;
	wire _networkUnits_101_io_addressIn_ready;
	wire _networkUnits_101_io_peAddress_ready;
	wire _networkUnits_101_io_addressOut_valid;
	wire [63:0] _networkUnits_101_io_addressOut_bits;
	wire _networkUnits_100_io_addressIn_ready;
	wire _networkUnits_100_io_peAddress_ready;
	wire _networkUnits_100_io_addressOut_valid;
	wire [63:0] _networkUnits_100_io_addressOut_bits;
	wire _networkUnits_99_io_addressIn_ready;
	wire _networkUnits_99_io_peAddress_ready;
	wire _networkUnits_99_io_addressOut_valid;
	wire [63:0] _networkUnits_99_io_addressOut_bits;
	wire _networkUnits_98_io_addressIn_ready;
	wire _networkUnits_98_io_peAddress_ready;
	wire _networkUnits_98_io_addressOut_valid;
	wire [63:0] _networkUnits_98_io_addressOut_bits;
	wire _networkUnits_97_io_addressIn_ready;
	wire _networkUnits_97_io_peAddress_ready;
	wire _networkUnits_97_io_addressOut_valid;
	wire [63:0] _networkUnits_97_io_addressOut_bits;
	wire _networkUnits_96_io_addressIn_ready;
	wire _networkUnits_96_io_peAddress_ready;
	wire _networkUnits_96_io_addressOut_valid;
	wire [63:0] _networkUnits_96_io_addressOut_bits;
	wire _networkUnits_95_io_addressIn_ready;
	wire _networkUnits_95_io_peAddress_ready;
	wire _networkUnits_95_io_addressOut_valid;
	wire [63:0] _networkUnits_95_io_addressOut_bits;
	wire _networkUnits_94_io_addressIn_ready;
	wire _networkUnits_94_io_peAddress_ready;
	wire _networkUnits_94_io_addressOut_valid;
	wire [63:0] _networkUnits_94_io_addressOut_bits;
	wire _networkUnits_93_io_addressIn_ready;
	wire _networkUnits_93_io_peAddress_ready;
	wire _networkUnits_93_io_addressOut_valid;
	wire [63:0] _networkUnits_93_io_addressOut_bits;
	wire _networkUnits_92_io_addressIn_ready;
	wire _networkUnits_92_io_peAddress_ready;
	wire _networkUnits_92_io_addressOut_valid;
	wire [63:0] _networkUnits_92_io_addressOut_bits;
	wire _networkUnits_91_io_addressIn_ready;
	wire _networkUnits_91_io_peAddress_ready;
	wire _networkUnits_91_io_addressOut_valid;
	wire [63:0] _networkUnits_91_io_addressOut_bits;
	wire _networkUnits_90_io_addressIn_ready;
	wire _networkUnits_90_io_peAddress_ready;
	wire _networkUnits_90_io_addressOut_valid;
	wire [63:0] _networkUnits_90_io_addressOut_bits;
	wire _networkUnits_89_io_addressIn_ready;
	wire _networkUnits_89_io_peAddress_ready;
	wire _networkUnits_89_io_addressOut_valid;
	wire [63:0] _networkUnits_89_io_addressOut_bits;
	wire _networkUnits_88_io_addressIn_ready;
	wire _networkUnits_88_io_peAddress_ready;
	wire _networkUnits_88_io_addressOut_valid;
	wire [63:0] _networkUnits_88_io_addressOut_bits;
	wire _networkUnits_87_io_addressIn_ready;
	wire _networkUnits_87_io_peAddress_ready;
	wire _networkUnits_87_io_addressOut_valid;
	wire [63:0] _networkUnits_87_io_addressOut_bits;
	wire _networkUnits_86_io_addressIn_ready;
	wire _networkUnits_86_io_peAddress_ready;
	wire _networkUnits_86_io_addressOut_valid;
	wire [63:0] _networkUnits_86_io_addressOut_bits;
	wire _networkUnits_85_io_addressIn_ready;
	wire _networkUnits_85_io_peAddress_ready;
	wire _networkUnits_85_io_addressOut_valid;
	wire [63:0] _networkUnits_85_io_addressOut_bits;
	wire _networkUnits_84_io_addressIn_ready;
	wire _networkUnits_84_io_peAddress_ready;
	wire _networkUnits_84_io_addressOut_valid;
	wire [63:0] _networkUnits_84_io_addressOut_bits;
	wire _networkUnits_83_io_addressIn_ready;
	wire _networkUnits_83_io_peAddress_ready;
	wire _networkUnits_83_io_addressOut_valid;
	wire [63:0] _networkUnits_83_io_addressOut_bits;
	wire _networkUnits_82_io_addressIn_ready;
	wire _networkUnits_82_io_peAddress_ready;
	wire _networkUnits_82_io_addressOut_valid;
	wire [63:0] _networkUnits_82_io_addressOut_bits;
	wire _networkUnits_81_io_addressIn_ready;
	wire _networkUnits_81_io_peAddress_ready;
	wire _networkUnits_81_io_addressOut_valid;
	wire [63:0] _networkUnits_81_io_addressOut_bits;
	wire _networkUnits_80_io_addressIn_ready;
	wire _networkUnits_80_io_peAddress_ready;
	wire _networkUnits_80_io_addressOut_valid;
	wire [63:0] _networkUnits_80_io_addressOut_bits;
	wire _networkUnits_79_io_addressIn_ready;
	wire _networkUnits_79_io_peAddress_ready;
	wire _networkUnits_79_io_addressOut_valid;
	wire [63:0] _networkUnits_79_io_addressOut_bits;
	wire _networkUnits_78_io_addressIn_ready;
	wire _networkUnits_78_io_peAddress_ready;
	wire _networkUnits_78_io_addressOut_valid;
	wire [63:0] _networkUnits_78_io_addressOut_bits;
	wire _networkUnits_77_io_addressIn_ready;
	wire _networkUnits_77_io_peAddress_ready;
	wire _networkUnits_77_io_addressOut_valid;
	wire [63:0] _networkUnits_77_io_addressOut_bits;
	wire _networkUnits_76_io_addressIn_ready;
	wire _networkUnits_76_io_peAddress_ready;
	wire _networkUnits_76_io_addressOut_valid;
	wire [63:0] _networkUnits_76_io_addressOut_bits;
	wire _networkUnits_75_io_addressIn_ready;
	wire _networkUnits_75_io_peAddress_ready;
	wire _networkUnits_75_io_addressOut_valid;
	wire [63:0] _networkUnits_75_io_addressOut_bits;
	wire _networkUnits_74_io_addressIn_ready;
	wire _networkUnits_74_io_peAddress_ready;
	wire _networkUnits_74_io_addressOut_valid;
	wire [63:0] _networkUnits_74_io_addressOut_bits;
	wire _networkUnits_73_io_addressIn_ready;
	wire _networkUnits_73_io_peAddress_ready;
	wire _networkUnits_73_io_addressOut_valid;
	wire [63:0] _networkUnits_73_io_addressOut_bits;
	wire _networkUnits_72_io_addressIn_ready;
	wire _networkUnits_72_io_peAddress_ready;
	wire _networkUnits_72_io_addressOut_valid;
	wire [63:0] _networkUnits_72_io_addressOut_bits;
	wire _networkUnits_71_io_addressIn_ready;
	wire _networkUnits_71_io_peAddress_ready;
	wire _networkUnits_71_io_addressOut_valid;
	wire [63:0] _networkUnits_71_io_addressOut_bits;
	wire _networkUnits_70_io_addressIn_ready;
	wire _networkUnits_70_io_peAddress_ready;
	wire _networkUnits_70_io_addressOut_valid;
	wire [63:0] _networkUnits_70_io_addressOut_bits;
	wire _networkUnits_69_io_addressIn_ready;
	wire _networkUnits_69_io_peAddress_ready;
	wire _networkUnits_69_io_addressOut_valid;
	wire [63:0] _networkUnits_69_io_addressOut_bits;
	wire _networkUnits_68_io_addressIn_ready;
	wire _networkUnits_68_io_peAddress_ready;
	wire _networkUnits_68_io_addressOut_valid;
	wire [63:0] _networkUnits_68_io_addressOut_bits;
	wire _networkUnits_67_io_addressIn_ready;
	wire _networkUnits_67_io_peAddress_ready;
	wire _networkUnits_67_io_addressOut_valid;
	wire [63:0] _networkUnits_67_io_addressOut_bits;
	wire _networkUnits_66_io_addressIn_ready;
	wire _networkUnits_66_io_peAddress_ready;
	wire _networkUnits_66_io_addressOut_valid;
	wire [63:0] _networkUnits_66_io_addressOut_bits;
	wire _networkUnits_65_io_addressIn_ready;
	wire _networkUnits_65_io_peAddress_ready;
	wire _networkUnits_65_io_addressOut_valid;
	wire [63:0] _networkUnits_65_io_addressOut_bits;
	wire _networkUnits_64_io_addressIn_ready;
	wire _networkUnits_64_io_peAddress_ready;
	wire _networkUnits_64_io_addressOut_valid;
	wire [63:0] _networkUnits_64_io_addressOut_bits;
	wire _networkUnits_63_io_addressIn_ready;
	wire _networkUnits_63_io_peAddress_ready;
	wire _networkUnits_63_io_addressOut_valid;
	wire [63:0] _networkUnits_63_io_addressOut_bits;
	wire _networkUnits_62_io_addressIn_ready;
	wire _networkUnits_62_io_peAddress_ready;
	wire _networkUnits_62_io_addressOut_valid;
	wire [63:0] _networkUnits_62_io_addressOut_bits;
	wire _networkUnits_61_io_addressIn_ready;
	wire _networkUnits_61_io_peAddress_ready;
	wire _networkUnits_61_io_addressOut_valid;
	wire [63:0] _networkUnits_61_io_addressOut_bits;
	wire _networkUnits_60_io_addressIn_ready;
	wire _networkUnits_60_io_peAddress_ready;
	wire _networkUnits_60_io_addressOut_valid;
	wire [63:0] _networkUnits_60_io_addressOut_bits;
	wire _networkUnits_59_io_addressIn_ready;
	wire _networkUnits_59_io_peAddress_ready;
	wire _networkUnits_59_io_addressOut_valid;
	wire [63:0] _networkUnits_59_io_addressOut_bits;
	wire _networkUnits_58_io_addressIn_ready;
	wire _networkUnits_58_io_peAddress_ready;
	wire _networkUnits_58_io_addressOut_valid;
	wire [63:0] _networkUnits_58_io_addressOut_bits;
	wire _networkUnits_57_io_addressIn_ready;
	wire _networkUnits_57_io_peAddress_ready;
	wire _networkUnits_57_io_addressOut_valid;
	wire [63:0] _networkUnits_57_io_addressOut_bits;
	wire _networkUnits_56_io_addressIn_ready;
	wire _networkUnits_56_io_peAddress_ready;
	wire _networkUnits_56_io_addressOut_valid;
	wire [63:0] _networkUnits_56_io_addressOut_bits;
	wire _networkUnits_55_io_addressIn_ready;
	wire _networkUnits_55_io_peAddress_ready;
	wire _networkUnits_55_io_addressOut_valid;
	wire [63:0] _networkUnits_55_io_addressOut_bits;
	wire _networkUnits_54_io_addressIn_ready;
	wire _networkUnits_54_io_peAddress_ready;
	wire _networkUnits_54_io_addressOut_valid;
	wire [63:0] _networkUnits_54_io_addressOut_bits;
	wire _networkUnits_53_io_addressIn_ready;
	wire _networkUnits_53_io_peAddress_ready;
	wire _networkUnits_53_io_addressOut_valid;
	wire [63:0] _networkUnits_53_io_addressOut_bits;
	wire _networkUnits_52_io_addressIn_ready;
	wire _networkUnits_52_io_peAddress_ready;
	wire _networkUnits_52_io_addressOut_valid;
	wire [63:0] _networkUnits_52_io_addressOut_bits;
	wire _networkUnits_51_io_addressIn_ready;
	wire _networkUnits_51_io_peAddress_ready;
	wire _networkUnits_51_io_addressOut_valid;
	wire [63:0] _networkUnits_51_io_addressOut_bits;
	wire _networkUnits_50_io_addressIn_ready;
	wire _networkUnits_50_io_peAddress_ready;
	wire _networkUnits_50_io_addressOut_valid;
	wire [63:0] _networkUnits_50_io_addressOut_bits;
	wire _networkUnits_49_io_addressIn_ready;
	wire _networkUnits_49_io_peAddress_ready;
	wire _networkUnits_49_io_addressOut_valid;
	wire [63:0] _networkUnits_49_io_addressOut_bits;
	wire _networkUnits_48_io_addressIn_ready;
	wire _networkUnits_48_io_peAddress_ready;
	wire _networkUnits_48_io_addressOut_valid;
	wire [63:0] _networkUnits_48_io_addressOut_bits;
	wire _networkUnits_47_io_addressIn_ready;
	wire _networkUnits_47_io_peAddress_ready;
	wire _networkUnits_47_io_addressOut_valid;
	wire [63:0] _networkUnits_47_io_addressOut_bits;
	wire _networkUnits_46_io_addressIn_ready;
	wire _networkUnits_46_io_peAddress_ready;
	wire _networkUnits_46_io_addressOut_valid;
	wire [63:0] _networkUnits_46_io_addressOut_bits;
	wire _networkUnits_45_io_addressIn_ready;
	wire _networkUnits_45_io_peAddress_ready;
	wire _networkUnits_45_io_addressOut_valid;
	wire [63:0] _networkUnits_45_io_addressOut_bits;
	wire _networkUnits_44_io_addressIn_ready;
	wire _networkUnits_44_io_peAddress_ready;
	wire _networkUnits_44_io_addressOut_valid;
	wire [63:0] _networkUnits_44_io_addressOut_bits;
	wire _networkUnits_43_io_addressIn_ready;
	wire _networkUnits_43_io_peAddress_ready;
	wire _networkUnits_43_io_addressOut_valid;
	wire [63:0] _networkUnits_43_io_addressOut_bits;
	wire _networkUnits_42_io_addressIn_ready;
	wire _networkUnits_42_io_peAddress_ready;
	wire _networkUnits_42_io_addressOut_valid;
	wire [63:0] _networkUnits_42_io_addressOut_bits;
	wire _networkUnits_41_io_addressIn_ready;
	wire _networkUnits_41_io_peAddress_ready;
	wire _networkUnits_41_io_addressOut_valid;
	wire [63:0] _networkUnits_41_io_addressOut_bits;
	wire _networkUnits_40_io_addressIn_ready;
	wire _networkUnits_40_io_peAddress_ready;
	wire _networkUnits_40_io_addressOut_valid;
	wire [63:0] _networkUnits_40_io_addressOut_bits;
	wire _networkUnits_39_io_addressIn_ready;
	wire _networkUnits_39_io_peAddress_ready;
	wire _networkUnits_39_io_addressOut_valid;
	wire [63:0] _networkUnits_39_io_addressOut_bits;
	wire _networkUnits_38_io_addressIn_ready;
	wire _networkUnits_38_io_peAddress_ready;
	wire _networkUnits_38_io_addressOut_valid;
	wire [63:0] _networkUnits_38_io_addressOut_bits;
	wire _networkUnits_37_io_addressIn_ready;
	wire _networkUnits_37_io_peAddress_ready;
	wire _networkUnits_37_io_addressOut_valid;
	wire [63:0] _networkUnits_37_io_addressOut_bits;
	wire _networkUnits_36_io_addressIn_ready;
	wire _networkUnits_36_io_peAddress_ready;
	wire _networkUnits_36_io_addressOut_valid;
	wire [63:0] _networkUnits_36_io_addressOut_bits;
	wire _networkUnits_35_io_addressIn_ready;
	wire _networkUnits_35_io_peAddress_ready;
	wire _networkUnits_35_io_addressOut_valid;
	wire [63:0] _networkUnits_35_io_addressOut_bits;
	wire _networkUnits_34_io_addressIn_ready;
	wire _networkUnits_34_io_peAddress_ready;
	wire _networkUnits_34_io_addressOut_valid;
	wire [63:0] _networkUnits_34_io_addressOut_bits;
	wire _networkUnits_33_io_addressIn_ready;
	wire _networkUnits_33_io_peAddress_ready;
	wire _networkUnits_33_io_addressOut_valid;
	wire [63:0] _networkUnits_33_io_addressOut_bits;
	wire _networkUnits_32_io_addressIn_ready;
	wire _networkUnits_32_io_peAddress_ready;
	wire _networkUnits_32_io_addressOut_valid;
	wire [63:0] _networkUnits_32_io_addressOut_bits;
	wire _networkUnits_31_io_addressIn_ready;
	wire _networkUnits_31_io_peAddress_ready;
	wire _networkUnits_31_io_addressOut_valid;
	wire [63:0] _networkUnits_31_io_addressOut_bits;
	wire _networkUnits_30_io_addressIn_ready;
	wire _networkUnits_30_io_peAddress_ready;
	wire _networkUnits_30_io_addressOut_valid;
	wire [63:0] _networkUnits_30_io_addressOut_bits;
	wire _networkUnits_29_io_addressIn_ready;
	wire _networkUnits_29_io_peAddress_ready;
	wire _networkUnits_29_io_addressOut_valid;
	wire [63:0] _networkUnits_29_io_addressOut_bits;
	wire _networkUnits_28_io_addressIn_ready;
	wire _networkUnits_28_io_peAddress_ready;
	wire _networkUnits_28_io_addressOut_valid;
	wire [63:0] _networkUnits_28_io_addressOut_bits;
	wire _networkUnits_27_io_addressIn_ready;
	wire _networkUnits_27_io_peAddress_ready;
	wire _networkUnits_27_io_addressOut_valid;
	wire [63:0] _networkUnits_27_io_addressOut_bits;
	wire _networkUnits_26_io_addressIn_ready;
	wire _networkUnits_26_io_peAddress_ready;
	wire _networkUnits_26_io_addressOut_valid;
	wire [63:0] _networkUnits_26_io_addressOut_bits;
	wire _networkUnits_25_io_addressIn_ready;
	wire _networkUnits_25_io_peAddress_ready;
	wire _networkUnits_25_io_addressOut_valid;
	wire [63:0] _networkUnits_25_io_addressOut_bits;
	wire _networkUnits_24_io_addressIn_ready;
	wire _networkUnits_24_io_peAddress_ready;
	wire _networkUnits_24_io_addressOut_valid;
	wire [63:0] _networkUnits_24_io_addressOut_bits;
	wire _networkUnits_23_io_addressIn_ready;
	wire _networkUnits_23_io_peAddress_ready;
	wire _networkUnits_23_io_addressOut_valid;
	wire [63:0] _networkUnits_23_io_addressOut_bits;
	wire _networkUnits_22_io_addressIn_ready;
	wire _networkUnits_22_io_peAddress_ready;
	wire _networkUnits_22_io_addressOut_valid;
	wire [63:0] _networkUnits_22_io_addressOut_bits;
	wire _networkUnits_21_io_addressIn_ready;
	wire _networkUnits_21_io_peAddress_ready;
	wire _networkUnits_21_io_addressOut_valid;
	wire [63:0] _networkUnits_21_io_addressOut_bits;
	wire _networkUnits_20_io_addressIn_ready;
	wire _networkUnits_20_io_peAddress_ready;
	wire _networkUnits_20_io_addressOut_valid;
	wire [63:0] _networkUnits_20_io_addressOut_bits;
	wire _networkUnits_19_io_addressIn_ready;
	wire _networkUnits_19_io_peAddress_ready;
	wire _networkUnits_19_io_addressOut_valid;
	wire [63:0] _networkUnits_19_io_addressOut_bits;
	wire _networkUnits_18_io_addressIn_ready;
	wire _networkUnits_18_io_peAddress_ready;
	wire _networkUnits_18_io_addressOut_valid;
	wire [63:0] _networkUnits_18_io_addressOut_bits;
	wire _networkUnits_17_io_addressIn_ready;
	wire _networkUnits_17_io_peAddress_ready;
	wire _networkUnits_17_io_addressOut_valid;
	wire [63:0] _networkUnits_17_io_addressOut_bits;
	wire _networkUnits_16_io_addressIn_ready;
	wire _networkUnits_16_io_peAddress_ready;
	wire _networkUnits_16_io_addressOut_valid;
	wire [63:0] _networkUnits_16_io_addressOut_bits;
	wire _networkUnits_15_io_addressIn_ready;
	wire _networkUnits_15_io_peAddress_ready;
	wire _networkUnits_15_io_addressOut_valid;
	wire [63:0] _networkUnits_15_io_addressOut_bits;
	wire _networkUnits_14_io_addressIn_ready;
	wire _networkUnits_14_io_peAddress_ready;
	wire _networkUnits_14_io_addressOut_valid;
	wire [63:0] _networkUnits_14_io_addressOut_bits;
	wire _networkUnits_13_io_addressIn_ready;
	wire _networkUnits_13_io_peAddress_ready;
	wire _networkUnits_13_io_addressOut_valid;
	wire [63:0] _networkUnits_13_io_addressOut_bits;
	wire _networkUnits_12_io_addressIn_ready;
	wire _networkUnits_12_io_peAddress_ready;
	wire _networkUnits_12_io_addressOut_valid;
	wire [63:0] _networkUnits_12_io_addressOut_bits;
	wire _networkUnits_11_io_addressIn_ready;
	wire _networkUnits_11_io_peAddress_ready;
	wire _networkUnits_11_io_addressOut_valid;
	wire [63:0] _networkUnits_11_io_addressOut_bits;
	wire _networkUnits_10_io_addressIn_ready;
	wire _networkUnits_10_io_peAddress_ready;
	wire _networkUnits_10_io_addressOut_valid;
	wire [63:0] _networkUnits_10_io_addressOut_bits;
	wire _networkUnits_9_io_addressIn_ready;
	wire _networkUnits_9_io_peAddress_ready;
	wire _networkUnits_9_io_addressOut_valid;
	wire [63:0] _networkUnits_9_io_addressOut_bits;
	wire _networkUnits_8_io_addressIn_ready;
	wire _networkUnits_8_io_peAddress_ready;
	wire _networkUnits_8_io_addressOut_valid;
	wire [63:0] _networkUnits_8_io_addressOut_bits;
	wire _networkUnits_7_io_addressIn_ready;
	wire _networkUnits_7_io_peAddress_ready;
	wire _networkUnits_7_io_addressOut_valid;
	wire [63:0] _networkUnits_7_io_addressOut_bits;
	wire _networkUnits_6_io_addressIn_ready;
	wire _networkUnits_6_io_peAddress_ready;
	wire _networkUnits_6_io_addressOut_valid;
	wire [63:0] _networkUnits_6_io_addressOut_bits;
	wire _networkUnits_5_io_addressIn_ready;
	wire _networkUnits_5_io_peAddress_ready;
	wire _networkUnits_5_io_addressOut_valid;
	wire [63:0] _networkUnits_5_io_addressOut_bits;
	wire _networkUnits_4_io_addressIn_ready;
	wire _networkUnits_4_io_peAddress_ready;
	wire _networkUnits_4_io_addressOut_valid;
	wire [63:0] _networkUnits_4_io_addressOut_bits;
	wire _networkUnits_3_io_addressIn_ready;
	wire _networkUnits_3_io_peAddress_ready;
	wire _networkUnits_3_io_addressOut_valid;
	wire [63:0] _networkUnits_3_io_addressOut_bits;
	wire _networkUnits_2_io_addressIn_ready;
	wire _networkUnits_2_io_peAddress_ready;
	wire _networkUnits_2_io_addressOut_valid;
	wire [63:0] _networkUnits_2_io_addressOut_bits;
	wire _networkUnits_1_io_addressIn_ready;
	wire _networkUnits_1_io_peAddress_ready;
	wire _networkUnits_1_io_addressOut_valid;
	wire [63:0] _networkUnits_1_io_addressOut_bits;
	wire _networkUnits_0_io_addressIn_ready;
	wire _networkUnits_0_io_peAddress_ready;
	wire _networkUnits_0_io_addressOut_valid;
	wire [63:0] _networkUnits_0_io_addressOut_bits;
	ArgumentNotifierNetworkUnit networkUnits_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_1_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_0_io_peAddress_ready),
		.io_peAddress_valid(_queues_0_io_addressOut_valid),
		.io_peAddress_bits(_queues_0_io_addressOut_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_15_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_0_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_2_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_1_io_peAddress_ready),
		.io_peAddress_valid(_queues_1_io_addressOut_valid),
		.io_peAddress_bits(_queues_1_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_1_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_3_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_2_io_peAddress_ready),
		.io_peAddress_valid(_queues_2_io_addressOut_valid),
		.io_peAddress_bits(_queues_2_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_2_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_4_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_3_io_peAddress_ready),
		.io_peAddress_valid(_queues_3_io_addressOut_valid),
		.io_peAddress_bits(_queues_3_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_3_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_5_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_4_io_peAddress_ready),
		.io_peAddress_valid(_queues_4_io_addressOut_valid),
		.io_peAddress_bits(_queues_4_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_4_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_6_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_5_io_peAddress_ready),
		.io_peAddress_valid(_queues_5_io_addressOut_valid),
		.io_peAddress_bits(_queues_5_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_5_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_7_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_6_io_peAddress_ready),
		.io_peAddress_valid(_queues_6_io_addressOut_valid),
		.io_peAddress_bits(_queues_6_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_6_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_8_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_7_io_peAddress_ready),
		.io_peAddress_valid(_queues_7_io_addressOut_valid),
		.io_peAddress_bits(_queues_7_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_7_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_9_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_8_io_peAddress_ready),
		.io_peAddress_valid(_queues_8_io_addressOut_valid),
		.io_peAddress_bits(_queues_8_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_8_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_10_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_9_io_peAddress_ready),
		.io_peAddress_valid(_queues_9_io_addressOut_valid),
		.io_peAddress_bits(_queues_9_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_9_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_11_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_10_io_peAddress_ready),
		.io_peAddress_valid(_queues_10_io_addressOut_valid),
		.io_peAddress_bits(_queues_10_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_10_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_12_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_11_io_peAddress_ready),
		.io_peAddress_valid(_queues_11_io_addressOut_valid),
		.io_peAddress_bits(_queues_11_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_11_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_13_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_12_io_peAddress_ready),
		.io_peAddress_valid(_queues_12_io_addressOut_valid),
		.io_peAddress_bits(_queues_12_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_12_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_14_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_13_io_peAddress_ready),
		.io_peAddress_valid(_queues_13_io_addressOut_valid),
		.io_peAddress_bits(_queues_13_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_13_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_15_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_14_io_peAddress_ready),
		.io_peAddress_valid(_queues_14_io_addressOut_valid),
		.io_peAddress_bits(_queues_14_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_14_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_16_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_15_io_peAddress_ready),
		.io_peAddress_valid(_queues_15_io_addressOut_valid),
		.io_peAddress_bits(_queues_15_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_15_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_17_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_16_io_peAddress_ready),
		.io_peAddress_valid(_queues_16_io_addressOut_valid),
		.io_peAddress_bits(_queues_16_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_16_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_18_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_17_io_peAddress_ready),
		.io_peAddress_valid(_queues_17_io_addressOut_valid),
		.io_peAddress_bits(_queues_17_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_17_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_19_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_18_io_peAddress_ready),
		.io_peAddress_valid(_queues_18_io_addressOut_valid),
		.io_peAddress_bits(_queues_18_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_18_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_20_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_19_io_peAddress_ready),
		.io_peAddress_valid(_queues_19_io_addressOut_valid),
		.io_peAddress_bits(_queues_19_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_19_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_21_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_20_io_peAddress_ready),
		.io_peAddress_valid(_queues_20_io_addressOut_valid),
		.io_peAddress_bits(_queues_20_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_20_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_22_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_21_io_peAddress_ready),
		.io_peAddress_valid(_queues_21_io_addressOut_valid),
		.io_peAddress_bits(_queues_21_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_21_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_23_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_22_io_peAddress_ready),
		.io_peAddress_valid(_queues_22_io_addressOut_valid),
		.io_peAddress_bits(_queues_22_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_22_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_24_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_23_io_peAddress_ready),
		.io_peAddress_valid(_queues_23_io_addressOut_valid),
		.io_peAddress_bits(_queues_23_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_23_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_25_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_24_io_peAddress_ready),
		.io_peAddress_valid(_queues_24_io_addressOut_valid),
		.io_peAddress_bits(_queues_24_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_24_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_26_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_25_io_peAddress_ready),
		.io_peAddress_valid(_queues_25_io_addressOut_valid),
		.io_peAddress_bits(_queues_25_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_25_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_27_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_26_io_peAddress_ready),
		.io_peAddress_valid(_queues_26_io_addressOut_valid),
		.io_peAddress_bits(_queues_26_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_26_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_28_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_27_io_peAddress_ready),
		.io_peAddress_valid(_queues_27_io_addressOut_valid),
		.io_peAddress_bits(_queues_27_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_27_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_29_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_28_io_peAddress_ready),
		.io_peAddress_valid(_queues_28_io_addressOut_valid),
		.io_peAddress_bits(_queues_28_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_28_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_30_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_29_io_peAddress_ready),
		.io_peAddress_valid(_queues_29_io_addressOut_valid),
		.io_peAddress_bits(_queues_29_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_29_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_31_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_30_io_peAddress_ready),
		.io_peAddress_valid(_queues_30_io_addressOut_valid),
		.io_peAddress_bits(_queues_30_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_30_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_32_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_31_io_peAddress_ready),
		.io_peAddress_valid(_queues_31_io_addressOut_valid),
		.io_peAddress_bits(_queues_31_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_31_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_33_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_32_io_peAddress_ready),
		.io_peAddress_valid(_queues_32_io_addressOut_valid),
		.io_peAddress_bits(_queues_32_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_32_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_34_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_33_io_peAddress_ready),
		.io_peAddress_valid(_queues_33_io_addressOut_valid),
		.io_peAddress_bits(_queues_33_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_33_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_35_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_34_io_peAddress_ready),
		.io_peAddress_valid(_queues_34_io_addressOut_valid),
		.io_peAddress_bits(_queues_34_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_34_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_36_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_35_io_peAddress_ready),
		.io_peAddress_valid(_queues_35_io_addressOut_valid),
		.io_peAddress_bits(_queues_35_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_35_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_37_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_36_io_peAddress_ready),
		.io_peAddress_valid(_queues_36_io_addressOut_valid),
		.io_peAddress_bits(_queues_36_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_36_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_38_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_37_io_peAddress_ready),
		.io_peAddress_valid(_queues_37_io_addressOut_valid),
		.io_peAddress_bits(_queues_37_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_37_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_39_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_38_io_peAddress_ready),
		.io_peAddress_valid(_queues_38_io_addressOut_valid),
		.io_peAddress_bits(_queues_38_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_38_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_40_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_39_io_peAddress_ready),
		.io_peAddress_valid(_queues_39_io_addressOut_valid),
		.io_peAddress_bits(_queues_39_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_39_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_41_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_40_io_peAddress_ready),
		.io_peAddress_valid(_queues_40_io_addressOut_valid),
		.io_peAddress_bits(_queues_40_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_40_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_42_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_41_io_peAddress_ready),
		.io_peAddress_valid(_queues_41_io_addressOut_valid),
		.io_peAddress_bits(_queues_41_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_41_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_43_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_42_io_peAddress_ready),
		.io_peAddress_valid(_queues_42_io_addressOut_valid),
		.io_peAddress_bits(_queues_42_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_42_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_44_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_43_io_peAddress_ready),
		.io_peAddress_valid(_queues_43_io_addressOut_valid),
		.io_peAddress_bits(_queues_43_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_43_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_45_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_44_io_peAddress_ready),
		.io_peAddress_valid(_queues_44_io_addressOut_valid),
		.io_peAddress_bits(_queues_44_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_44_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_46_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_45_io_peAddress_ready),
		.io_peAddress_valid(_queues_45_io_addressOut_valid),
		.io_peAddress_bits(_queues_45_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_45_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_47_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_46_io_peAddress_ready),
		.io_peAddress_valid(_queues_46_io_addressOut_valid),
		.io_peAddress_bits(_queues_46_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_46_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_48_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_47_io_peAddress_ready),
		.io_peAddress_valid(_queues_47_io_addressOut_valid),
		.io_peAddress_bits(_queues_47_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_47_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_49_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_48_io_peAddress_ready),
		.io_peAddress_valid(_queues_48_io_addressOut_valid),
		.io_peAddress_bits(_queues_48_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_48_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_50_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_49_io_peAddress_ready),
		.io_peAddress_valid(_queues_49_io_addressOut_valid),
		.io_peAddress_bits(_queues_49_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_49_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_51_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_50_io_peAddress_ready),
		.io_peAddress_valid(_queues_50_io_addressOut_valid),
		.io_peAddress_bits(_queues_50_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_50_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_52_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_51_io_peAddress_ready),
		.io_peAddress_valid(_queues_51_io_addressOut_valid),
		.io_peAddress_bits(_queues_51_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_51_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_53_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_52_io_peAddress_ready),
		.io_peAddress_valid(_queues_52_io_addressOut_valid),
		.io_peAddress_bits(_queues_52_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_52_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_54_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_53_io_peAddress_ready),
		.io_peAddress_valid(_queues_53_io_addressOut_valid),
		.io_peAddress_bits(_queues_53_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_53_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_55_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_54_io_peAddress_ready),
		.io_peAddress_valid(_queues_54_io_addressOut_valid),
		.io_peAddress_bits(_queues_54_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_54_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_56_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_55_io_peAddress_ready),
		.io_peAddress_valid(_queues_55_io_addressOut_valid),
		.io_peAddress_bits(_queues_55_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_55_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_57_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_56_io_peAddress_ready),
		.io_peAddress_valid(_queues_56_io_addressOut_valid),
		.io_peAddress_bits(_queues_56_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_56_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_58_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_57_io_peAddress_ready),
		.io_peAddress_valid(_queues_57_io_addressOut_valid),
		.io_peAddress_bits(_queues_57_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_57_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_59_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_58_io_peAddress_ready),
		.io_peAddress_valid(_queues_58_io_addressOut_valid),
		.io_peAddress_bits(_queues_58_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_58_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_60_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_59_io_peAddress_ready),
		.io_peAddress_valid(_queues_59_io_addressOut_valid),
		.io_peAddress_bits(_queues_59_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_59_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_61_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_60_io_peAddress_ready),
		.io_peAddress_valid(_queues_60_io_addressOut_valid),
		.io_peAddress_bits(_queues_60_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_60_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_62_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_61_io_peAddress_ready),
		.io_peAddress_valid(_queues_61_io_addressOut_valid),
		.io_peAddress_bits(_queues_61_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_61_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_63_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_63_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_62_io_peAddress_ready),
		.io_peAddress_valid(_queues_62_io_addressOut_valid),
		.io_peAddress_bits(_queues_62_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_62_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_64_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_64_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_63_io_peAddress_ready),
		.io_peAddress_valid(_queues_63_io_addressOut_valid),
		.io_peAddress_bits(_queues_63_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_63_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_63_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_64(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_64_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_65_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_65_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_64_io_peAddress_ready),
		.io_peAddress_valid(_queues_64_io_addressOut_valid),
		.io_peAddress_bits(_queues_64_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_64_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_64_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_65(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_65_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_66_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_66_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_65_io_peAddress_ready),
		.io_peAddress_valid(_queues_65_io_addressOut_valid),
		.io_peAddress_bits(_queues_65_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_64_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_65_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_65_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_66(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_66_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_67_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_67_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_66_io_peAddress_ready),
		.io_peAddress_valid(_queues_66_io_addressOut_valid),
		.io_peAddress_bits(_queues_66_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_65_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_66_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_66_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_67(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_67_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_68_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_68_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_67_io_peAddress_ready),
		.io_peAddress_valid(_queues_67_io_addressOut_valid),
		.io_peAddress_bits(_queues_67_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_66_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_67_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_67_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_68(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_68_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_69_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_69_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_68_io_peAddress_ready),
		.io_peAddress_valid(_queues_68_io_addressOut_valid),
		.io_peAddress_bits(_queues_68_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_67_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_68_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_68_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_69(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_69_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_70_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_70_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_69_io_peAddress_ready),
		.io_peAddress_valid(_queues_69_io_addressOut_valid),
		.io_peAddress_bits(_queues_69_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_68_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_69_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_69_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_70(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_70_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_71_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_71_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_70_io_peAddress_ready),
		.io_peAddress_valid(_queues_70_io_addressOut_valid),
		.io_peAddress_bits(_queues_70_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_69_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_70_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_70_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_71(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_71_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_72_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_72_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_71_io_peAddress_ready),
		.io_peAddress_valid(_queues_71_io_addressOut_valid),
		.io_peAddress_bits(_queues_71_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_70_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_71_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_71_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_72(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_72_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_73_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_73_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_72_io_peAddress_ready),
		.io_peAddress_valid(_queues_72_io_addressOut_valid),
		.io_peAddress_bits(_queues_72_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_71_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_72_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_72_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_73(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_73_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_74_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_74_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_73_io_peAddress_ready),
		.io_peAddress_valid(_queues_73_io_addressOut_valid),
		.io_peAddress_bits(_queues_73_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_72_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_73_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_73_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_74(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_74_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_75_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_75_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_74_io_peAddress_ready),
		.io_peAddress_valid(_queues_74_io_addressOut_valid),
		.io_peAddress_bits(_queues_74_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_73_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_74_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_74_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_75(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_75_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_76_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_76_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_75_io_peAddress_ready),
		.io_peAddress_valid(_queues_75_io_addressOut_valid),
		.io_peAddress_bits(_queues_75_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_74_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_75_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_75_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_76(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_76_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_77_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_77_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_76_io_peAddress_ready),
		.io_peAddress_valid(_queues_76_io_addressOut_valid),
		.io_peAddress_bits(_queues_76_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_75_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_76_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_76_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_77(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_77_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_78_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_78_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_77_io_peAddress_ready),
		.io_peAddress_valid(_queues_77_io_addressOut_valid),
		.io_peAddress_bits(_queues_77_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_76_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_77_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_77_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_78(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_78_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_79_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_79_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_78_io_peAddress_ready),
		.io_peAddress_valid(_queues_78_io_addressOut_valid),
		.io_peAddress_bits(_queues_78_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_77_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_78_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_78_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_79(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_79_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_80_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_80_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_79_io_peAddress_ready),
		.io_peAddress_valid(_queues_79_io_addressOut_valid),
		.io_peAddress_bits(_queues_79_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_78_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_79_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_79_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_80(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_80_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_81_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_81_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_80_io_peAddress_ready),
		.io_peAddress_valid(_queues_80_io_addressOut_valid),
		.io_peAddress_bits(_queues_80_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_79_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_80_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_80_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_81(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_81_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_82_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_82_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_81_io_peAddress_ready),
		.io_peAddress_valid(_queues_81_io_addressOut_valid),
		.io_peAddress_bits(_queues_81_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_80_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_81_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_81_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_82(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_82_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_83_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_83_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_82_io_peAddress_ready),
		.io_peAddress_valid(_queues_82_io_addressOut_valid),
		.io_peAddress_bits(_queues_82_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_81_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_82_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_82_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_83(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_83_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_84_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_84_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_83_io_peAddress_ready),
		.io_peAddress_valid(_queues_83_io_addressOut_valid),
		.io_peAddress_bits(_queues_83_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_82_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_83_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_83_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_84(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_84_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_85_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_85_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_84_io_peAddress_ready),
		.io_peAddress_valid(_queues_84_io_addressOut_valid),
		.io_peAddress_bits(_queues_84_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_83_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_84_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_84_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_85(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_85_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_86_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_86_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_85_io_peAddress_ready),
		.io_peAddress_valid(_queues_85_io_addressOut_valid),
		.io_peAddress_bits(_queues_85_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_84_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_85_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_85_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_86(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_86_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_87_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_87_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_86_io_peAddress_ready),
		.io_peAddress_valid(_queues_86_io_addressOut_valid),
		.io_peAddress_bits(_queues_86_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_85_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_86_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_86_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_87(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_87_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_88_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_88_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_87_io_peAddress_ready),
		.io_peAddress_valid(_queues_87_io_addressOut_valid),
		.io_peAddress_bits(_queues_87_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_86_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_87_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_87_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_88(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_88_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_89_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_89_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_88_io_peAddress_ready),
		.io_peAddress_valid(_queues_88_io_addressOut_valid),
		.io_peAddress_bits(_queues_88_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_87_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_88_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_88_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_89(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_89_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_90_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_90_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_89_io_peAddress_ready),
		.io_peAddress_valid(_queues_89_io_addressOut_valid),
		.io_peAddress_bits(_queues_89_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_88_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_89_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_89_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_90(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_90_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_91_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_91_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_90_io_peAddress_ready),
		.io_peAddress_valid(_queues_90_io_addressOut_valid),
		.io_peAddress_bits(_queues_90_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_89_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_90_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_90_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_91(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_91_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_92_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_92_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_91_io_peAddress_ready),
		.io_peAddress_valid(_queues_91_io_addressOut_valid),
		.io_peAddress_bits(_queues_91_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_90_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_91_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_91_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_92(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_92_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_93_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_93_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_92_io_peAddress_ready),
		.io_peAddress_valid(_queues_92_io_addressOut_valid),
		.io_peAddress_bits(_queues_92_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_91_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_92_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_92_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_93(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_93_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_94_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_94_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_93_io_peAddress_ready),
		.io_peAddress_valid(_queues_93_io_addressOut_valid),
		.io_peAddress_bits(_queues_93_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_92_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_93_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_93_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_94(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_94_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_95_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_95_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_94_io_peAddress_ready),
		.io_peAddress_valid(_queues_94_io_addressOut_valid),
		.io_peAddress_bits(_queues_94_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_93_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_94_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_94_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_95(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_95_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_96_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_96_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_95_io_peAddress_ready),
		.io_peAddress_valid(_queues_95_io_addressOut_valid),
		.io_peAddress_bits(_queues_95_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_94_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_95_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_95_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_96(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_96_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_97_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_97_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_96_io_peAddress_ready),
		.io_peAddress_valid(_queues_96_io_addressOut_valid),
		.io_peAddress_bits(_queues_96_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_95_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_96_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_96_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_97(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_97_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_98_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_98_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_97_io_peAddress_ready),
		.io_peAddress_valid(_queues_97_io_addressOut_valid),
		.io_peAddress_bits(_queues_97_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_96_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_97_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_97_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_98(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_98_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_99_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_99_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_98_io_peAddress_ready),
		.io_peAddress_valid(_queues_98_io_addressOut_valid),
		.io_peAddress_bits(_queues_98_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_97_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_98_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_98_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_99(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_99_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_100_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_100_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_99_io_peAddress_ready),
		.io_peAddress_valid(_queues_99_io_addressOut_valid),
		.io_peAddress_bits(_queues_99_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_98_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_99_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_99_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_100(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_100_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_101_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_101_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_100_io_peAddress_ready),
		.io_peAddress_valid(_queues_100_io_addressOut_valid),
		.io_peAddress_bits(_queues_100_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_99_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_100_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_100_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_101(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_101_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_102_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_102_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_101_io_peAddress_ready),
		.io_peAddress_valid(_queues_101_io_addressOut_valid),
		.io_peAddress_bits(_queues_101_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_100_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_101_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_101_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_102(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_102_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_103_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_103_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_102_io_peAddress_ready),
		.io_peAddress_valid(_queues_102_io_addressOut_valid),
		.io_peAddress_bits(_queues_102_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_101_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_102_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_102_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_103(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_103_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_104_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_104_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_103_io_peAddress_ready),
		.io_peAddress_valid(_queues_103_io_addressOut_valid),
		.io_peAddress_bits(_queues_103_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_102_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_103_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_103_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_104(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_104_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_105_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_105_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_104_io_peAddress_ready),
		.io_peAddress_valid(_queues_104_io_addressOut_valid),
		.io_peAddress_bits(_queues_104_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_103_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_104_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_104_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_105(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_105_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_106_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_106_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_105_io_peAddress_ready),
		.io_peAddress_valid(_queues_105_io_addressOut_valid),
		.io_peAddress_bits(_queues_105_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_104_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_105_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_105_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_106(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_106_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_107_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_107_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_106_io_peAddress_ready),
		.io_peAddress_valid(_queues_106_io_addressOut_valid),
		.io_peAddress_bits(_queues_106_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_105_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_106_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_106_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_107(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_107_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_108_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_108_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_107_io_peAddress_ready),
		.io_peAddress_valid(_queues_107_io_addressOut_valid),
		.io_peAddress_bits(_queues_107_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_106_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_107_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_107_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_108(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_108_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_109_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_109_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_108_io_peAddress_ready),
		.io_peAddress_valid(_queues_108_io_addressOut_valid),
		.io_peAddress_bits(_queues_108_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_107_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_108_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_108_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_109(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_109_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_110_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_110_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_109_io_peAddress_ready),
		.io_peAddress_valid(_queues_109_io_addressOut_valid),
		.io_peAddress_bits(_queues_109_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_108_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_109_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_109_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_110(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_110_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_111_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_111_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_110_io_peAddress_ready),
		.io_peAddress_valid(_queues_110_io_addressOut_valid),
		.io_peAddress_bits(_queues_110_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_109_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_110_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_110_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_111(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_111_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_112_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_112_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_111_io_peAddress_ready),
		.io_peAddress_valid(_queues_111_io_addressOut_valid),
		.io_peAddress_bits(_queues_111_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_110_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_111_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_111_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_112(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_112_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_113_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_113_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_112_io_peAddress_ready),
		.io_peAddress_valid(_queues_112_io_addressOut_valid),
		.io_peAddress_bits(_queues_112_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_111_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_112_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_112_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_113(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_113_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_114_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_114_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_113_io_peAddress_ready),
		.io_peAddress_valid(_queues_113_io_addressOut_valid),
		.io_peAddress_bits(_queues_113_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_112_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_113_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_113_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_114(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_114_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_115_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_115_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_114_io_peAddress_ready),
		.io_peAddress_valid(_queues_114_io_addressOut_valid),
		.io_peAddress_bits(_queues_114_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_113_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_114_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_114_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_115(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_115_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_116_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_116_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_115_io_peAddress_ready),
		.io_peAddress_valid(_queues_115_io_addressOut_valid),
		.io_peAddress_bits(_queues_115_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_114_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_115_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_115_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_116(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_116_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_117_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_117_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_116_io_peAddress_ready),
		.io_peAddress_valid(_queues_116_io_addressOut_valid),
		.io_peAddress_bits(_queues_116_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_115_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_116_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_116_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_117(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_117_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_118_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_118_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_117_io_peAddress_ready),
		.io_peAddress_valid(_queues_117_io_addressOut_valid),
		.io_peAddress_bits(_queues_117_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_116_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_117_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_117_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_118(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_118_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_119_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_119_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_118_io_peAddress_ready),
		.io_peAddress_valid(_queues_118_io_addressOut_valid),
		.io_peAddress_bits(_queues_118_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_117_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_118_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_118_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_119(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_119_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_120_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_120_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_119_io_peAddress_ready),
		.io_peAddress_valid(_queues_119_io_addressOut_valid),
		.io_peAddress_bits(_queues_119_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_118_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_119_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_119_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_120(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_120_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_121_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_121_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_120_io_peAddress_ready),
		.io_peAddress_valid(_queues_120_io_addressOut_valid),
		.io_peAddress_bits(_queues_120_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_119_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_120_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_120_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_121(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_121_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_122_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_122_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_121_io_peAddress_ready),
		.io_peAddress_valid(_queues_121_io_addressOut_valid),
		.io_peAddress_bits(_queues_121_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_120_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_121_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_121_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_122(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_122_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_123_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_123_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_122_io_peAddress_ready),
		.io_peAddress_valid(_queues_122_io_addressOut_valid),
		.io_peAddress_bits(_queues_122_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_121_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_122_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_122_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_123(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_123_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_124_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_124_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_123_io_peAddress_ready),
		.io_peAddress_valid(_queues_123_io_addressOut_valid),
		.io_peAddress_bits(_queues_123_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_122_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_123_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_123_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_124(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_124_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_125_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_125_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_124_io_peAddress_ready),
		.io_peAddress_valid(_queues_124_io_addressOut_valid),
		.io_peAddress_bits(_queues_124_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_123_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_124_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_124_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_125(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_125_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_126_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_126_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_125_io_peAddress_ready),
		.io_peAddress_valid(_queues_125_io_addressOut_valid),
		.io_peAddress_bits(_queues_125_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_124_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_125_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_125_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_126(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_126_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_127_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_127_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_126_io_peAddress_ready),
		.io_peAddress_valid(_queues_126_io_addressOut_valid),
		.io_peAddress_bits(_queues_126_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_125_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_126_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_126_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_127(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(),
		.io_addressIn_valid(1'h0),
		.io_addressIn_bits(64'h0000000000000000),
		.io_peAddress_ready(_networkUnits_127_io_peAddress_ready),
		.io_peAddress_valid(_queues_127_io_addressOut_valid),
		.io_peAddress_bits(_queues_127_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_126_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_127_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_127_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit ArgumentNotifierServerNetworkUnit(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_0_ready),
		.io_vasAddressOut_valid(io_connVAS_0_valid),
		.io_vasAddressOut_bits(io_connVAS_0_bits)
	);
	ArgumentNotifierServerNetworkUnit_1 ArgumentNotifierServerNetworkUnit_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_1_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_1_ready),
		.io_vasAddressOut_valid(io_connVAS_1_valid),
		.io_vasAddressOut_bits(io_connVAS_1_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_2 ArgumentNotifierServerNetworkUnit_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_2_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_2_ready),
		.io_vasAddressOut_valid(io_connVAS_2_valid),
		.io_vasAddressOut_bits(io_connVAS_2_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_1_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_3 ArgumentNotifierServerNetworkUnit_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_3_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_3_ready),
		.io_vasAddressOut_valid(io_connVAS_3_valid),
		.io_vasAddressOut_bits(io_connVAS_3_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_2_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_4 ArgumentNotifierServerNetworkUnit_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_4_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_4_ready),
		.io_vasAddressOut_valid(io_connVAS_4_valid),
		.io_vasAddressOut_bits(io_connVAS_4_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_3_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_5 ArgumentNotifierServerNetworkUnit_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_5_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_5_ready),
		.io_vasAddressOut_valid(io_connVAS_5_valid),
		.io_vasAddressOut_bits(io_connVAS_5_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_4_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_6 ArgumentNotifierServerNetworkUnit_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_6_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_6_ready),
		.io_vasAddressOut_valid(io_connVAS_6_valid),
		.io_vasAddressOut_bits(io_connVAS_6_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_5_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_7 ArgumentNotifierServerNetworkUnit_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_7_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_7_ready),
		.io_vasAddressOut_valid(io_connVAS_7_valid),
		.io_vasAddressOut_bits(io_connVAS_7_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_6_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_8 ArgumentNotifierServerNetworkUnit_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_8_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_8_ready),
		.io_vasAddressOut_valid(io_connVAS_8_valid),
		.io_vasAddressOut_bits(io_connVAS_8_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_7_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_9 ArgumentNotifierServerNetworkUnit_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_9_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_9_ready),
		.io_vasAddressOut_valid(io_connVAS_9_valid),
		.io_vasAddressOut_bits(io_connVAS_9_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_8_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_10 ArgumentNotifierServerNetworkUnit_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_10_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_10_ready),
		.io_vasAddressOut_valid(io_connVAS_10_valid),
		.io_vasAddressOut_bits(io_connVAS_10_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_9_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_11 ArgumentNotifierServerNetworkUnit_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_11_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_11_ready),
		.io_vasAddressOut_valid(io_connVAS_11_valid),
		.io_vasAddressOut_bits(io_connVAS_11_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_10_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_12 ArgumentNotifierServerNetworkUnit_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_12_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_12_ready),
		.io_vasAddressOut_valid(io_connVAS_12_valid),
		.io_vasAddressOut_bits(io_connVAS_12_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_11_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_13 ArgumentNotifierServerNetworkUnit_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_13_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_13_ready),
		.io_vasAddressOut_valid(io_connVAS_13_valid),
		.io_vasAddressOut_bits(io_connVAS_13_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_12_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_14 ArgumentNotifierServerNetworkUnit_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_14_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_14_ready),
		.io_vasAddressOut_valid(io_connVAS_14_valid),
		.io_vasAddressOut_bits(io_connVAS_14_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_13_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_15 ArgumentNotifierServerNetworkUnit_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_0_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_15_ready),
		.io_vasAddressOut_valid(io_connVAS_15_valid),
		.io_vasAddressOut_bits(io_connVAS_15_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_14_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_0_ready),
		.io_addressIn_valid(io_connPE_0_valid),
		.io_addressIn_bits(io_connPE_0_bits),
		.io_addressOut_ready(_networkUnits_0_io_peAddress_ready),
		.io_addressOut_valid(_queues_0_io_addressOut_valid),
		.io_addressOut_bits(_queues_0_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_1_ready),
		.io_addressIn_valid(io_connPE_1_valid),
		.io_addressIn_bits(io_connPE_1_bits),
		.io_addressOut_ready(_networkUnits_1_io_peAddress_ready),
		.io_addressOut_valid(_queues_1_io_addressOut_valid),
		.io_addressOut_bits(_queues_1_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_2_ready),
		.io_addressIn_valid(io_connPE_2_valid),
		.io_addressIn_bits(io_connPE_2_bits),
		.io_addressOut_ready(_networkUnits_2_io_peAddress_ready),
		.io_addressOut_valid(_queues_2_io_addressOut_valid),
		.io_addressOut_bits(_queues_2_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_3_ready),
		.io_addressIn_valid(io_connPE_3_valid),
		.io_addressIn_bits(io_connPE_3_bits),
		.io_addressOut_ready(_networkUnits_3_io_peAddress_ready),
		.io_addressOut_valid(_queues_3_io_addressOut_valid),
		.io_addressOut_bits(_queues_3_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_4_ready),
		.io_addressIn_valid(io_connPE_4_valid),
		.io_addressIn_bits(io_connPE_4_bits),
		.io_addressOut_ready(_networkUnits_4_io_peAddress_ready),
		.io_addressOut_valid(_queues_4_io_addressOut_valid),
		.io_addressOut_bits(_queues_4_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_5_ready),
		.io_addressIn_valid(io_connPE_5_valid),
		.io_addressIn_bits(io_connPE_5_bits),
		.io_addressOut_ready(_networkUnits_5_io_peAddress_ready),
		.io_addressOut_valid(_queues_5_io_addressOut_valid),
		.io_addressOut_bits(_queues_5_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_6_ready),
		.io_addressIn_valid(io_connPE_6_valid),
		.io_addressIn_bits(io_connPE_6_bits),
		.io_addressOut_ready(_networkUnits_6_io_peAddress_ready),
		.io_addressOut_valid(_queues_6_io_addressOut_valid),
		.io_addressOut_bits(_queues_6_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_7_ready),
		.io_addressIn_valid(io_connPE_7_valid),
		.io_addressIn_bits(io_connPE_7_bits),
		.io_addressOut_ready(_networkUnits_7_io_peAddress_ready),
		.io_addressOut_valid(_queues_7_io_addressOut_valid),
		.io_addressOut_bits(_queues_7_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_8_ready),
		.io_addressIn_valid(io_connPE_8_valid),
		.io_addressIn_bits(io_connPE_8_bits),
		.io_addressOut_ready(_networkUnits_8_io_peAddress_ready),
		.io_addressOut_valid(_queues_8_io_addressOut_valid),
		.io_addressOut_bits(_queues_8_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_9_ready),
		.io_addressIn_valid(io_connPE_9_valid),
		.io_addressIn_bits(io_connPE_9_bits),
		.io_addressOut_ready(_networkUnits_9_io_peAddress_ready),
		.io_addressOut_valid(_queues_9_io_addressOut_valid),
		.io_addressOut_bits(_queues_9_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_10_ready),
		.io_addressIn_valid(io_connPE_10_valid),
		.io_addressIn_bits(io_connPE_10_bits),
		.io_addressOut_ready(_networkUnits_10_io_peAddress_ready),
		.io_addressOut_valid(_queues_10_io_addressOut_valid),
		.io_addressOut_bits(_queues_10_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_11_ready),
		.io_addressIn_valid(io_connPE_11_valid),
		.io_addressIn_bits(io_connPE_11_bits),
		.io_addressOut_ready(_networkUnits_11_io_peAddress_ready),
		.io_addressOut_valid(_queues_11_io_addressOut_valid),
		.io_addressOut_bits(_queues_11_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_12_ready),
		.io_addressIn_valid(io_connPE_12_valid),
		.io_addressIn_bits(io_connPE_12_bits),
		.io_addressOut_ready(_networkUnits_12_io_peAddress_ready),
		.io_addressOut_valid(_queues_12_io_addressOut_valid),
		.io_addressOut_bits(_queues_12_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_13_ready),
		.io_addressIn_valid(io_connPE_13_valid),
		.io_addressIn_bits(io_connPE_13_bits),
		.io_addressOut_ready(_networkUnits_13_io_peAddress_ready),
		.io_addressOut_valid(_queues_13_io_addressOut_valid),
		.io_addressOut_bits(_queues_13_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_14_ready),
		.io_addressIn_valid(io_connPE_14_valid),
		.io_addressIn_bits(io_connPE_14_bits),
		.io_addressOut_ready(_networkUnits_14_io_peAddress_ready),
		.io_addressOut_valid(_queues_14_io_addressOut_valid),
		.io_addressOut_bits(_queues_14_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_15_ready),
		.io_addressIn_valid(io_connPE_15_valid),
		.io_addressIn_bits(io_connPE_15_bits),
		.io_addressOut_ready(_networkUnits_15_io_peAddress_ready),
		.io_addressOut_valid(_queues_15_io_addressOut_valid),
		.io_addressOut_bits(_queues_15_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_16_ready),
		.io_addressIn_valid(io_connPE_16_valid),
		.io_addressIn_bits(io_connPE_16_bits),
		.io_addressOut_ready(_networkUnits_16_io_peAddress_ready),
		.io_addressOut_valid(_queues_16_io_addressOut_valid),
		.io_addressOut_bits(_queues_16_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_17_ready),
		.io_addressIn_valid(io_connPE_17_valid),
		.io_addressIn_bits(io_connPE_17_bits),
		.io_addressOut_ready(_networkUnits_17_io_peAddress_ready),
		.io_addressOut_valid(_queues_17_io_addressOut_valid),
		.io_addressOut_bits(_queues_17_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_18_ready),
		.io_addressIn_valid(io_connPE_18_valid),
		.io_addressIn_bits(io_connPE_18_bits),
		.io_addressOut_ready(_networkUnits_18_io_peAddress_ready),
		.io_addressOut_valid(_queues_18_io_addressOut_valid),
		.io_addressOut_bits(_queues_18_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_19_ready),
		.io_addressIn_valid(io_connPE_19_valid),
		.io_addressIn_bits(io_connPE_19_bits),
		.io_addressOut_ready(_networkUnits_19_io_peAddress_ready),
		.io_addressOut_valid(_queues_19_io_addressOut_valid),
		.io_addressOut_bits(_queues_19_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_20_ready),
		.io_addressIn_valid(io_connPE_20_valid),
		.io_addressIn_bits(io_connPE_20_bits),
		.io_addressOut_ready(_networkUnits_20_io_peAddress_ready),
		.io_addressOut_valid(_queues_20_io_addressOut_valid),
		.io_addressOut_bits(_queues_20_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_21_ready),
		.io_addressIn_valid(io_connPE_21_valid),
		.io_addressIn_bits(io_connPE_21_bits),
		.io_addressOut_ready(_networkUnits_21_io_peAddress_ready),
		.io_addressOut_valid(_queues_21_io_addressOut_valid),
		.io_addressOut_bits(_queues_21_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_22_ready),
		.io_addressIn_valid(io_connPE_22_valid),
		.io_addressIn_bits(io_connPE_22_bits),
		.io_addressOut_ready(_networkUnits_22_io_peAddress_ready),
		.io_addressOut_valid(_queues_22_io_addressOut_valid),
		.io_addressOut_bits(_queues_22_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_23_ready),
		.io_addressIn_valid(io_connPE_23_valid),
		.io_addressIn_bits(io_connPE_23_bits),
		.io_addressOut_ready(_networkUnits_23_io_peAddress_ready),
		.io_addressOut_valid(_queues_23_io_addressOut_valid),
		.io_addressOut_bits(_queues_23_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_24_ready),
		.io_addressIn_valid(io_connPE_24_valid),
		.io_addressIn_bits(io_connPE_24_bits),
		.io_addressOut_ready(_networkUnits_24_io_peAddress_ready),
		.io_addressOut_valid(_queues_24_io_addressOut_valid),
		.io_addressOut_bits(_queues_24_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_25_ready),
		.io_addressIn_valid(io_connPE_25_valid),
		.io_addressIn_bits(io_connPE_25_bits),
		.io_addressOut_ready(_networkUnits_25_io_peAddress_ready),
		.io_addressOut_valid(_queues_25_io_addressOut_valid),
		.io_addressOut_bits(_queues_25_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_26_ready),
		.io_addressIn_valid(io_connPE_26_valid),
		.io_addressIn_bits(io_connPE_26_bits),
		.io_addressOut_ready(_networkUnits_26_io_peAddress_ready),
		.io_addressOut_valid(_queues_26_io_addressOut_valid),
		.io_addressOut_bits(_queues_26_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_27_ready),
		.io_addressIn_valid(io_connPE_27_valid),
		.io_addressIn_bits(io_connPE_27_bits),
		.io_addressOut_ready(_networkUnits_27_io_peAddress_ready),
		.io_addressOut_valid(_queues_27_io_addressOut_valid),
		.io_addressOut_bits(_queues_27_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_28_ready),
		.io_addressIn_valid(io_connPE_28_valid),
		.io_addressIn_bits(io_connPE_28_bits),
		.io_addressOut_ready(_networkUnits_28_io_peAddress_ready),
		.io_addressOut_valid(_queues_28_io_addressOut_valid),
		.io_addressOut_bits(_queues_28_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_29_ready),
		.io_addressIn_valid(io_connPE_29_valid),
		.io_addressIn_bits(io_connPE_29_bits),
		.io_addressOut_ready(_networkUnits_29_io_peAddress_ready),
		.io_addressOut_valid(_queues_29_io_addressOut_valid),
		.io_addressOut_bits(_queues_29_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_30_ready),
		.io_addressIn_valid(io_connPE_30_valid),
		.io_addressIn_bits(io_connPE_30_bits),
		.io_addressOut_ready(_networkUnits_30_io_peAddress_ready),
		.io_addressOut_valid(_queues_30_io_addressOut_valid),
		.io_addressOut_bits(_queues_30_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_31_ready),
		.io_addressIn_valid(io_connPE_31_valid),
		.io_addressIn_bits(io_connPE_31_bits),
		.io_addressOut_ready(_networkUnits_31_io_peAddress_ready),
		.io_addressOut_valid(_queues_31_io_addressOut_valid),
		.io_addressOut_bits(_queues_31_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_32_ready),
		.io_addressIn_valid(io_connPE_32_valid),
		.io_addressIn_bits(io_connPE_32_bits),
		.io_addressOut_ready(_networkUnits_32_io_peAddress_ready),
		.io_addressOut_valid(_queues_32_io_addressOut_valid),
		.io_addressOut_bits(_queues_32_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_33_ready),
		.io_addressIn_valid(io_connPE_33_valid),
		.io_addressIn_bits(io_connPE_33_bits),
		.io_addressOut_ready(_networkUnits_33_io_peAddress_ready),
		.io_addressOut_valid(_queues_33_io_addressOut_valid),
		.io_addressOut_bits(_queues_33_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_34_ready),
		.io_addressIn_valid(io_connPE_34_valid),
		.io_addressIn_bits(io_connPE_34_bits),
		.io_addressOut_ready(_networkUnits_34_io_peAddress_ready),
		.io_addressOut_valid(_queues_34_io_addressOut_valid),
		.io_addressOut_bits(_queues_34_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_35_ready),
		.io_addressIn_valid(io_connPE_35_valid),
		.io_addressIn_bits(io_connPE_35_bits),
		.io_addressOut_ready(_networkUnits_35_io_peAddress_ready),
		.io_addressOut_valid(_queues_35_io_addressOut_valid),
		.io_addressOut_bits(_queues_35_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_36_ready),
		.io_addressIn_valid(io_connPE_36_valid),
		.io_addressIn_bits(io_connPE_36_bits),
		.io_addressOut_ready(_networkUnits_36_io_peAddress_ready),
		.io_addressOut_valid(_queues_36_io_addressOut_valid),
		.io_addressOut_bits(_queues_36_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_37_ready),
		.io_addressIn_valid(io_connPE_37_valid),
		.io_addressIn_bits(io_connPE_37_bits),
		.io_addressOut_ready(_networkUnits_37_io_peAddress_ready),
		.io_addressOut_valid(_queues_37_io_addressOut_valid),
		.io_addressOut_bits(_queues_37_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_38_ready),
		.io_addressIn_valid(io_connPE_38_valid),
		.io_addressIn_bits(io_connPE_38_bits),
		.io_addressOut_ready(_networkUnits_38_io_peAddress_ready),
		.io_addressOut_valid(_queues_38_io_addressOut_valid),
		.io_addressOut_bits(_queues_38_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_39_ready),
		.io_addressIn_valid(io_connPE_39_valid),
		.io_addressIn_bits(io_connPE_39_bits),
		.io_addressOut_ready(_networkUnits_39_io_peAddress_ready),
		.io_addressOut_valid(_queues_39_io_addressOut_valid),
		.io_addressOut_bits(_queues_39_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_40_ready),
		.io_addressIn_valid(io_connPE_40_valid),
		.io_addressIn_bits(io_connPE_40_bits),
		.io_addressOut_ready(_networkUnits_40_io_peAddress_ready),
		.io_addressOut_valid(_queues_40_io_addressOut_valid),
		.io_addressOut_bits(_queues_40_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_41_ready),
		.io_addressIn_valid(io_connPE_41_valid),
		.io_addressIn_bits(io_connPE_41_bits),
		.io_addressOut_ready(_networkUnits_41_io_peAddress_ready),
		.io_addressOut_valid(_queues_41_io_addressOut_valid),
		.io_addressOut_bits(_queues_41_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_42_ready),
		.io_addressIn_valid(io_connPE_42_valid),
		.io_addressIn_bits(io_connPE_42_bits),
		.io_addressOut_ready(_networkUnits_42_io_peAddress_ready),
		.io_addressOut_valid(_queues_42_io_addressOut_valid),
		.io_addressOut_bits(_queues_42_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_43_ready),
		.io_addressIn_valid(io_connPE_43_valid),
		.io_addressIn_bits(io_connPE_43_bits),
		.io_addressOut_ready(_networkUnits_43_io_peAddress_ready),
		.io_addressOut_valid(_queues_43_io_addressOut_valid),
		.io_addressOut_bits(_queues_43_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_44_ready),
		.io_addressIn_valid(io_connPE_44_valid),
		.io_addressIn_bits(io_connPE_44_bits),
		.io_addressOut_ready(_networkUnits_44_io_peAddress_ready),
		.io_addressOut_valid(_queues_44_io_addressOut_valid),
		.io_addressOut_bits(_queues_44_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_45_ready),
		.io_addressIn_valid(io_connPE_45_valid),
		.io_addressIn_bits(io_connPE_45_bits),
		.io_addressOut_ready(_networkUnits_45_io_peAddress_ready),
		.io_addressOut_valid(_queues_45_io_addressOut_valid),
		.io_addressOut_bits(_queues_45_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_46_ready),
		.io_addressIn_valid(io_connPE_46_valid),
		.io_addressIn_bits(io_connPE_46_bits),
		.io_addressOut_ready(_networkUnits_46_io_peAddress_ready),
		.io_addressOut_valid(_queues_46_io_addressOut_valid),
		.io_addressOut_bits(_queues_46_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_47_ready),
		.io_addressIn_valid(io_connPE_47_valid),
		.io_addressIn_bits(io_connPE_47_bits),
		.io_addressOut_ready(_networkUnits_47_io_peAddress_ready),
		.io_addressOut_valid(_queues_47_io_addressOut_valid),
		.io_addressOut_bits(_queues_47_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_48_ready),
		.io_addressIn_valid(io_connPE_48_valid),
		.io_addressIn_bits(io_connPE_48_bits),
		.io_addressOut_ready(_networkUnits_48_io_peAddress_ready),
		.io_addressOut_valid(_queues_48_io_addressOut_valid),
		.io_addressOut_bits(_queues_48_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_49_ready),
		.io_addressIn_valid(io_connPE_49_valid),
		.io_addressIn_bits(io_connPE_49_bits),
		.io_addressOut_ready(_networkUnits_49_io_peAddress_ready),
		.io_addressOut_valid(_queues_49_io_addressOut_valid),
		.io_addressOut_bits(_queues_49_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_50_ready),
		.io_addressIn_valid(io_connPE_50_valid),
		.io_addressIn_bits(io_connPE_50_bits),
		.io_addressOut_ready(_networkUnits_50_io_peAddress_ready),
		.io_addressOut_valid(_queues_50_io_addressOut_valid),
		.io_addressOut_bits(_queues_50_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_51_ready),
		.io_addressIn_valid(io_connPE_51_valid),
		.io_addressIn_bits(io_connPE_51_bits),
		.io_addressOut_ready(_networkUnits_51_io_peAddress_ready),
		.io_addressOut_valid(_queues_51_io_addressOut_valid),
		.io_addressOut_bits(_queues_51_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_52_ready),
		.io_addressIn_valid(io_connPE_52_valid),
		.io_addressIn_bits(io_connPE_52_bits),
		.io_addressOut_ready(_networkUnits_52_io_peAddress_ready),
		.io_addressOut_valid(_queues_52_io_addressOut_valid),
		.io_addressOut_bits(_queues_52_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_53_ready),
		.io_addressIn_valid(io_connPE_53_valid),
		.io_addressIn_bits(io_connPE_53_bits),
		.io_addressOut_ready(_networkUnits_53_io_peAddress_ready),
		.io_addressOut_valid(_queues_53_io_addressOut_valid),
		.io_addressOut_bits(_queues_53_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_54_ready),
		.io_addressIn_valid(io_connPE_54_valid),
		.io_addressIn_bits(io_connPE_54_bits),
		.io_addressOut_ready(_networkUnits_54_io_peAddress_ready),
		.io_addressOut_valid(_queues_54_io_addressOut_valid),
		.io_addressOut_bits(_queues_54_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_55_ready),
		.io_addressIn_valid(io_connPE_55_valid),
		.io_addressIn_bits(io_connPE_55_bits),
		.io_addressOut_ready(_networkUnits_55_io_peAddress_ready),
		.io_addressOut_valid(_queues_55_io_addressOut_valid),
		.io_addressOut_bits(_queues_55_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_56_ready),
		.io_addressIn_valid(io_connPE_56_valid),
		.io_addressIn_bits(io_connPE_56_bits),
		.io_addressOut_ready(_networkUnits_56_io_peAddress_ready),
		.io_addressOut_valid(_queues_56_io_addressOut_valid),
		.io_addressOut_bits(_queues_56_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_57_ready),
		.io_addressIn_valid(io_connPE_57_valid),
		.io_addressIn_bits(io_connPE_57_bits),
		.io_addressOut_ready(_networkUnits_57_io_peAddress_ready),
		.io_addressOut_valid(_queues_57_io_addressOut_valid),
		.io_addressOut_bits(_queues_57_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_58_ready),
		.io_addressIn_valid(io_connPE_58_valid),
		.io_addressIn_bits(io_connPE_58_bits),
		.io_addressOut_ready(_networkUnits_58_io_peAddress_ready),
		.io_addressOut_valid(_queues_58_io_addressOut_valid),
		.io_addressOut_bits(_queues_58_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_59_ready),
		.io_addressIn_valid(io_connPE_59_valid),
		.io_addressIn_bits(io_connPE_59_bits),
		.io_addressOut_ready(_networkUnits_59_io_peAddress_ready),
		.io_addressOut_valid(_queues_59_io_addressOut_valid),
		.io_addressOut_bits(_queues_59_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_60_ready),
		.io_addressIn_valid(io_connPE_60_valid),
		.io_addressIn_bits(io_connPE_60_bits),
		.io_addressOut_ready(_networkUnits_60_io_peAddress_ready),
		.io_addressOut_valid(_queues_60_io_addressOut_valid),
		.io_addressOut_bits(_queues_60_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_61_ready),
		.io_addressIn_valid(io_connPE_61_valid),
		.io_addressIn_bits(io_connPE_61_bits),
		.io_addressOut_ready(_networkUnits_61_io_peAddress_ready),
		.io_addressOut_valid(_queues_61_io_addressOut_valid),
		.io_addressOut_bits(_queues_61_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_62_ready),
		.io_addressIn_valid(io_connPE_62_valid),
		.io_addressIn_bits(io_connPE_62_bits),
		.io_addressOut_ready(_networkUnits_62_io_peAddress_ready),
		.io_addressOut_valid(_queues_62_io_addressOut_valid),
		.io_addressOut_bits(_queues_62_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_63_ready),
		.io_addressIn_valid(io_connPE_63_valid),
		.io_addressIn_bits(io_connPE_63_bits),
		.io_addressOut_ready(_networkUnits_63_io_peAddress_ready),
		.io_addressOut_valid(_queues_63_io_addressOut_valid),
		.io_addressOut_bits(_queues_63_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_64(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_64_ready),
		.io_addressIn_valid(io_connPE_64_valid),
		.io_addressIn_bits(io_connPE_64_bits),
		.io_addressOut_ready(_networkUnits_64_io_peAddress_ready),
		.io_addressOut_valid(_queues_64_io_addressOut_valid),
		.io_addressOut_bits(_queues_64_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_65(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_65_ready),
		.io_addressIn_valid(io_connPE_65_valid),
		.io_addressIn_bits(io_connPE_65_bits),
		.io_addressOut_ready(_networkUnits_65_io_peAddress_ready),
		.io_addressOut_valid(_queues_65_io_addressOut_valid),
		.io_addressOut_bits(_queues_65_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_66(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_66_ready),
		.io_addressIn_valid(io_connPE_66_valid),
		.io_addressIn_bits(io_connPE_66_bits),
		.io_addressOut_ready(_networkUnits_66_io_peAddress_ready),
		.io_addressOut_valid(_queues_66_io_addressOut_valid),
		.io_addressOut_bits(_queues_66_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_67(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_67_ready),
		.io_addressIn_valid(io_connPE_67_valid),
		.io_addressIn_bits(io_connPE_67_bits),
		.io_addressOut_ready(_networkUnits_67_io_peAddress_ready),
		.io_addressOut_valid(_queues_67_io_addressOut_valid),
		.io_addressOut_bits(_queues_67_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_68(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_68_ready),
		.io_addressIn_valid(io_connPE_68_valid),
		.io_addressIn_bits(io_connPE_68_bits),
		.io_addressOut_ready(_networkUnits_68_io_peAddress_ready),
		.io_addressOut_valid(_queues_68_io_addressOut_valid),
		.io_addressOut_bits(_queues_68_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_69(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_69_ready),
		.io_addressIn_valid(io_connPE_69_valid),
		.io_addressIn_bits(io_connPE_69_bits),
		.io_addressOut_ready(_networkUnits_69_io_peAddress_ready),
		.io_addressOut_valid(_queues_69_io_addressOut_valid),
		.io_addressOut_bits(_queues_69_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_70(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_70_ready),
		.io_addressIn_valid(io_connPE_70_valid),
		.io_addressIn_bits(io_connPE_70_bits),
		.io_addressOut_ready(_networkUnits_70_io_peAddress_ready),
		.io_addressOut_valid(_queues_70_io_addressOut_valid),
		.io_addressOut_bits(_queues_70_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_71(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_71_ready),
		.io_addressIn_valid(io_connPE_71_valid),
		.io_addressIn_bits(io_connPE_71_bits),
		.io_addressOut_ready(_networkUnits_71_io_peAddress_ready),
		.io_addressOut_valid(_queues_71_io_addressOut_valid),
		.io_addressOut_bits(_queues_71_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_72(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_72_ready),
		.io_addressIn_valid(io_connPE_72_valid),
		.io_addressIn_bits(io_connPE_72_bits),
		.io_addressOut_ready(_networkUnits_72_io_peAddress_ready),
		.io_addressOut_valid(_queues_72_io_addressOut_valid),
		.io_addressOut_bits(_queues_72_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_73(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_73_ready),
		.io_addressIn_valid(io_connPE_73_valid),
		.io_addressIn_bits(io_connPE_73_bits),
		.io_addressOut_ready(_networkUnits_73_io_peAddress_ready),
		.io_addressOut_valid(_queues_73_io_addressOut_valid),
		.io_addressOut_bits(_queues_73_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_74(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_74_ready),
		.io_addressIn_valid(io_connPE_74_valid),
		.io_addressIn_bits(io_connPE_74_bits),
		.io_addressOut_ready(_networkUnits_74_io_peAddress_ready),
		.io_addressOut_valid(_queues_74_io_addressOut_valid),
		.io_addressOut_bits(_queues_74_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_75(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_75_ready),
		.io_addressIn_valid(io_connPE_75_valid),
		.io_addressIn_bits(io_connPE_75_bits),
		.io_addressOut_ready(_networkUnits_75_io_peAddress_ready),
		.io_addressOut_valid(_queues_75_io_addressOut_valid),
		.io_addressOut_bits(_queues_75_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_76(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_76_ready),
		.io_addressIn_valid(io_connPE_76_valid),
		.io_addressIn_bits(io_connPE_76_bits),
		.io_addressOut_ready(_networkUnits_76_io_peAddress_ready),
		.io_addressOut_valid(_queues_76_io_addressOut_valid),
		.io_addressOut_bits(_queues_76_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_77(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_77_ready),
		.io_addressIn_valid(io_connPE_77_valid),
		.io_addressIn_bits(io_connPE_77_bits),
		.io_addressOut_ready(_networkUnits_77_io_peAddress_ready),
		.io_addressOut_valid(_queues_77_io_addressOut_valid),
		.io_addressOut_bits(_queues_77_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_78(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_78_ready),
		.io_addressIn_valid(io_connPE_78_valid),
		.io_addressIn_bits(io_connPE_78_bits),
		.io_addressOut_ready(_networkUnits_78_io_peAddress_ready),
		.io_addressOut_valid(_queues_78_io_addressOut_valid),
		.io_addressOut_bits(_queues_78_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_79(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_79_ready),
		.io_addressIn_valid(io_connPE_79_valid),
		.io_addressIn_bits(io_connPE_79_bits),
		.io_addressOut_ready(_networkUnits_79_io_peAddress_ready),
		.io_addressOut_valid(_queues_79_io_addressOut_valid),
		.io_addressOut_bits(_queues_79_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_80(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_80_ready),
		.io_addressIn_valid(io_connPE_80_valid),
		.io_addressIn_bits(io_connPE_80_bits),
		.io_addressOut_ready(_networkUnits_80_io_peAddress_ready),
		.io_addressOut_valid(_queues_80_io_addressOut_valid),
		.io_addressOut_bits(_queues_80_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_81(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_81_ready),
		.io_addressIn_valid(io_connPE_81_valid),
		.io_addressIn_bits(io_connPE_81_bits),
		.io_addressOut_ready(_networkUnits_81_io_peAddress_ready),
		.io_addressOut_valid(_queues_81_io_addressOut_valid),
		.io_addressOut_bits(_queues_81_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_82(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_82_ready),
		.io_addressIn_valid(io_connPE_82_valid),
		.io_addressIn_bits(io_connPE_82_bits),
		.io_addressOut_ready(_networkUnits_82_io_peAddress_ready),
		.io_addressOut_valid(_queues_82_io_addressOut_valid),
		.io_addressOut_bits(_queues_82_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_83(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_83_ready),
		.io_addressIn_valid(io_connPE_83_valid),
		.io_addressIn_bits(io_connPE_83_bits),
		.io_addressOut_ready(_networkUnits_83_io_peAddress_ready),
		.io_addressOut_valid(_queues_83_io_addressOut_valid),
		.io_addressOut_bits(_queues_83_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_84(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_84_ready),
		.io_addressIn_valid(io_connPE_84_valid),
		.io_addressIn_bits(io_connPE_84_bits),
		.io_addressOut_ready(_networkUnits_84_io_peAddress_ready),
		.io_addressOut_valid(_queues_84_io_addressOut_valid),
		.io_addressOut_bits(_queues_84_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_85(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_85_ready),
		.io_addressIn_valid(io_connPE_85_valid),
		.io_addressIn_bits(io_connPE_85_bits),
		.io_addressOut_ready(_networkUnits_85_io_peAddress_ready),
		.io_addressOut_valid(_queues_85_io_addressOut_valid),
		.io_addressOut_bits(_queues_85_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_86(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_86_ready),
		.io_addressIn_valid(io_connPE_86_valid),
		.io_addressIn_bits(io_connPE_86_bits),
		.io_addressOut_ready(_networkUnits_86_io_peAddress_ready),
		.io_addressOut_valid(_queues_86_io_addressOut_valid),
		.io_addressOut_bits(_queues_86_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_87(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_87_ready),
		.io_addressIn_valid(io_connPE_87_valid),
		.io_addressIn_bits(io_connPE_87_bits),
		.io_addressOut_ready(_networkUnits_87_io_peAddress_ready),
		.io_addressOut_valid(_queues_87_io_addressOut_valid),
		.io_addressOut_bits(_queues_87_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_88(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_88_ready),
		.io_addressIn_valid(io_connPE_88_valid),
		.io_addressIn_bits(io_connPE_88_bits),
		.io_addressOut_ready(_networkUnits_88_io_peAddress_ready),
		.io_addressOut_valid(_queues_88_io_addressOut_valid),
		.io_addressOut_bits(_queues_88_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_89(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_89_ready),
		.io_addressIn_valid(io_connPE_89_valid),
		.io_addressIn_bits(io_connPE_89_bits),
		.io_addressOut_ready(_networkUnits_89_io_peAddress_ready),
		.io_addressOut_valid(_queues_89_io_addressOut_valid),
		.io_addressOut_bits(_queues_89_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_90(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_90_ready),
		.io_addressIn_valid(io_connPE_90_valid),
		.io_addressIn_bits(io_connPE_90_bits),
		.io_addressOut_ready(_networkUnits_90_io_peAddress_ready),
		.io_addressOut_valid(_queues_90_io_addressOut_valid),
		.io_addressOut_bits(_queues_90_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_91(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_91_ready),
		.io_addressIn_valid(io_connPE_91_valid),
		.io_addressIn_bits(io_connPE_91_bits),
		.io_addressOut_ready(_networkUnits_91_io_peAddress_ready),
		.io_addressOut_valid(_queues_91_io_addressOut_valid),
		.io_addressOut_bits(_queues_91_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_92(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_92_ready),
		.io_addressIn_valid(io_connPE_92_valid),
		.io_addressIn_bits(io_connPE_92_bits),
		.io_addressOut_ready(_networkUnits_92_io_peAddress_ready),
		.io_addressOut_valid(_queues_92_io_addressOut_valid),
		.io_addressOut_bits(_queues_92_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_93(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_93_ready),
		.io_addressIn_valid(io_connPE_93_valid),
		.io_addressIn_bits(io_connPE_93_bits),
		.io_addressOut_ready(_networkUnits_93_io_peAddress_ready),
		.io_addressOut_valid(_queues_93_io_addressOut_valid),
		.io_addressOut_bits(_queues_93_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_94(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_94_ready),
		.io_addressIn_valid(io_connPE_94_valid),
		.io_addressIn_bits(io_connPE_94_bits),
		.io_addressOut_ready(_networkUnits_94_io_peAddress_ready),
		.io_addressOut_valid(_queues_94_io_addressOut_valid),
		.io_addressOut_bits(_queues_94_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_95(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_95_ready),
		.io_addressIn_valid(io_connPE_95_valid),
		.io_addressIn_bits(io_connPE_95_bits),
		.io_addressOut_ready(_networkUnits_95_io_peAddress_ready),
		.io_addressOut_valid(_queues_95_io_addressOut_valid),
		.io_addressOut_bits(_queues_95_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_96(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_96_ready),
		.io_addressIn_valid(io_connPE_96_valid),
		.io_addressIn_bits(io_connPE_96_bits),
		.io_addressOut_ready(_networkUnits_96_io_peAddress_ready),
		.io_addressOut_valid(_queues_96_io_addressOut_valid),
		.io_addressOut_bits(_queues_96_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_97(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_97_ready),
		.io_addressIn_valid(io_connPE_97_valid),
		.io_addressIn_bits(io_connPE_97_bits),
		.io_addressOut_ready(_networkUnits_97_io_peAddress_ready),
		.io_addressOut_valid(_queues_97_io_addressOut_valid),
		.io_addressOut_bits(_queues_97_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_98(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_98_ready),
		.io_addressIn_valid(io_connPE_98_valid),
		.io_addressIn_bits(io_connPE_98_bits),
		.io_addressOut_ready(_networkUnits_98_io_peAddress_ready),
		.io_addressOut_valid(_queues_98_io_addressOut_valid),
		.io_addressOut_bits(_queues_98_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_99(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_99_ready),
		.io_addressIn_valid(io_connPE_99_valid),
		.io_addressIn_bits(io_connPE_99_bits),
		.io_addressOut_ready(_networkUnits_99_io_peAddress_ready),
		.io_addressOut_valid(_queues_99_io_addressOut_valid),
		.io_addressOut_bits(_queues_99_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_100(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_100_ready),
		.io_addressIn_valid(io_connPE_100_valid),
		.io_addressIn_bits(io_connPE_100_bits),
		.io_addressOut_ready(_networkUnits_100_io_peAddress_ready),
		.io_addressOut_valid(_queues_100_io_addressOut_valid),
		.io_addressOut_bits(_queues_100_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_101(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_101_ready),
		.io_addressIn_valid(io_connPE_101_valid),
		.io_addressIn_bits(io_connPE_101_bits),
		.io_addressOut_ready(_networkUnits_101_io_peAddress_ready),
		.io_addressOut_valid(_queues_101_io_addressOut_valid),
		.io_addressOut_bits(_queues_101_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_102(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_102_ready),
		.io_addressIn_valid(io_connPE_102_valid),
		.io_addressIn_bits(io_connPE_102_bits),
		.io_addressOut_ready(_networkUnits_102_io_peAddress_ready),
		.io_addressOut_valid(_queues_102_io_addressOut_valid),
		.io_addressOut_bits(_queues_102_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_103(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_103_ready),
		.io_addressIn_valid(io_connPE_103_valid),
		.io_addressIn_bits(io_connPE_103_bits),
		.io_addressOut_ready(_networkUnits_103_io_peAddress_ready),
		.io_addressOut_valid(_queues_103_io_addressOut_valid),
		.io_addressOut_bits(_queues_103_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_104(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_104_ready),
		.io_addressIn_valid(io_connPE_104_valid),
		.io_addressIn_bits(io_connPE_104_bits),
		.io_addressOut_ready(_networkUnits_104_io_peAddress_ready),
		.io_addressOut_valid(_queues_104_io_addressOut_valid),
		.io_addressOut_bits(_queues_104_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_105(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_105_ready),
		.io_addressIn_valid(io_connPE_105_valid),
		.io_addressIn_bits(io_connPE_105_bits),
		.io_addressOut_ready(_networkUnits_105_io_peAddress_ready),
		.io_addressOut_valid(_queues_105_io_addressOut_valid),
		.io_addressOut_bits(_queues_105_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_106(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_106_ready),
		.io_addressIn_valid(io_connPE_106_valid),
		.io_addressIn_bits(io_connPE_106_bits),
		.io_addressOut_ready(_networkUnits_106_io_peAddress_ready),
		.io_addressOut_valid(_queues_106_io_addressOut_valid),
		.io_addressOut_bits(_queues_106_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_107(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_107_ready),
		.io_addressIn_valid(io_connPE_107_valid),
		.io_addressIn_bits(io_connPE_107_bits),
		.io_addressOut_ready(_networkUnits_107_io_peAddress_ready),
		.io_addressOut_valid(_queues_107_io_addressOut_valid),
		.io_addressOut_bits(_queues_107_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_108(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_108_ready),
		.io_addressIn_valid(io_connPE_108_valid),
		.io_addressIn_bits(io_connPE_108_bits),
		.io_addressOut_ready(_networkUnits_108_io_peAddress_ready),
		.io_addressOut_valid(_queues_108_io_addressOut_valid),
		.io_addressOut_bits(_queues_108_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_109(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_109_ready),
		.io_addressIn_valid(io_connPE_109_valid),
		.io_addressIn_bits(io_connPE_109_bits),
		.io_addressOut_ready(_networkUnits_109_io_peAddress_ready),
		.io_addressOut_valid(_queues_109_io_addressOut_valid),
		.io_addressOut_bits(_queues_109_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_110(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_110_ready),
		.io_addressIn_valid(io_connPE_110_valid),
		.io_addressIn_bits(io_connPE_110_bits),
		.io_addressOut_ready(_networkUnits_110_io_peAddress_ready),
		.io_addressOut_valid(_queues_110_io_addressOut_valid),
		.io_addressOut_bits(_queues_110_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_111(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_111_ready),
		.io_addressIn_valid(io_connPE_111_valid),
		.io_addressIn_bits(io_connPE_111_bits),
		.io_addressOut_ready(_networkUnits_111_io_peAddress_ready),
		.io_addressOut_valid(_queues_111_io_addressOut_valid),
		.io_addressOut_bits(_queues_111_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_112(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_112_ready),
		.io_addressIn_valid(io_connPE_112_valid),
		.io_addressIn_bits(io_connPE_112_bits),
		.io_addressOut_ready(_networkUnits_112_io_peAddress_ready),
		.io_addressOut_valid(_queues_112_io_addressOut_valid),
		.io_addressOut_bits(_queues_112_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_113(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_113_ready),
		.io_addressIn_valid(io_connPE_113_valid),
		.io_addressIn_bits(io_connPE_113_bits),
		.io_addressOut_ready(_networkUnits_113_io_peAddress_ready),
		.io_addressOut_valid(_queues_113_io_addressOut_valid),
		.io_addressOut_bits(_queues_113_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_114(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_114_ready),
		.io_addressIn_valid(io_connPE_114_valid),
		.io_addressIn_bits(io_connPE_114_bits),
		.io_addressOut_ready(_networkUnits_114_io_peAddress_ready),
		.io_addressOut_valid(_queues_114_io_addressOut_valid),
		.io_addressOut_bits(_queues_114_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_115(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_115_ready),
		.io_addressIn_valid(io_connPE_115_valid),
		.io_addressIn_bits(io_connPE_115_bits),
		.io_addressOut_ready(_networkUnits_115_io_peAddress_ready),
		.io_addressOut_valid(_queues_115_io_addressOut_valid),
		.io_addressOut_bits(_queues_115_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_116(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_116_ready),
		.io_addressIn_valid(io_connPE_116_valid),
		.io_addressIn_bits(io_connPE_116_bits),
		.io_addressOut_ready(_networkUnits_116_io_peAddress_ready),
		.io_addressOut_valid(_queues_116_io_addressOut_valid),
		.io_addressOut_bits(_queues_116_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_117(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_117_ready),
		.io_addressIn_valid(io_connPE_117_valid),
		.io_addressIn_bits(io_connPE_117_bits),
		.io_addressOut_ready(_networkUnits_117_io_peAddress_ready),
		.io_addressOut_valid(_queues_117_io_addressOut_valid),
		.io_addressOut_bits(_queues_117_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_118(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_118_ready),
		.io_addressIn_valid(io_connPE_118_valid),
		.io_addressIn_bits(io_connPE_118_bits),
		.io_addressOut_ready(_networkUnits_118_io_peAddress_ready),
		.io_addressOut_valid(_queues_118_io_addressOut_valid),
		.io_addressOut_bits(_queues_118_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_119(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_119_ready),
		.io_addressIn_valid(io_connPE_119_valid),
		.io_addressIn_bits(io_connPE_119_bits),
		.io_addressOut_ready(_networkUnits_119_io_peAddress_ready),
		.io_addressOut_valid(_queues_119_io_addressOut_valid),
		.io_addressOut_bits(_queues_119_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_120(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_120_ready),
		.io_addressIn_valid(io_connPE_120_valid),
		.io_addressIn_bits(io_connPE_120_bits),
		.io_addressOut_ready(_networkUnits_120_io_peAddress_ready),
		.io_addressOut_valid(_queues_120_io_addressOut_valid),
		.io_addressOut_bits(_queues_120_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_121(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_121_ready),
		.io_addressIn_valid(io_connPE_121_valid),
		.io_addressIn_bits(io_connPE_121_bits),
		.io_addressOut_ready(_networkUnits_121_io_peAddress_ready),
		.io_addressOut_valid(_queues_121_io_addressOut_valid),
		.io_addressOut_bits(_queues_121_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_122(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_122_ready),
		.io_addressIn_valid(io_connPE_122_valid),
		.io_addressIn_bits(io_connPE_122_bits),
		.io_addressOut_ready(_networkUnits_122_io_peAddress_ready),
		.io_addressOut_valid(_queues_122_io_addressOut_valid),
		.io_addressOut_bits(_queues_122_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_123(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_123_ready),
		.io_addressIn_valid(io_connPE_123_valid),
		.io_addressIn_bits(io_connPE_123_bits),
		.io_addressOut_ready(_networkUnits_123_io_peAddress_ready),
		.io_addressOut_valid(_queues_123_io_addressOut_valid),
		.io_addressOut_bits(_queues_123_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_124(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_124_ready),
		.io_addressIn_valid(io_connPE_124_valid),
		.io_addressIn_bits(io_connPE_124_bits),
		.io_addressOut_ready(_networkUnits_124_io_peAddress_ready),
		.io_addressOut_valid(_queues_124_io_addressOut_valid),
		.io_addressOut_bits(_queues_124_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_125(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_125_ready),
		.io_addressIn_valid(io_connPE_125_valid),
		.io_addressIn_bits(io_connPE_125_bits),
		.io_addressOut_ready(_networkUnits_125_io_peAddress_ready),
		.io_addressOut_valid(_queues_125_io_addressOut_valid),
		.io_addressOut_bits(_queues_125_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_126(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_126_ready),
		.io_addressIn_valid(io_connPE_126_valid),
		.io_addressIn_bits(io_connPE_126_bits),
		.io_addressOut_ready(_networkUnits_126_io_peAddress_ready),
		.io_addressOut_valid(_queues_126_io_addressOut_valid),
		.io_addressOut_bits(_queues_126_io_addressOut_bits)
	);
	AllocatorBuffer_64 queues_127(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_127_ready),
		.io_addressIn_valid(io_connPE_127_valid),
		.io_addressIn_bits(io_connPE_127_bits),
		.io_addressOut_ready(_networkUnits_127_io_peAddress_ready),
		.io_addressOut_valid(_queues_127_io_addressOut_valid),
		.io_addressOut_bits(_queues_127_io_addressOut_bits)
	);
endmodule
module ArgumentServer (
	clock,
	reset,
	io_connNetwork_ready,
	io_connNetwork_valid,
	io_connNetwork_bits,
	io_connStealNtw_ctrl_serveStealReq_valid,
	io_connStealNtw_ctrl_serveStealReq_ready,
	io_connStealNtw_data_qOutTask_ready,
	io_connStealNtw_data_qOutTask_valid,
	io_connStealNtw_data_qOutTask_bits,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_read_address_task_ready,
	io_read_address_task_valid,
	io_read_address_task_bits,
	io_read_data_task_ready,
	io_read_data_task_valid,
	io_read_data_task_bits
);
	input clock;
	input reset;
	output wire io_connNetwork_ready;
	input io_connNetwork_valid;
	input [63:0] io_connNetwork_bits;
	output wire io_connStealNtw_ctrl_serveStealReq_valid;
	input io_connStealNtw_ctrl_serveStealReq_ready;
	input io_connStealNtw_data_qOutTask_ready;
	output wire io_connStealNtw_data_qOutTask_valid;
	output wire [255:0] io_connStealNtw_data_qOutTask_bits;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [31:0] io_read_data_bits;
	input io_write_address_ready;
	output wire io_write_address_valid;
	output wire [63:0] io_write_address_bits;
	input io_write_data_ready;
	output wire io_write_data_valid;
	output wire [31:0] io_write_data_bits;
	input io_read_address_task_ready;
	output wire io_read_address_task_valid;
	output wire [63:0] io_read_address_task_bits;
	output wire io_read_data_task_ready;
	input io_read_data_task_valid;
	input [31:0] io_read_data_task_bits;
	wire _readyTasksQueue_io_enq_ready;
	wire _readyTasksQueue_io_deq_valid;
	wire [255:0] _readyTasksQueue_io_deq_bits;
	wire _addressesOfReadyTasks_io_enq_ready;
	wire _addressesOfReadyTasks_io_deq_valid;
	wire [63:0] _addressesOfReadyTasks_io_deq_bits;
	wire _addrNtwInQueue_io_deq_valid;
	wire [63:0] _addrNtwInQueue_io_deq_bits;
	reg [3:0] counterStateReg;
	reg [63:0] counterReg;
	reg [63:0] currReadAddr;
	reg [63:0] counterAddr;
	reg [63:0] addrMask;
	reg helpGarbageCollector;
	wire _GEN = counterStateReg == 4'h1;
	wire _GEN_0 = counterStateReg == 4'h2;
	wire _GEN_1 = counterStateReg == 4'h3;
	wire _GEN_2 = _GEN | _GEN_0;
	wire _GEN_3 = counterStateReg == 4'h4;
	wire _GEN_4 = counterStateReg == 4'h5;
	wire _GEN_5 = counterStateReg == 4'h7;
	wire _GEN_6 = ((_GEN | _GEN_0) | _GEN_1) | _GEN_3;
	reg [3:0] taskReadAddressStateReg;
	reg [63:0] taskAddr;
	wire _GEN_7 = taskReadAddressStateReg == 4'h6;
	wire _GEN_8 = taskReadAddressStateReg == 4'h8;
	reg [3:0] taskReadStateReg;
	reg [2:0] taskReadCount;
	reg [31:0] taskRegisters_0;
	reg [31:0] taskRegisters_1;
	reg [31:0] taskRegisters_2;
	reg [31:0] taskRegisters_3;
	reg [31:0] taskRegisters_4;
	reg [31:0] taskRegisters_5;
	reg [31:0] taskRegisters_6;
	reg [31:0] taskRegisters_7;
	wire io_read_data_task_ready_0 = taskReadStateReg == 4'h9;
	wire _GEN_9 = taskReadStateReg == 4'ha;
	reg [31:0] tasksGivenAwayCount;
	reg [255:0] taskReg;
	reg [3:0] taskWriteStateReg;
	wire _GEN_10 = taskWriteStateReg == 4'hb;
	wire _GEN_11 = taskWriteStateReg == 4'hc;
	wire io_connStealNtw_ctrl_serveStealReq_valid_0 = |tasksGivenAwayCount & (taskWriteStateReg != 4'hc);
	always @(posedge clock)
		if (reset) begin
			counterStateReg <= 4'h1;
			counterReg <= 64'h0000000000000000;
			currReadAddr <= 64'h0000000000000000;
			counterAddr <= 64'h0000000000000000;
			addrMask <= 64'h0000000000000000;
			helpGarbageCollector <= 1'h0;
			taskReadAddressStateReg <= 4'h6;
			taskAddr <= 64'h0000000000000000;
			taskReadStateReg <= 4'h9;
			taskReadCount <= 3'h7;
			taskRegisters_0 <= 32'h00000000;
			taskRegisters_1 <= 32'h00000000;
			taskRegisters_2 <= 32'h00000000;
			taskRegisters_3 <= 32'h00000000;
			taskRegisters_4 <= 32'h00000000;
			taskRegisters_5 <= 32'h00000000;
			taskRegisters_6 <= 32'h00000000;
			taskRegisters_7 <= 32'h00000000;
			tasksGivenAwayCount <= 32'h00000000;
			taskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			taskWriteStateReg <= 4'hb;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_12;
			reg _GEN_13;
			reg [2:0] _taskReadCount_T;
			reg _GEN_14;
			_GEN_12 = io_read_data_valid & (io_read_data_bits == 32'h00000001);
			_GEN_13 = _GEN_5 & _addressesOfReadyTasks_io_enq_ready;
			_taskReadCount_T = taskReadCount - 3'h1;
			_GEN_14 = _GEN_11 & io_connStealNtw_data_qOutTask_ready;
			if (_GEN) begin
				if (_addrNtwInQueue_io_deq_valid)
					counterStateReg <= 4'h2;
			end
			else if (_GEN_0) begin
				if (io_read_address_ready)
					counterStateReg <= 4'h3;
			end
			else if (_GEN_1) begin
				if (_GEN_12)
					counterStateReg <= 4'h7;
				else if (io_read_data_valid)
					counterStateReg <= 4'h4;
			end
			else if (_GEN_3) begin
				if (io_write_address_ready)
					counterStateReg <= 4'h5;
			end
			else if (_GEN_4) begin
				if (io_write_data_ready)
					counterStateReg <= 4'h1;
			end
			else if (_GEN_13)
				counterStateReg <= 4'h4;
			if (((_GEN_2 | ~_GEN_1) | _GEN_12) | ~io_read_data_valid)
				;
			else
				counterReg <= {32'h00000000, io_read_data_bits - 32'h00000001};
			if (_GEN_2 | ~(_GEN_1 & _GEN_12))
				;
			else
				currReadAddr <= counterAddr + 64'h0000000000000004;
			if (_GEN & _addrNtwInQueue_io_deq_valid)
				counterAddr <= _addrNtwInQueue_io_deq_bits & addrMask;
			addrMask <= 64'hffffffffffffffe0;
			if (~_GEN_6) begin
				if (_GEN_4)
					helpGarbageCollector <= ~io_write_data_ready & helpGarbageCollector;
				else
					helpGarbageCollector <= _GEN_13 | helpGarbageCollector;
			end
			if (_GEN_7) begin
				if (_addressesOfReadyTasks_io_deq_valid)
					taskReadAddressStateReg <= 4'h8;
			end
			else if (_GEN_8 & io_read_address_task_ready)
				taskReadAddressStateReg <= 4'h6;
			if (_GEN_7 & _addressesOfReadyTasks_io_deq_valid)
				taskAddr <= _addressesOfReadyTasks_io_deq_bits;
			if (io_read_data_task_ready_0) begin
				if ((taskReadCount == 3'h1) & io_read_data_task_valid)
					taskReadStateReg <= 4'ha;
				if (io_read_data_task_valid)
					taskReadCount <= _taskReadCount_T;
			end
			else if (_GEN_9 & _readyTasksQueue_io_enq_ready) begin
				taskReadStateReg <= 4'h9;
				taskReadCount <= 3'h7;
			end
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h0))
				taskRegisters_0 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h1))
				taskRegisters_1 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h2))
				taskRegisters_2 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h3))
				taskRegisters_3 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h4))
				taskRegisters_4 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h5))
				taskRegisters_5 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 3'h6))
				taskRegisters_6 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (&_taskReadCount_T))
				taskRegisters_7 <= io_read_data_task_bits;
			if (io_connStealNtw_ctrl_serveStealReq_valid_0 & io_connStealNtw_ctrl_serveStealReq_ready)
				tasksGivenAwayCount <= tasksGivenAwayCount - 32'h00000001;
			else if (_GEN_10 | ~_GEN_14)
				;
			else
				tasksGivenAwayCount <= tasksGivenAwayCount + 32'h00000001;
			if (_GEN_10 & _readyTasksQueue_io_deq_valid)
				taskReg <= _readyTasksQueue_io_deq_bits;
			if (_GEN_10) begin
				if (_readyTasksQueue_io_deq_valid)
					taskWriteStateReg <= 4'hc;
			end
			else if (_GEN_14)
				taskWriteStateReg <= 4'hb;
		end
	Queue16_UInt_4 addrNtwInQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_connNetwork_ready),
		.io_enq_valid(io_connNetwork_valid),
		.io_enq_bits(io_connNetwork_bits),
		.io_deq_ready(_GEN),
		.io_deq_valid(_addrNtwInQueue_io_deq_valid),
		.io_deq_bits(_addrNtwInQueue_io_deq_bits)
	);
	Queue16_UInt_4 addressesOfReadyTasks(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_addressesOfReadyTasks_io_enq_ready),
		.io_enq_valid(~((((_GEN | _GEN_0) | _GEN_1) | _GEN_3) | _GEN_4) & _GEN_5),
		.io_enq_bits(currReadAddr),
		.io_deq_ready(_GEN_7),
		.io_deq_valid(_addressesOfReadyTasks_io_deq_valid),
		.io_deq_bits(_addressesOfReadyTasks_io_deq_bits)
	);
	Queue16_UInt_2 readyTasksQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_readyTasksQueue_io_enq_ready),
		.io_enq_valid(~io_read_data_task_ready_0 & _GEN_9),
		.io_enq_bits({taskRegisters_0, taskRegisters_1, taskRegisters_2, taskRegisters_3, taskRegisters_4, taskRegisters_5, taskRegisters_6, taskRegisters_7}),
		.io_deq_ready(_GEN_10),
		.io_deq_valid(_readyTasksQueue_io_deq_valid),
		.io_deq_bits(_readyTasksQueue_io_deq_bits),
		.io_count()
	);
	assign io_connStealNtw_ctrl_serveStealReq_valid = io_connStealNtw_ctrl_serveStealReq_valid_0;
	assign io_connStealNtw_data_qOutTask_valid = ~_GEN_10 & _GEN_11;
	assign io_connStealNtw_data_qOutTask_bits = taskReg;
	assign io_read_address_valid = ~_GEN & _GEN_0;
	assign io_read_address_bits = counterAddr;
	assign io_read_data_ready = ~_GEN_2 & _GEN_1;
	assign io_write_address_valid = ~((_GEN | _GEN_0) | _GEN_1) & _GEN_3;
	assign io_write_address_bits = counterAddr;
	assign io_write_data_valid = ~_GEN_6 & _GEN_4;
	assign io_write_data_bits = (helpGarbageCollector ? 32'h01000000 : counterReg[31:0]);
	assign io_read_address_task_valid = ~_GEN_7 & _GEN_8;
	assign io_read_address_task_bits = (_GEN_7 | ~_GEN_8 ? 64'h0000000000000000 : taskAddr);
	assign io_read_data_task_ready = io_read_data_task_ready_0;
endmodule
module RVtoAXIBridge_8 (
	clock,
	reset,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data,
	axi_aw_ready,
	axi_aw_valid,
	axi_aw_bits_addr,
	axi_w_ready,
	axi_w_valid,
	axi_w_bits_data,
	axi_b_valid
);
	input clock;
	input reset;
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [31:0] io_read_data_bits;
	output wire io_write_address_ready;
	input io_write_address_valid;
	input [63:0] io_write_address_bits;
	output wire io_write_data_ready;
	input io_write_data_valid;
	input [31:0] io_write_data_bits;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire axi_r_ready;
	input axi_r_valid;
	input [31:0] axi_r_bits_data;
	input axi_aw_ready;
	output wire axi_aw_valid;
	output wire [63:0] axi_aw_bits_addr;
	input axi_w_ready;
	output wire axi_w_valid;
	output wire [31:0] axi_w_bits_data;
	input axi_b_valid;
	reg [1:0] writeDataDone;
	reg writeHandshakeDetector;
	wire axi_w_valid_0 = (io_write_data_valid & axi_w_ready) & ~writeHandshakeDetector;
	always @(posedge clock)
		if (reset) begin
			writeDataDone <= 2'h0;
			writeHandshakeDetector <= 1'h0;
		end
		else begin
			if ((writeDataDone == 2'h0) & axi_w_ready)
				writeDataDone <= 2'h1;
			else if ((writeDataDone == 2'h1) & axi_b_valid)
				writeDataDone <= 2'h0;
			writeHandshakeDetector <= axi_w_valid_0 | (~axi_b_valid & writeHandshakeDetector);
		end
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign io_write_address_ready = axi_aw_ready;
	assign io_write_data_ready = (writeDataDone == 2'h1) & axi_b_valid;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_r_ready = io_read_data_ready;
	assign axi_aw_valid = io_write_address_valid;
	assign axi_aw_bits_addr = io_write_address_bits;
	assign axi_w_valid = axi_w_valid_0;
	assign axi_w_bits_data = io_write_data_bits;
endmodule
module RVtoAXIBridge_24 (
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data
);
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [31:0] io_read_data_bits;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire axi_r_ready;
	input axi_r_valid;
	input [31:0] axi_r_bits_data;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_r_ready = io_read_data_ready;
endmodule
module ram_2x32 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [31:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [31:0] W0_data;
	reg [31:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel_16 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [31:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [31:0] io_deq_bits_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x32 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_data)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module ram_2x37 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [36:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [36:0] W0_data;
	reg [36:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 37'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteDataChannel_16 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [31:0] io_enq_bits_data;
	input [3:0] io_enq_bits_strb;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [31:0] io_deq_bits_data;
	output wire [3:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	wire [36:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_deq == do_enq))
				maybe_full <= do_enq;
		end
	ram_2x37 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_strb, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[31:0];
	assign io_deq_bits_strb = _ram_ext_R0_data[35:32];
	assign io_deq_bits_last = _ram_ext_R0_data[36];
endmodule
module Queue2_WriteResponseChannel_16 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_deq_ready,
	io_deq_valid
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_deq_ready;
	output wire io_deq_valid;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_enq;
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			do_enq = ~full & io_enq_valid;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module ram_2x98 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [97:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [97:0] W0_data;
	reg [97:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 98'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadAddressChannel_43 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [4:0] io_enq_bits_id;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [4:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [97:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x98 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[4:0];
	assign io_deq_bits_addr = _ram_ext_R0_data[68:5];
	assign io_deq_bits_len = _ram_ext_R0_data[76:69];
	assign io_deq_bits_size = _ram_ext_R0_data[79:77];
	assign io_deq_bits_burst = _ram_ext_R0_data[81:80];
	assign io_deq_bits_lock = _ram_ext_R0_data[82];
	assign io_deq_bits_cache = _ram_ext_R0_data[86:83];
	assign io_deq_bits_prot = _ram_ext_R0_data[89:87];
	assign io_deq_bits_qos = _ram_ext_R0_data[93:90];
	assign io_deq_bits_region = _ram_ext_R0_data[97:94];
endmodule
module ram_2x40 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [39:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [39:0] W0_data;
	reg [39:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel_48 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_data,
	io_deq_bits_resp,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [4:0] io_enq_bits_id;
	input [31:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [4:0] io_deq_bits_id;
	output wire [31:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	output wire io_deq_bits_last;
	wire [39:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x40 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_last, io_enq_bits_resp, io_enq_bits_data, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[4:0];
	assign io_deq_bits_data = _ram_ext_R0_data[36:5];
	assign io_deq_bits_resp = _ram_ext_R0_data[38:37];
	assign io_deq_bits_last = _ram_ext_R0_data[39];
endmodule
module Queue2_WriteAddressChannel_43 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_enq_bits_lock,
	io_enq_bits_cache,
	io_enq_bits_prot,
	io_enq_bits_qos,
	io_enq_bits_region,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [4:0] io_enq_bits_id;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_enq_bits_lock;
	input [3:0] io_enq_bits_cache;
	input [2:0] io_enq_bits_prot;
	input [3:0] io_enq_bits_qos;
	input [3:0] io_enq_bits_region;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [4:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [97:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x98 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_region, io_enq_bits_qos, io_enq_bits_prot, io_enq_bits_cache, io_enq_bits_lock, io_enq_bits_burst, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr, io_enq_bits_id})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_id = _ram_ext_R0_data[4:0];
	assign io_deq_bits_addr = _ram_ext_R0_data[68:5];
	assign io_deq_bits_len = _ram_ext_R0_data[76:69];
	assign io_deq_bits_size = _ram_ext_R0_data[79:77];
	assign io_deq_bits_burst = _ram_ext_R0_data[81:80];
	assign io_deq_bits_lock = _ram_ext_R0_data[82];
	assign io_deq_bits_cache = _ram_ext_R0_data[86:83];
	assign io_deq_bits_prot = _ram_ext_R0_data[89:87];
	assign io_deq_bits_qos = _ram_ext_R0_data[93:90];
	assign io_deq_bits_region = _ram_ext_R0_data[97:94];
endmodule
module ram_2x5 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [4:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [4:0] W0_data;
	reg [4:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 5'bxxxxx);
endmodule
module Queue2_WriteResponseChannel_48 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [4:0] io_enq_bits_id;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [4:0] io_deq_bits_id;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x5 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_id),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_id)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module elasticArbiter_6 (
	clock,
	reset,
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_addr,
	io_sources_0_bits_len,
	io_sources_0_bits_size,
	io_sources_0_bits_burst,
	io_sources_0_bits_lock,
	io_sources_0_bits_cache,
	io_sources_0_bits_prot,
	io_sources_0_bits_qos,
	io_sources_0_bits_region,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_addr,
	io_sources_1_bits_len,
	io_sources_1_bits_size,
	io_sources_1_bits_burst,
	io_sources_1_bits_lock,
	io_sources_1_bits_cache,
	io_sources_1_bits_prot,
	io_sources_1_bits_qos,
	io_sources_1_bits_region,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_addr,
	io_sources_2_bits_len,
	io_sources_2_bits_size,
	io_sources_2_bits_burst,
	io_sources_2_bits_lock,
	io_sources_2_bits_cache,
	io_sources_2_bits_prot,
	io_sources_2_bits_qos,
	io_sources_2_bits_region,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_addr,
	io_sources_3_bits_len,
	io_sources_3_bits_size,
	io_sources_3_bits_burst,
	io_sources_3_bits_lock,
	io_sources_3_bits_cache,
	io_sources_3_bits_prot,
	io_sources_3_bits_qos,
	io_sources_3_bits_region,
	io_sources_4_ready,
	io_sources_4_valid,
	io_sources_4_bits_addr,
	io_sources_4_bits_len,
	io_sources_4_bits_size,
	io_sources_4_bits_burst,
	io_sources_4_bits_lock,
	io_sources_4_bits_cache,
	io_sources_4_bits_prot,
	io_sources_4_bits_qos,
	io_sources_4_bits_region,
	io_sources_5_ready,
	io_sources_5_valid,
	io_sources_5_bits_addr,
	io_sources_5_bits_len,
	io_sources_5_bits_size,
	io_sources_5_bits_burst,
	io_sources_5_bits_lock,
	io_sources_5_bits_cache,
	io_sources_5_bits_prot,
	io_sources_5_bits_qos,
	io_sources_5_bits_region,
	io_sources_6_ready,
	io_sources_6_valid,
	io_sources_6_bits_addr,
	io_sources_6_bits_len,
	io_sources_6_bits_size,
	io_sources_6_bits_burst,
	io_sources_6_bits_lock,
	io_sources_6_bits_cache,
	io_sources_6_bits_prot,
	io_sources_6_bits_qos,
	io_sources_6_bits_region,
	io_sources_7_ready,
	io_sources_7_valid,
	io_sources_7_bits_addr,
	io_sources_7_bits_len,
	io_sources_7_bits_size,
	io_sources_7_bits_burst,
	io_sources_7_bits_lock,
	io_sources_7_bits_cache,
	io_sources_7_bits_prot,
	io_sources_7_bits_qos,
	io_sources_7_bits_region,
	io_sources_8_ready,
	io_sources_8_valid,
	io_sources_8_bits_addr,
	io_sources_8_bits_len,
	io_sources_8_bits_size,
	io_sources_8_bits_burst,
	io_sources_8_bits_lock,
	io_sources_8_bits_cache,
	io_sources_8_bits_prot,
	io_sources_8_bits_qos,
	io_sources_8_bits_region,
	io_sources_9_ready,
	io_sources_9_valid,
	io_sources_9_bits_addr,
	io_sources_9_bits_len,
	io_sources_9_bits_size,
	io_sources_9_bits_burst,
	io_sources_9_bits_lock,
	io_sources_9_bits_cache,
	io_sources_9_bits_prot,
	io_sources_9_bits_qos,
	io_sources_9_bits_region,
	io_sources_10_ready,
	io_sources_10_valid,
	io_sources_10_bits_addr,
	io_sources_10_bits_len,
	io_sources_10_bits_size,
	io_sources_10_bits_burst,
	io_sources_10_bits_lock,
	io_sources_10_bits_cache,
	io_sources_10_bits_prot,
	io_sources_10_bits_qos,
	io_sources_10_bits_region,
	io_sources_11_ready,
	io_sources_11_valid,
	io_sources_11_bits_addr,
	io_sources_11_bits_len,
	io_sources_11_bits_size,
	io_sources_11_bits_burst,
	io_sources_11_bits_lock,
	io_sources_11_bits_cache,
	io_sources_11_bits_prot,
	io_sources_11_bits_qos,
	io_sources_11_bits_region,
	io_sources_12_ready,
	io_sources_12_valid,
	io_sources_12_bits_addr,
	io_sources_12_bits_len,
	io_sources_12_bits_size,
	io_sources_12_bits_burst,
	io_sources_12_bits_lock,
	io_sources_12_bits_cache,
	io_sources_12_bits_prot,
	io_sources_12_bits_qos,
	io_sources_12_bits_region,
	io_sources_13_ready,
	io_sources_13_valid,
	io_sources_13_bits_addr,
	io_sources_13_bits_len,
	io_sources_13_bits_size,
	io_sources_13_bits_burst,
	io_sources_13_bits_lock,
	io_sources_13_bits_cache,
	io_sources_13_bits_prot,
	io_sources_13_bits_qos,
	io_sources_13_bits_region,
	io_sources_14_ready,
	io_sources_14_valid,
	io_sources_14_bits_addr,
	io_sources_14_bits_len,
	io_sources_14_bits_size,
	io_sources_14_bits_burst,
	io_sources_14_bits_lock,
	io_sources_14_bits_cache,
	io_sources_14_bits_prot,
	io_sources_14_bits_qos,
	io_sources_14_bits_region,
	io_sources_15_ready,
	io_sources_15_valid,
	io_sources_15_bits_addr,
	io_sources_15_bits_len,
	io_sources_15_bits_size,
	io_sources_15_bits_burst,
	io_sources_15_bits_lock,
	io_sources_15_bits_cache,
	io_sources_15_bits_prot,
	io_sources_15_bits_qos,
	io_sources_15_bits_region,
	io_sources_16_ready,
	io_sources_16_valid,
	io_sources_16_bits_addr,
	io_sources_16_bits_len,
	io_sources_16_bits_size,
	io_sources_16_bits_burst,
	io_sources_16_bits_lock,
	io_sources_16_bits_cache,
	io_sources_16_bits_prot,
	io_sources_16_bits_qos,
	io_sources_16_bits_region,
	io_sources_17_ready,
	io_sources_17_valid,
	io_sources_17_bits_addr,
	io_sources_17_bits_len,
	io_sources_17_bits_size,
	io_sources_17_bits_burst,
	io_sources_17_bits_lock,
	io_sources_17_bits_cache,
	io_sources_17_bits_prot,
	io_sources_17_bits_qos,
	io_sources_17_bits_region,
	io_sources_18_ready,
	io_sources_18_valid,
	io_sources_18_bits_addr,
	io_sources_18_bits_len,
	io_sources_18_bits_size,
	io_sources_18_bits_burst,
	io_sources_18_bits_lock,
	io_sources_18_bits_cache,
	io_sources_18_bits_prot,
	io_sources_18_bits_qos,
	io_sources_18_bits_region,
	io_sources_19_ready,
	io_sources_19_valid,
	io_sources_19_bits_addr,
	io_sources_19_bits_len,
	io_sources_19_bits_size,
	io_sources_19_bits_burst,
	io_sources_19_bits_lock,
	io_sources_19_bits_cache,
	io_sources_19_bits_prot,
	io_sources_19_bits_qos,
	io_sources_19_bits_region,
	io_sources_20_ready,
	io_sources_20_valid,
	io_sources_20_bits_addr,
	io_sources_20_bits_len,
	io_sources_20_bits_size,
	io_sources_20_bits_burst,
	io_sources_20_bits_lock,
	io_sources_20_bits_cache,
	io_sources_20_bits_prot,
	io_sources_20_bits_qos,
	io_sources_20_bits_region,
	io_sources_21_ready,
	io_sources_21_valid,
	io_sources_21_bits_addr,
	io_sources_21_bits_len,
	io_sources_21_bits_size,
	io_sources_21_bits_burst,
	io_sources_21_bits_lock,
	io_sources_21_bits_cache,
	io_sources_21_bits_prot,
	io_sources_21_bits_qos,
	io_sources_21_bits_region,
	io_sources_22_ready,
	io_sources_22_valid,
	io_sources_22_bits_addr,
	io_sources_22_bits_len,
	io_sources_22_bits_size,
	io_sources_22_bits_burst,
	io_sources_22_bits_lock,
	io_sources_22_bits_cache,
	io_sources_22_bits_prot,
	io_sources_22_bits_qos,
	io_sources_22_bits_region,
	io_sources_23_ready,
	io_sources_23_valid,
	io_sources_23_bits_addr,
	io_sources_23_bits_len,
	io_sources_23_bits_size,
	io_sources_23_bits_burst,
	io_sources_23_bits_lock,
	io_sources_23_bits_cache,
	io_sources_23_bits_prot,
	io_sources_23_bits_qos,
	io_sources_23_bits_region,
	io_sources_24_ready,
	io_sources_24_valid,
	io_sources_24_bits_addr,
	io_sources_24_bits_len,
	io_sources_24_bits_size,
	io_sources_24_bits_burst,
	io_sources_24_bits_lock,
	io_sources_24_bits_cache,
	io_sources_24_bits_prot,
	io_sources_24_bits_qos,
	io_sources_24_bits_region,
	io_sources_25_ready,
	io_sources_25_valid,
	io_sources_25_bits_addr,
	io_sources_25_bits_len,
	io_sources_25_bits_size,
	io_sources_25_bits_burst,
	io_sources_25_bits_lock,
	io_sources_25_bits_cache,
	io_sources_25_bits_prot,
	io_sources_25_bits_qos,
	io_sources_25_bits_region,
	io_sources_26_ready,
	io_sources_26_valid,
	io_sources_26_bits_addr,
	io_sources_26_bits_len,
	io_sources_26_bits_size,
	io_sources_26_bits_burst,
	io_sources_26_bits_lock,
	io_sources_26_bits_cache,
	io_sources_26_bits_prot,
	io_sources_26_bits_qos,
	io_sources_26_bits_region,
	io_sources_27_ready,
	io_sources_27_valid,
	io_sources_27_bits_addr,
	io_sources_27_bits_len,
	io_sources_27_bits_size,
	io_sources_27_bits_burst,
	io_sources_27_bits_lock,
	io_sources_27_bits_cache,
	io_sources_27_bits_prot,
	io_sources_27_bits_qos,
	io_sources_27_bits_region,
	io_sources_28_ready,
	io_sources_28_valid,
	io_sources_28_bits_addr,
	io_sources_28_bits_len,
	io_sources_28_bits_size,
	io_sources_28_bits_burst,
	io_sources_28_bits_lock,
	io_sources_28_bits_cache,
	io_sources_28_bits_prot,
	io_sources_28_bits_qos,
	io_sources_28_bits_region,
	io_sources_29_ready,
	io_sources_29_valid,
	io_sources_29_bits_addr,
	io_sources_29_bits_len,
	io_sources_29_bits_size,
	io_sources_29_bits_burst,
	io_sources_29_bits_lock,
	io_sources_29_bits_cache,
	io_sources_29_bits_prot,
	io_sources_29_bits_qos,
	io_sources_29_bits_region,
	io_sources_30_ready,
	io_sources_30_valid,
	io_sources_30_bits_addr,
	io_sources_30_bits_len,
	io_sources_30_bits_size,
	io_sources_30_bits_burst,
	io_sources_30_bits_lock,
	io_sources_30_bits_cache,
	io_sources_30_bits_prot,
	io_sources_30_bits_qos,
	io_sources_30_bits_region,
	io_sources_31_ready,
	io_sources_31_valid,
	io_sources_31_bits_addr,
	io_sources_31_bits_len,
	io_sources_31_bits_size,
	io_sources_31_bits_burst,
	io_sources_31_bits_lock,
	io_sources_31_bits_cache,
	io_sources_31_bits_prot,
	io_sources_31_bits_qos,
	io_sources_31_bits_region,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_id,
	io_sink_bits_addr,
	io_sink_bits_len,
	io_sink_bits_size,
	io_sink_bits_burst,
	io_sink_bits_lock,
	io_sink_bits_cache,
	io_sink_bits_prot,
	io_sink_bits_qos,
	io_sink_bits_region,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	input clock;
	input reset;
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [63:0] io_sources_0_bits_addr;
	input [7:0] io_sources_0_bits_len;
	input [2:0] io_sources_0_bits_size;
	input [1:0] io_sources_0_bits_burst;
	input io_sources_0_bits_lock;
	input [3:0] io_sources_0_bits_cache;
	input [2:0] io_sources_0_bits_prot;
	input [3:0] io_sources_0_bits_qos;
	input [3:0] io_sources_0_bits_region;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [63:0] io_sources_1_bits_addr;
	input [7:0] io_sources_1_bits_len;
	input [2:0] io_sources_1_bits_size;
	input [1:0] io_sources_1_bits_burst;
	input io_sources_1_bits_lock;
	input [3:0] io_sources_1_bits_cache;
	input [2:0] io_sources_1_bits_prot;
	input [3:0] io_sources_1_bits_qos;
	input [3:0] io_sources_1_bits_region;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [63:0] io_sources_2_bits_addr;
	input [7:0] io_sources_2_bits_len;
	input [2:0] io_sources_2_bits_size;
	input [1:0] io_sources_2_bits_burst;
	input io_sources_2_bits_lock;
	input [3:0] io_sources_2_bits_cache;
	input [2:0] io_sources_2_bits_prot;
	input [3:0] io_sources_2_bits_qos;
	input [3:0] io_sources_2_bits_region;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [63:0] io_sources_3_bits_addr;
	input [7:0] io_sources_3_bits_len;
	input [2:0] io_sources_3_bits_size;
	input [1:0] io_sources_3_bits_burst;
	input io_sources_3_bits_lock;
	input [3:0] io_sources_3_bits_cache;
	input [2:0] io_sources_3_bits_prot;
	input [3:0] io_sources_3_bits_qos;
	input [3:0] io_sources_3_bits_region;
	output wire io_sources_4_ready;
	input io_sources_4_valid;
	input [63:0] io_sources_4_bits_addr;
	input [7:0] io_sources_4_bits_len;
	input [2:0] io_sources_4_bits_size;
	input [1:0] io_sources_4_bits_burst;
	input io_sources_4_bits_lock;
	input [3:0] io_sources_4_bits_cache;
	input [2:0] io_sources_4_bits_prot;
	input [3:0] io_sources_4_bits_qos;
	input [3:0] io_sources_4_bits_region;
	output wire io_sources_5_ready;
	input io_sources_5_valid;
	input [63:0] io_sources_5_bits_addr;
	input [7:0] io_sources_5_bits_len;
	input [2:0] io_sources_5_bits_size;
	input [1:0] io_sources_5_bits_burst;
	input io_sources_5_bits_lock;
	input [3:0] io_sources_5_bits_cache;
	input [2:0] io_sources_5_bits_prot;
	input [3:0] io_sources_5_bits_qos;
	input [3:0] io_sources_5_bits_region;
	output wire io_sources_6_ready;
	input io_sources_6_valid;
	input [63:0] io_sources_6_bits_addr;
	input [7:0] io_sources_6_bits_len;
	input [2:0] io_sources_6_bits_size;
	input [1:0] io_sources_6_bits_burst;
	input io_sources_6_bits_lock;
	input [3:0] io_sources_6_bits_cache;
	input [2:0] io_sources_6_bits_prot;
	input [3:0] io_sources_6_bits_qos;
	input [3:0] io_sources_6_bits_region;
	output wire io_sources_7_ready;
	input io_sources_7_valid;
	input [63:0] io_sources_7_bits_addr;
	input [7:0] io_sources_7_bits_len;
	input [2:0] io_sources_7_bits_size;
	input [1:0] io_sources_7_bits_burst;
	input io_sources_7_bits_lock;
	input [3:0] io_sources_7_bits_cache;
	input [2:0] io_sources_7_bits_prot;
	input [3:0] io_sources_7_bits_qos;
	input [3:0] io_sources_7_bits_region;
	output wire io_sources_8_ready;
	input io_sources_8_valid;
	input [63:0] io_sources_8_bits_addr;
	input [7:0] io_sources_8_bits_len;
	input [2:0] io_sources_8_bits_size;
	input [1:0] io_sources_8_bits_burst;
	input io_sources_8_bits_lock;
	input [3:0] io_sources_8_bits_cache;
	input [2:0] io_sources_8_bits_prot;
	input [3:0] io_sources_8_bits_qos;
	input [3:0] io_sources_8_bits_region;
	output wire io_sources_9_ready;
	input io_sources_9_valid;
	input [63:0] io_sources_9_bits_addr;
	input [7:0] io_sources_9_bits_len;
	input [2:0] io_sources_9_bits_size;
	input [1:0] io_sources_9_bits_burst;
	input io_sources_9_bits_lock;
	input [3:0] io_sources_9_bits_cache;
	input [2:0] io_sources_9_bits_prot;
	input [3:0] io_sources_9_bits_qos;
	input [3:0] io_sources_9_bits_region;
	output wire io_sources_10_ready;
	input io_sources_10_valid;
	input [63:0] io_sources_10_bits_addr;
	input [7:0] io_sources_10_bits_len;
	input [2:0] io_sources_10_bits_size;
	input [1:0] io_sources_10_bits_burst;
	input io_sources_10_bits_lock;
	input [3:0] io_sources_10_bits_cache;
	input [2:0] io_sources_10_bits_prot;
	input [3:0] io_sources_10_bits_qos;
	input [3:0] io_sources_10_bits_region;
	output wire io_sources_11_ready;
	input io_sources_11_valid;
	input [63:0] io_sources_11_bits_addr;
	input [7:0] io_sources_11_bits_len;
	input [2:0] io_sources_11_bits_size;
	input [1:0] io_sources_11_bits_burst;
	input io_sources_11_bits_lock;
	input [3:0] io_sources_11_bits_cache;
	input [2:0] io_sources_11_bits_prot;
	input [3:0] io_sources_11_bits_qos;
	input [3:0] io_sources_11_bits_region;
	output wire io_sources_12_ready;
	input io_sources_12_valid;
	input [63:0] io_sources_12_bits_addr;
	input [7:0] io_sources_12_bits_len;
	input [2:0] io_sources_12_bits_size;
	input [1:0] io_sources_12_bits_burst;
	input io_sources_12_bits_lock;
	input [3:0] io_sources_12_bits_cache;
	input [2:0] io_sources_12_bits_prot;
	input [3:0] io_sources_12_bits_qos;
	input [3:0] io_sources_12_bits_region;
	output wire io_sources_13_ready;
	input io_sources_13_valid;
	input [63:0] io_sources_13_bits_addr;
	input [7:0] io_sources_13_bits_len;
	input [2:0] io_sources_13_bits_size;
	input [1:0] io_sources_13_bits_burst;
	input io_sources_13_bits_lock;
	input [3:0] io_sources_13_bits_cache;
	input [2:0] io_sources_13_bits_prot;
	input [3:0] io_sources_13_bits_qos;
	input [3:0] io_sources_13_bits_region;
	output wire io_sources_14_ready;
	input io_sources_14_valid;
	input [63:0] io_sources_14_bits_addr;
	input [7:0] io_sources_14_bits_len;
	input [2:0] io_sources_14_bits_size;
	input [1:0] io_sources_14_bits_burst;
	input io_sources_14_bits_lock;
	input [3:0] io_sources_14_bits_cache;
	input [2:0] io_sources_14_bits_prot;
	input [3:0] io_sources_14_bits_qos;
	input [3:0] io_sources_14_bits_region;
	output wire io_sources_15_ready;
	input io_sources_15_valid;
	input [63:0] io_sources_15_bits_addr;
	input [7:0] io_sources_15_bits_len;
	input [2:0] io_sources_15_bits_size;
	input [1:0] io_sources_15_bits_burst;
	input io_sources_15_bits_lock;
	input [3:0] io_sources_15_bits_cache;
	input [2:0] io_sources_15_bits_prot;
	input [3:0] io_sources_15_bits_qos;
	input [3:0] io_sources_15_bits_region;
	output wire io_sources_16_ready;
	input io_sources_16_valid;
	input [63:0] io_sources_16_bits_addr;
	input [7:0] io_sources_16_bits_len;
	input [2:0] io_sources_16_bits_size;
	input [1:0] io_sources_16_bits_burst;
	input io_sources_16_bits_lock;
	input [3:0] io_sources_16_bits_cache;
	input [2:0] io_sources_16_bits_prot;
	input [3:0] io_sources_16_bits_qos;
	input [3:0] io_sources_16_bits_region;
	output wire io_sources_17_ready;
	input io_sources_17_valid;
	input [63:0] io_sources_17_bits_addr;
	input [7:0] io_sources_17_bits_len;
	input [2:0] io_sources_17_bits_size;
	input [1:0] io_sources_17_bits_burst;
	input io_sources_17_bits_lock;
	input [3:0] io_sources_17_bits_cache;
	input [2:0] io_sources_17_bits_prot;
	input [3:0] io_sources_17_bits_qos;
	input [3:0] io_sources_17_bits_region;
	output wire io_sources_18_ready;
	input io_sources_18_valid;
	input [63:0] io_sources_18_bits_addr;
	input [7:0] io_sources_18_bits_len;
	input [2:0] io_sources_18_bits_size;
	input [1:0] io_sources_18_bits_burst;
	input io_sources_18_bits_lock;
	input [3:0] io_sources_18_bits_cache;
	input [2:0] io_sources_18_bits_prot;
	input [3:0] io_sources_18_bits_qos;
	input [3:0] io_sources_18_bits_region;
	output wire io_sources_19_ready;
	input io_sources_19_valid;
	input [63:0] io_sources_19_bits_addr;
	input [7:0] io_sources_19_bits_len;
	input [2:0] io_sources_19_bits_size;
	input [1:0] io_sources_19_bits_burst;
	input io_sources_19_bits_lock;
	input [3:0] io_sources_19_bits_cache;
	input [2:0] io_sources_19_bits_prot;
	input [3:0] io_sources_19_bits_qos;
	input [3:0] io_sources_19_bits_region;
	output wire io_sources_20_ready;
	input io_sources_20_valid;
	input [63:0] io_sources_20_bits_addr;
	input [7:0] io_sources_20_bits_len;
	input [2:0] io_sources_20_bits_size;
	input [1:0] io_sources_20_bits_burst;
	input io_sources_20_bits_lock;
	input [3:0] io_sources_20_bits_cache;
	input [2:0] io_sources_20_bits_prot;
	input [3:0] io_sources_20_bits_qos;
	input [3:0] io_sources_20_bits_region;
	output wire io_sources_21_ready;
	input io_sources_21_valid;
	input [63:0] io_sources_21_bits_addr;
	input [7:0] io_sources_21_bits_len;
	input [2:0] io_sources_21_bits_size;
	input [1:0] io_sources_21_bits_burst;
	input io_sources_21_bits_lock;
	input [3:0] io_sources_21_bits_cache;
	input [2:0] io_sources_21_bits_prot;
	input [3:0] io_sources_21_bits_qos;
	input [3:0] io_sources_21_bits_region;
	output wire io_sources_22_ready;
	input io_sources_22_valid;
	input [63:0] io_sources_22_bits_addr;
	input [7:0] io_sources_22_bits_len;
	input [2:0] io_sources_22_bits_size;
	input [1:0] io_sources_22_bits_burst;
	input io_sources_22_bits_lock;
	input [3:0] io_sources_22_bits_cache;
	input [2:0] io_sources_22_bits_prot;
	input [3:0] io_sources_22_bits_qos;
	input [3:0] io_sources_22_bits_region;
	output wire io_sources_23_ready;
	input io_sources_23_valid;
	input [63:0] io_sources_23_bits_addr;
	input [7:0] io_sources_23_bits_len;
	input [2:0] io_sources_23_bits_size;
	input [1:0] io_sources_23_bits_burst;
	input io_sources_23_bits_lock;
	input [3:0] io_sources_23_bits_cache;
	input [2:0] io_sources_23_bits_prot;
	input [3:0] io_sources_23_bits_qos;
	input [3:0] io_sources_23_bits_region;
	output wire io_sources_24_ready;
	input io_sources_24_valid;
	input [63:0] io_sources_24_bits_addr;
	input [7:0] io_sources_24_bits_len;
	input [2:0] io_sources_24_bits_size;
	input [1:0] io_sources_24_bits_burst;
	input io_sources_24_bits_lock;
	input [3:0] io_sources_24_bits_cache;
	input [2:0] io_sources_24_bits_prot;
	input [3:0] io_sources_24_bits_qos;
	input [3:0] io_sources_24_bits_region;
	output wire io_sources_25_ready;
	input io_sources_25_valid;
	input [63:0] io_sources_25_bits_addr;
	input [7:0] io_sources_25_bits_len;
	input [2:0] io_sources_25_bits_size;
	input [1:0] io_sources_25_bits_burst;
	input io_sources_25_bits_lock;
	input [3:0] io_sources_25_bits_cache;
	input [2:0] io_sources_25_bits_prot;
	input [3:0] io_sources_25_bits_qos;
	input [3:0] io_sources_25_bits_region;
	output wire io_sources_26_ready;
	input io_sources_26_valid;
	input [63:0] io_sources_26_bits_addr;
	input [7:0] io_sources_26_bits_len;
	input [2:0] io_sources_26_bits_size;
	input [1:0] io_sources_26_bits_burst;
	input io_sources_26_bits_lock;
	input [3:0] io_sources_26_bits_cache;
	input [2:0] io_sources_26_bits_prot;
	input [3:0] io_sources_26_bits_qos;
	input [3:0] io_sources_26_bits_region;
	output wire io_sources_27_ready;
	input io_sources_27_valid;
	input [63:0] io_sources_27_bits_addr;
	input [7:0] io_sources_27_bits_len;
	input [2:0] io_sources_27_bits_size;
	input [1:0] io_sources_27_bits_burst;
	input io_sources_27_bits_lock;
	input [3:0] io_sources_27_bits_cache;
	input [2:0] io_sources_27_bits_prot;
	input [3:0] io_sources_27_bits_qos;
	input [3:0] io_sources_27_bits_region;
	output wire io_sources_28_ready;
	input io_sources_28_valid;
	input [63:0] io_sources_28_bits_addr;
	input [7:0] io_sources_28_bits_len;
	input [2:0] io_sources_28_bits_size;
	input [1:0] io_sources_28_bits_burst;
	input io_sources_28_bits_lock;
	input [3:0] io_sources_28_bits_cache;
	input [2:0] io_sources_28_bits_prot;
	input [3:0] io_sources_28_bits_qos;
	input [3:0] io_sources_28_bits_region;
	output wire io_sources_29_ready;
	input io_sources_29_valid;
	input [63:0] io_sources_29_bits_addr;
	input [7:0] io_sources_29_bits_len;
	input [2:0] io_sources_29_bits_size;
	input [1:0] io_sources_29_bits_burst;
	input io_sources_29_bits_lock;
	input [3:0] io_sources_29_bits_cache;
	input [2:0] io_sources_29_bits_prot;
	input [3:0] io_sources_29_bits_qos;
	input [3:0] io_sources_29_bits_region;
	output wire io_sources_30_ready;
	input io_sources_30_valid;
	input [63:0] io_sources_30_bits_addr;
	input [7:0] io_sources_30_bits_len;
	input [2:0] io_sources_30_bits_size;
	input [1:0] io_sources_30_bits_burst;
	input io_sources_30_bits_lock;
	input [3:0] io_sources_30_bits_cache;
	input [2:0] io_sources_30_bits_prot;
	input [3:0] io_sources_30_bits_qos;
	input [3:0] io_sources_30_bits_region;
	output wire io_sources_31_ready;
	input io_sources_31_valid;
	input [63:0] io_sources_31_bits_addr;
	input [7:0] io_sources_31_bits_len;
	input [2:0] io_sources_31_bits_size;
	input [1:0] io_sources_31_bits_burst;
	input io_sources_31_bits_lock;
	input [3:0] io_sources_31_bits_cache;
	input [2:0] io_sources_31_bits_prot;
	input [3:0] io_sources_31_bits_qos;
	input [3:0] io_sources_31_bits_region;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [4:0] io_sink_bits_id;
	output wire [63:0] io_sink_bits_addr;
	output wire [7:0] io_sink_bits_len;
	output wire [2:0] io_sink_bits_size;
	output wire [1:0] io_sink_bits_burst;
	output wire io_sink_bits_lock;
	output wire [3:0] io_sink_bits_cache;
	output wire [2:0] io_sink_bits_prot;
	output wire [3:0] io_sink_bits_qos;
	output wire [3:0] io_sink_bits_region;
	input io_select_ready;
	output wire io_select_valid;
	output wire [4:0] io_select_bits;
	wire sourceReady;
	wire [159:0] _GEN = 160'hffbbcdeb38bdab49ca307b9ac5a928398a418820;
	reg [4:0] chooser_lastChoice;
	wire _chooser_rrChoice_T_4 = (chooser_lastChoice == 5'h00) & io_sources_1_valid;
	wire _chooser_rrChoice_T_6 = (chooser_lastChoice < 5'h02) & io_sources_2_valid;
	wire _chooser_rrChoice_T_8 = (chooser_lastChoice < 5'h03) & io_sources_3_valid;
	wire _chooser_rrChoice_T_10 = (chooser_lastChoice < 5'h04) & io_sources_4_valid;
	wire _chooser_rrChoice_T_12 = (chooser_lastChoice < 5'h05) & io_sources_5_valid;
	wire _chooser_rrChoice_T_14 = (chooser_lastChoice < 5'h06) & io_sources_6_valid;
	wire _chooser_rrChoice_T_16 = (chooser_lastChoice < 5'h07) & io_sources_7_valid;
	wire _chooser_rrChoice_T_18 = (chooser_lastChoice < 5'h08) & io_sources_8_valid;
	wire _chooser_rrChoice_T_20 = (chooser_lastChoice < 5'h09) & io_sources_9_valid;
	wire _chooser_rrChoice_T_22 = (chooser_lastChoice < 5'h0a) & io_sources_10_valid;
	wire _chooser_rrChoice_T_24 = (chooser_lastChoice < 5'h0b) & io_sources_11_valid;
	wire _chooser_rrChoice_T_26 = (chooser_lastChoice < 5'h0c) & io_sources_12_valid;
	wire _chooser_rrChoice_T_28 = (chooser_lastChoice < 5'h0d) & io_sources_13_valid;
	wire _chooser_rrChoice_T_30 = (chooser_lastChoice < 5'h0e) & io_sources_14_valid;
	wire _chooser_rrChoice_T_32 = (chooser_lastChoice < 5'h0f) & io_sources_15_valid;
	wire _chooser_rrChoice_T_34 = ~chooser_lastChoice[4] & io_sources_16_valid;
	wire _chooser_rrChoice_T_36 = (chooser_lastChoice < 5'h11) & io_sources_17_valid;
	wire _chooser_rrChoice_T_38 = (chooser_lastChoice < 5'h12) & io_sources_18_valid;
	wire _chooser_rrChoice_T_40 = (chooser_lastChoice < 5'h13) & io_sources_19_valid;
	wire _chooser_rrChoice_T_42 = (chooser_lastChoice < 5'h14) & io_sources_20_valid;
	wire _chooser_rrChoice_T_44 = (chooser_lastChoice < 5'h15) & io_sources_21_valid;
	wire _chooser_rrChoice_T_46 = (chooser_lastChoice < 5'h16) & io_sources_22_valid;
	wire _chooser_rrChoice_T_48 = (chooser_lastChoice < 5'h17) & io_sources_23_valid;
	wire _chooser_rrChoice_T_50 = (chooser_lastChoice[4:3] != 2'h3) & io_sources_24_valid;
	wire _chooser_rrChoice_T_52 = (chooser_lastChoice < 5'h19) & io_sources_25_valid;
	wire _chooser_rrChoice_T_54 = (chooser_lastChoice < 5'h1a) & io_sources_26_valid;
	wire _chooser_rrChoice_T_56 = (chooser_lastChoice < 5'h1b) & io_sources_27_valid;
	wire _chooser_rrChoice_T_58 = (chooser_lastChoice[4:2] != 3'h7) & io_sources_28_valid;
	wire _chooser_rrChoice_T_60 = (chooser_lastChoice < 5'h1d) & io_sources_29_valid;
	wire [4:0] _chooser_rrChoice_T_65 = {4'hf, ~((chooser_lastChoice[4:1] != 4'hf) & io_sources_30_valid)};
	wire [4:0] chooser_rrChoice = (&chooser_lastChoice ? 5'h00 : (_chooser_rrChoice_T_4 ? 5'h01 : (_chooser_rrChoice_T_6 ? 5'h02 : (_chooser_rrChoice_T_8 ? 5'h03 : (_chooser_rrChoice_T_10 ? 5'h04 : (_chooser_rrChoice_T_12 ? 5'h05 : (_chooser_rrChoice_T_14 ? 5'h06 : (_chooser_rrChoice_T_16 ? 5'h07 : (_chooser_rrChoice_T_18 ? 5'h08 : (_chooser_rrChoice_T_20 ? 5'h09 : (_chooser_rrChoice_T_22 ? 5'h0a : (_chooser_rrChoice_T_24 ? 5'h0b : (_chooser_rrChoice_T_26 ? 5'h0c : (_chooser_rrChoice_T_28 ? 5'h0d : (_chooser_rrChoice_T_30 ? 5'h0e : (_chooser_rrChoice_T_32 ? 5'h0f : (_chooser_rrChoice_T_34 ? 5'h10 : (_chooser_rrChoice_T_36 ? 5'h11 : (_chooser_rrChoice_T_38 ? 5'h12 : (_chooser_rrChoice_T_40 ? 5'h13 : (_chooser_rrChoice_T_42 ? 5'h14 : (_chooser_rrChoice_T_44 ? 5'h15 : (_chooser_rrChoice_T_46 ? 5'h16 : (_chooser_rrChoice_T_48 ? 5'h17 : (_chooser_rrChoice_T_50 ? 5'h18 : (_chooser_rrChoice_T_52 ? 5'h19 : (_chooser_rrChoice_T_54 ? 5'h1a : (_chooser_rrChoice_T_56 ? 5'h1b : (_chooser_rrChoice_T_58 ? 5'h1c : (_chooser_rrChoice_T_60 ? 5'h1d : _chooser_rrChoice_T_65))))))))))))))))))))))))))))));
	wire [4:0] chooser_priorityChoice = (io_sources_0_valid ? 5'h00 : (io_sources_1_valid ? 5'h01 : (io_sources_2_valid ? 5'h02 : (io_sources_3_valid ? 5'h03 : (io_sources_4_valid ? 5'h04 : (io_sources_5_valid ? 5'h05 : (io_sources_6_valid ? 5'h06 : (io_sources_7_valid ? 5'h07 : (io_sources_8_valid ? 5'h08 : (io_sources_9_valid ? 5'h09 : (io_sources_10_valid ? 5'h0a : (io_sources_11_valid ? 5'h0b : (io_sources_12_valid ? 5'h0c : (io_sources_13_valid ? 5'h0d : (io_sources_14_valid ? 5'h0e : (io_sources_15_valid ? 5'h0f : (io_sources_16_valid ? 5'h10 : (io_sources_17_valid ? 5'h11 : (io_sources_18_valid ? 5'h12 : (io_sources_19_valid ? 5'h13 : (io_sources_20_valid ? 5'h14 : (io_sources_21_valid ? 5'h15 : (io_sources_22_valid ? 5'h16 : (io_sources_23_valid ? 5'h17 : (io_sources_24_valid ? 5'h18 : (io_sources_25_valid ? 5'h19 : (io_sources_26_valid ? 5'h1a : (io_sources_27_valid ? 5'h1b : (io_sources_28_valid ? 5'h1c : (io_sources_29_valid ? 5'h1d : {4'hf, ~io_sources_30_valid}))))))))))))))))))))))))))))));
	wire [31:0] _GEN_0 = {io_sources_31_valid, io_sources_30_valid, io_sources_29_valid, io_sources_28_valid, io_sources_27_valid, io_sources_26_valid, io_sources_25_valid, io_sources_24_valid, io_sources_23_valid, io_sources_22_valid, io_sources_21_valid, io_sources_20_valid, io_sources_19_valid, io_sources_18_valid, io_sources_17_valid, io_sources_16_valid, io_sources_15_valid, io_sources_14_valid, io_sources_13_valid, io_sources_12_valid, io_sources_11_valid, io_sources_10_valid, io_sources_9_valid, io_sources_8_valid, io_sources_7_valid, io_sources_6_valid, io_sources_5_valid, io_sources_4_valid, io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [4:0] io_select_bits_0 = (_GEN_0[chooser_rrChoice] ? chooser_rrChoice : chooser_priorityChoice);
	wire [2047:0] _GEN_1 = {io_sources_31_bits_addr, io_sources_30_bits_addr, io_sources_29_bits_addr, io_sources_28_bits_addr, io_sources_27_bits_addr, io_sources_26_bits_addr, io_sources_25_bits_addr, io_sources_24_bits_addr, io_sources_23_bits_addr, io_sources_22_bits_addr, io_sources_21_bits_addr, io_sources_20_bits_addr, io_sources_19_bits_addr, io_sources_18_bits_addr, io_sources_17_bits_addr, io_sources_16_bits_addr, io_sources_15_bits_addr, io_sources_14_bits_addr, io_sources_13_bits_addr, io_sources_12_bits_addr, io_sources_11_bits_addr, io_sources_10_bits_addr, io_sources_9_bits_addr, io_sources_8_bits_addr, io_sources_7_bits_addr, io_sources_6_bits_addr, io_sources_5_bits_addr, io_sources_4_bits_addr, io_sources_3_bits_addr, io_sources_2_bits_addr, io_sources_1_bits_addr, io_sources_0_bits_addr};
	wire [255:0] _GEN_2 = {io_sources_31_bits_len, io_sources_30_bits_len, io_sources_29_bits_len, io_sources_28_bits_len, io_sources_27_bits_len, io_sources_26_bits_len, io_sources_25_bits_len, io_sources_24_bits_len, io_sources_23_bits_len, io_sources_22_bits_len, io_sources_21_bits_len, io_sources_20_bits_len, io_sources_19_bits_len, io_sources_18_bits_len, io_sources_17_bits_len, io_sources_16_bits_len, io_sources_15_bits_len, io_sources_14_bits_len, io_sources_13_bits_len, io_sources_12_bits_len, io_sources_11_bits_len, io_sources_10_bits_len, io_sources_9_bits_len, io_sources_8_bits_len, io_sources_7_bits_len, io_sources_6_bits_len, io_sources_5_bits_len, io_sources_4_bits_len, io_sources_3_bits_len, io_sources_2_bits_len, io_sources_1_bits_len, io_sources_0_bits_len};
	wire [95:0] _GEN_3 = {io_sources_31_bits_size, io_sources_30_bits_size, io_sources_29_bits_size, io_sources_28_bits_size, io_sources_27_bits_size, io_sources_26_bits_size, io_sources_25_bits_size, io_sources_24_bits_size, io_sources_23_bits_size, io_sources_22_bits_size, io_sources_21_bits_size, io_sources_20_bits_size, io_sources_19_bits_size, io_sources_18_bits_size, io_sources_17_bits_size, io_sources_16_bits_size, io_sources_15_bits_size, io_sources_14_bits_size, io_sources_13_bits_size, io_sources_12_bits_size, io_sources_11_bits_size, io_sources_10_bits_size, io_sources_9_bits_size, io_sources_8_bits_size, io_sources_7_bits_size, io_sources_6_bits_size, io_sources_5_bits_size, io_sources_4_bits_size, io_sources_3_bits_size, io_sources_2_bits_size, io_sources_1_bits_size, io_sources_0_bits_size};
	wire [63:0] _GEN_4 = {io_sources_31_bits_burst, io_sources_30_bits_burst, io_sources_29_bits_burst, io_sources_28_bits_burst, io_sources_27_bits_burst, io_sources_26_bits_burst, io_sources_25_bits_burst, io_sources_24_bits_burst, io_sources_23_bits_burst, io_sources_22_bits_burst, io_sources_21_bits_burst, io_sources_20_bits_burst, io_sources_19_bits_burst, io_sources_18_bits_burst, io_sources_17_bits_burst, io_sources_16_bits_burst, io_sources_15_bits_burst, io_sources_14_bits_burst, io_sources_13_bits_burst, io_sources_12_bits_burst, io_sources_11_bits_burst, io_sources_10_bits_burst, io_sources_9_bits_burst, io_sources_8_bits_burst, io_sources_7_bits_burst, io_sources_6_bits_burst, io_sources_5_bits_burst, io_sources_4_bits_burst, io_sources_3_bits_burst, io_sources_2_bits_burst, io_sources_1_bits_burst, io_sources_0_bits_burst};
	wire [31:0] _GEN_5 = {io_sources_31_bits_lock, io_sources_30_bits_lock, io_sources_29_bits_lock, io_sources_28_bits_lock, io_sources_27_bits_lock, io_sources_26_bits_lock, io_sources_25_bits_lock, io_sources_24_bits_lock, io_sources_23_bits_lock, io_sources_22_bits_lock, io_sources_21_bits_lock, io_sources_20_bits_lock, io_sources_19_bits_lock, io_sources_18_bits_lock, io_sources_17_bits_lock, io_sources_16_bits_lock, io_sources_15_bits_lock, io_sources_14_bits_lock, io_sources_13_bits_lock, io_sources_12_bits_lock, io_sources_11_bits_lock, io_sources_10_bits_lock, io_sources_9_bits_lock, io_sources_8_bits_lock, io_sources_7_bits_lock, io_sources_6_bits_lock, io_sources_5_bits_lock, io_sources_4_bits_lock, io_sources_3_bits_lock, io_sources_2_bits_lock, io_sources_1_bits_lock, io_sources_0_bits_lock};
	wire [127:0] _GEN_6 = {io_sources_31_bits_cache, io_sources_30_bits_cache, io_sources_29_bits_cache, io_sources_28_bits_cache, io_sources_27_bits_cache, io_sources_26_bits_cache, io_sources_25_bits_cache, io_sources_24_bits_cache, io_sources_23_bits_cache, io_sources_22_bits_cache, io_sources_21_bits_cache, io_sources_20_bits_cache, io_sources_19_bits_cache, io_sources_18_bits_cache, io_sources_17_bits_cache, io_sources_16_bits_cache, io_sources_15_bits_cache, io_sources_14_bits_cache, io_sources_13_bits_cache, io_sources_12_bits_cache, io_sources_11_bits_cache, io_sources_10_bits_cache, io_sources_9_bits_cache, io_sources_8_bits_cache, io_sources_7_bits_cache, io_sources_6_bits_cache, io_sources_5_bits_cache, io_sources_4_bits_cache, io_sources_3_bits_cache, io_sources_2_bits_cache, io_sources_1_bits_cache, io_sources_0_bits_cache};
	wire [95:0] _GEN_7 = {io_sources_31_bits_prot, io_sources_30_bits_prot, io_sources_29_bits_prot, io_sources_28_bits_prot, io_sources_27_bits_prot, io_sources_26_bits_prot, io_sources_25_bits_prot, io_sources_24_bits_prot, io_sources_23_bits_prot, io_sources_22_bits_prot, io_sources_21_bits_prot, io_sources_20_bits_prot, io_sources_19_bits_prot, io_sources_18_bits_prot, io_sources_17_bits_prot, io_sources_16_bits_prot, io_sources_15_bits_prot, io_sources_14_bits_prot, io_sources_13_bits_prot, io_sources_12_bits_prot, io_sources_11_bits_prot, io_sources_10_bits_prot, io_sources_9_bits_prot, io_sources_8_bits_prot, io_sources_7_bits_prot, io_sources_6_bits_prot, io_sources_5_bits_prot, io_sources_4_bits_prot, io_sources_3_bits_prot, io_sources_2_bits_prot, io_sources_1_bits_prot, io_sources_0_bits_prot};
	wire [127:0] _GEN_8 = {io_sources_31_bits_qos, io_sources_30_bits_qos, io_sources_29_bits_qos, io_sources_28_bits_qos, io_sources_27_bits_qos, io_sources_26_bits_qos, io_sources_25_bits_qos, io_sources_24_bits_qos, io_sources_23_bits_qos, io_sources_22_bits_qos, io_sources_21_bits_qos, io_sources_20_bits_qos, io_sources_19_bits_qos, io_sources_18_bits_qos, io_sources_17_bits_qos, io_sources_16_bits_qos, io_sources_15_bits_qos, io_sources_14_bits_qos, io_sources_13_bits_qos, io_sources_12_bits_qos, io_sources_11_bits_qos, io_sources_10_bits_qos, io_sources_9_bits_qos, io_sources_8_bits_qos, io_sources_7_bits_qos, io_sources_6_bits_qos, io_sources_5_bits_qos, io_sources_4_bits_qos, io_sources_3_bits_qos, io_sources_2_bits_qos, io_sources_1_bits_qos, io_sources_0_bits_qos};
	wire [127:0] _GEN_9 = {io_sources_31_bits_region, io_sources_30_bits_region, io_sources_29_bits_region, io_sources_28_bits_region, io_sources_27_bits_region, io_sources_26_bits_region, io_sources_25_bits_region, io_sources_24_bits_region, io_sources_23_bits_region, io_sources_22_bits_region, io_sources_21_bits_region, io_sources_20_bits_region, io_sources_19_bits_region, io_sources_18_bits_region, io_sources_17_bits_region, io_sources_16_bits_region, io_sources_15_bits_region, io_sources_14_bits_region, io_sources_13_bits_region, io_sources_12_bits_region, io_sources_11_bits_region, io_sources_10_bits_region, io_sources_9_bits_region, io_sources_8_bits_region, io_sources_7_bits_region, io_sources_6_bits_region, io_sources_5_bits_region, io_sources_4_bits_region, io_sources_3_bits_region, io_sources_2_bits_region, io_sources_1_bits_region, io_sources_0_bits_region};
	reg sinkSent;
	reg selectSent;
	assign sourceReady = (sinkSent | io_sink_ready) & (selectSent | io_select_ready);
	always @(posedge clock)
		if (reset) begin
			chooser_lastChoice <= 5'h00;
			sinkSent <= 1'h0;
			selectSent <= 1'h0;
		end
		else begin
			if (_GEN_0[io_select_bits_0] & sourceReady) begin
				if (_GEN_0[chooser_rrChoice]) begin
					if (&chooser_lastChoice)
						chooser_lastChoice <= 5'h00;
					else if (_chooser_rrChoice_T_4)
						chooser_lastChoice <= 5'h01;
					else if (_chooser_rrChoice_T_6)
						chooser_lastChoice <= 5'h02;
					else if (_chooser_rrChoice_T_8)
						chooser_lastChoice <= 5'h03;
					else if (_chooser_rrChoice_T_10)
						chooser_lastChoice <= 5'h04;
					else if (_chooser_rrChoice_T_12)
						chooser_lastChoice <= 5'h05;
					else if (_chooser_rrChoice_T_14)
						chooser_lastChoice <= 5'h06;
					else if (_chooser_rrChoice_T_16)
						chooser_lastChoice <= 5'h07;
					else if (_chooser_rrChoice_T_18)
						chooser_lastChoice <= 5'h08;
					else if (_chooser_rrChoice_T_20)
						chooser_lastChoice <= 5'h09;
					else if (_chooser_rrChoice_T_22)
						chooser_lastChoice <= 5'h0a;
					else if (_chooser_rrChoice_T_24)
						chooser_lastChoice <= 5'h0b;
					else if (_chooser_rrChoice_T_26)
						chooser_lastChoice <= 5'h0c;
					else if (_chooser_rrChoice_T_28)
						chooser_lastChoice <= 5'h0d;
					else if (_chooser_rrChoice_T_30)
						chooser_lastChoice <= 5'h0e;
					else if (_chooser_rrChoice_T_32)
						chooser_lastChoice <= 5'h0f;
					else if (_chooser_rrChoice_T_34)
						chooser_lastChoice <= 5'h10;
					else if (_chooser_rrChoice_T_36)
						chooser_lastChoice <= 5'h11;
					else if (_chooser_rrChoice_T_38)
						chooser_lastChoice <= 5'h12;
					else if (_chooser_rrChoice_T_40)
						chooser_lastChoice <= 5'h13;
					else if (_chooser_rrChoice_T_42)
						chooser_lastChoice <= 5'h14;
					else if (_chooser_rrChoice_T_44)
						chooser_lastChoice <= 5'h15;
					else if (_chooser_rrChoice_T_46)
						chooser_lastChoice <= 5'h16;
					else if (_chooser_rrChoice_T_48)
						chooser_lastChoice <= 5'h17;
					else if (_chooser_rrChoice_T_50)
						chooser_lastChoice <= 5'h18;
					else if (_chooser_rrChoice_T_52)
						chooser_lastChoice <= 5'h19;
					else if (_chooser_rrChoice_T_54)
						chooser_lastChoice <= 5'h1a;
					else if (_chooser_rrChoice_T_56)
						chooser_lastChoice <= 5'h1b;
					else if (_chooser_rrChoice_T_58)
						chooser_lastChoice <= 5'h1c;
					else if (_chooser_rrChoice_T_60)
						chooser_lastChoice <= 5'h1d;
					else
						chooser_lastChoice <= _chooser_rrChoice_T_65;
				end
				else
					chooser_lastChoice <= chooser_priorityChoice;
			end
			sinkSent <= ((io_sink_ready | sinkSent) & _GEN_0[io_select_bits_0]) & ~sourceReady;
			selectSent <= ((io_select_ready | selectSent) & _GEN_0[io_select_bits_0]) & ~sourceReady;
		end
	assign io_sources_0_ready = sourceReady & (io_select_bits_0 == 5'h00);
	assign io_sources_1_ready = sourceReady & (io_select_bits_0 == 5'h01);
	assign io_sources_2_ready = sourceReady & (io_select_bits_0 == 5'h02);
	assign io_sources_3_ready = sourceReady & (io_select_bits_0 == 5'h03);
	assign io_sources_4_ready = sourceReady & (io_select_bits_0 == 5'h04);
	assign io_sources_5_ready = sourceReady & (io_select_bits_0 == 5'h05);
	assign io_sources_6_ready = sourceReady & (io_select_bits_0 == 5'h06);
	assign io_sources_7_ready = sourceReady & (io_select_bits_0 == 5'h07);
	assign io_sources_8_ready = sourceReady & (io_select_bits_0 == 5'h08);
	assign io_sources_9_ready = sourceReady & (io_select_bits_0 == 5'h09);
	assign io_sources_10_ready = sourceReady & (io_select_bits_0 == 5'h0a);
	assign io_sources_11_ready = sourceReady & (io_select_bits_0 == 5'h0b);
	assign io_sources_12_ready = sourceReady & (io_select_bits_0 == 5'h0c);
	assign io_sources_13_ready = sourceReady & (io_select_bits_0 == 5'h0d);
	assign io_sources_14_ready = sourceReady & (io_select_bits_0 == 5'h0e);
	assign io_sources_15_ready = sourceReady & (io_select_bits_0 == 5'h0f);
	assign io_sources_16_ready = sourceReady & (io_select_bits_0 == 5'h10);
	assign io_sources_17_ready = sourceReady & (io_select_bits_0 == 5'h11);
	assign io_sources_18_ready = sourceReady & (io_select_bits_0 == 5'h12);
	assign io_sources_19_ready = sourceReady & (io_select_bits_0 == 5'h13);
	assign io_sources_20_ready = sourceReady & (io_select_bits_0 == 5'h14);
	assign io_sources_21_ready = sourceReady & (io_select_bits_0 == 5'h15);
	assign io_sources_22_ready = sourceReady & (io_select_bits_0 == 5'h16);
	assign io_sources_23_ready = sourceReady & (io_select_bits_0 == 5'h17);
	assign io_sources_24_ready = sourceReady & (io_select_bits_0 == 5'h18);
	assign io_sources_25_ready = sourceReady & (io_select_bits_0 == 5'h19);
	assign io_sources_26_ready = sourceReady & (io_select_bits_0 == 5'h1a);
	assign io_sources_27_ready = sourceReady & (io_select_bits_0 == 5'h1b);
	assign io_sources_28_ready = sourceReady & (io_select_bits_0 == 5'h1c);
	assign io_sources_29_ready = sourceReady & (io_select_bits_0 == 5'h1d);
	assign io_sources_30_ready = sourceReady & (io_select_bits_0 == 5'h1e);
	assign io_sources_31_ready = sourceReady & (&io_select_bits_0);
	assign io_sink_valid = _GEN_0[io_select_bits_0] & ~sinkSent;
	assign io_sink_bits_id = _GEN[io_select_bits_0 * 5+:5];
	assign io_sink_bits_addr = _GEN_1[io_select_bits_0 * 64+:64];
	assign io_sink_bits_len = _GEN_2[io_select_bits_0 * 8+:8];
	assign io_sink_bits_size = _GEN_3[io_select_bits_0 * 3+:3];
	assign io_sink_bits_burst = _GEN_4[io_select_bits_0 * 2+:2];
	assign io_sink_bits_lock = _GEN_5[io_select_bits_0];
	assign io_sink_bits_cache = _GEN_6[io_select_bits_0 * 4+:4];
	assign io_sink_bits_prot = _GEN_7[io_select_bits_0 * 3+:3];
	assign io_sink_bits_qos = _GEN_8[io_select_bits_0 * 4+:4];
	assign io_sink_bits_region = _GEN_9[io_select_bits_0 * 4+:4];
	assign io_select_valid = _GEN_0[io_select_bits_0] & ~selectSent;
	assign io_select_bits = io_select_bits_0;
endmodule
module elasticDemux_9 (
	io_source_ready,
	io_source_valid,
	io_source_bits_data,
	io_source_bits_resp,
	io_source_bits_last,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_data,
	io_sinks_0_bits_resp,
	io_sinks_0_bits_last,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_data,
	io_sinks_1_bits_resp,
	io_sinks_1_bits_last,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_2_bits_data,
	io_sinks_2_bits_resp,
	io_sinks_2_bits_last,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_3_bits_data,
	io_sinks_3_bits_resp,
	io_sinks_3_bits_last,
	io_sinks_4_ready,
	io_sinks_4_valid,
	io_sinks_4_bits_data,
	io_sinks_4_bits_resp,
	io_sinks_4_bits_last,
	io_sinks_5_ready,
	io_sinks_5_valid,
	io_sinks_5_bits_data,
	io_sinks_5_bits_resp,
	io_sinks_5_bits_last,
	io_sinks_6_ready,
	io_sinks_6_valid,
	io_sinks_6_bits_data,
	io_sinks_6_bits_resp,
	io_sinks_6_bits_last,
	io_sinks_7_ready,
	io_sinks_7_valid,
	io_sinks_7_bits_data,
	io_sinks_7_bits_resp,
	io_sinks_7_bits_last,
	io_sinks_8_ready,
	io_sinks_8_valid,
	io_sinks_8_bits_data,
	io_sinks_8_bits_resp,
	io_sinks_8_bits_last,
	io_sinks_9_ready,
	io_sinks_9_valid,
	io_sinks_9_bits_data,
	io_sinks_9_bits_resp,
	io_sinks_9_bits_last,
	io_sinks_10_ready,
	io_sinks_10_valid,
	io_sinks_10_bits_data,
	io_sinks_10_bits_resp,
	io_sinks_10_bits_last,
	io_sinks_11_ready,
	io_sinks_11_valid,
	io_sinks_11_bits_data,
	io_sinks_11_bits_resp,
	io_sinks_11_bits_last,
	io_sinks_12_ready,
	io_sinks_12_valid,
	io_sinks_12_bits_data,
	io_sinks_12_bits_resp,
	io_sinks_12_bits_last,
	io_sinks_13_ready,
	io_sinks_13_valid,
	io_sinks_13_bits_data,
	io_sinks_13_bits_resp,
	io_sinks_13_bits_last,
	io_sinks_14_ready,
	io_sinks_14_valid,
	io_sinks_14_bits_data,
	io_sinks_14_bits_resp,
	io_sinks_14_bits_last,
	io_sinks_15_ready,
	io_sinks_15_valid,
	io_sinks_15_bits_data,
	io_sinks_15_bits_resp,
	io_sinks_15_bits_last,
	io_sinks_16_ready,
	io_sinks_16_valid,
	io_sinks_16_bits_data,
	io_sinks_16_bits_resp,
	io_sinks_16_bits_last,
	io_sinks_17_ready,
	io_sinks_17_valid,
	io_sinks_17_bits_data,
	io_sinks_17_bits_resp,
	io_sinks_17_bits_last,
	io_sinks_18_ready,
	io_sinks_18_valid,
	io_sinks_18_bits_data,
	io_sinks_18_bits_resp,
	io_sinks_18_bits_last,
	io_sinks_19_ready,
	io_sinks_19_valid,
	io_sinks_19_bits_data,
	io_sinks_19_bits_resp,
	io_sinks_19_bits_last,
	io_sinks_20_ready,
	io_sinks_20_valid,
	io_sinks_20_bits_data,
	io_sinks_20_bits_resp,
	io_sinks_20_bits_last,
	io_sinks_21_ready,
	io_sinks_21_valid,
	io_sinks_21_bits_data,
	io_sinks_21_bits_resp,
	io_sinks_21_bits_last,
	io_sinks_22_ready,
	io_sinks_22_valid,
	io_sinks_22_bits_data,
	io_sinks_22_bits_resp,
	io_sinks_22_bits_last,
	io_sinks_23_ready,
	io_sinks_23_valid,
	io_sinks_23_bits_data,
	io_sinks_23_bits_resp,
	io_sinks_23_bits_last,
	io_sinks_24_ready,
	io_sinks_24_valid,
	io_sinks_24_bits_data,
	io_sinks_24_bits_resp,
	io_sinks_24_bits_last,
	io_sinks_25_ready,
	io_sinks_25_valid,
	io_sinks_25_bits_data,
	io_sinks_25_bits_resp,
	io_sinks_25_bits_last,
	io_sinks_26_ready,
	io_sinks_26_valid,
	io_sinks_26_bits_data,
	io_sinks_26_bits_resp,
	io_sinks_26_bits_last,
	io_sinks_27_ready,
	io_sinks_27_valid,
	io_sinks_27_bits_data,
	io_sinks_27_bits_resp,
	io_sinks_27_bits_last,
	io_sinks_28_ready,
	io_sinks_28_valid,
	io_sinks_28_bits_data,
	io_sinks_28_bits_resp,
	io_sinks_28_bits_last,
	io_sinks_29_ready,
	io_sinks_29_valid,
	io_sinks_29_bits_data,
	io_sinks_29_bits_resp,
	io_sinks_29_bits_last,
	io_sinks_30_ready,
	io_sinks_30_valid,
	io_sinks_30_bits_data,
	io_sinks_30_bits_resp,
	io_sinks_30_bits_last,
	io_sinks_31_ready,
	io_sinks_31_valid,
	io_sinks_31_bits_data,
	io_sinks_31_bits_resp,
	io_sinks_31_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [31:0] io_source_bits_data;
	input [1:0] io_source_bits_resp;
	input io_source_bits_last;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [31:0] io_sinks_0_bits_data;
	output wire [1:0] io_sinks_0_bits_resp;
	output wire io_sinks_0_bits_last;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [31:0] io_sinks_1_bits_data;
	output wire [1:0] io_sinks_1_bits_resp;
	output wire io_sinks_1_bits_last;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	output wire [31:0] io_sinks_2_bits_data;
	output wire [1:0] io_sinks_2_bits_resp;
	output wire io_sinks_2_bits_last;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire [31:0] io_sinks_3_bits_data;
	output wire [1:0] io_sinks_3_bits_resp;
	output wire io_sinks_3_bits_last;
	input io_sinks_4_ready;
	output wire io_sinks_4_valid;
	output wire [31:0] io_sinks_4_bits_data;
	output wire [1:0] io_sinks_4_bits_resp;
	output wire io_sinks_4_bits_last;
	input io_sinks_5_ready;
	output wire io_sinks_5_valid;
	output wire [31:0] io_sinks_5_bits_data;
	output wire [1:0] io_sinks_5_bits_resp;
	output wire io_sinks_5_bits_last;
	input io_sinks_6_ready;
	output wire io_sinks_6_valid;
	output wire [31:0] io_sinks_6_bits_data;
	output wire [1:0] io_sinks_6_bits_resp;
	output wire io_sinks_6_bits_last;
	input io_sinks_7_ready;
	output wire io_sinks_7_valid;
	output wire [31:0] io_sinks_7_bits_data;
	output wire [1:0] io_sinks_7_bits_resp;
	output wire io_sinks_7_bits_last;
	input io_sinks_8_ready;
	output wire io_sinks_8_valid;
	output wire [31:0] io_sinks_8_bits_data;
	output wire [1:0] io_sinks_8_bits_resp;
	output wire io_sinks_8_bits_last;
	input io_sinks_9_ready;
	output wire io_sinks_9_valid;
	output wire [31:0] io_sinks_9_bits_data;
	output wire [1:0] io_sinks_9_bits_resp;
	output wire io_sinks_9_bits_last;
	input io_sinks_10_ready;
	output wire io_sinks_10_valid;
	output wire [31:0] io_sinks_10_bits_data;
	output wire [1:0] io_sinks_10_bits_resp;
	output wire io_sinks_10_bits_last;
	input io_sinks_11_ready;
	output wire io_sinks_11_valid;
	output wire [31:0] io_sinks_11_bits_data;
	output wire [1:0] io_sinks_11_bits_resp;
	output wire io_sinks_11_bits_last;
	input io_sinks_12_ready;
	output wire io_sinks_12_valid;
	output wire [31:0] io_sinks_12_bits_data;
	output wire [1:0] io_sinks_12_bits_resp;
	output wire io_sinks_12_bits_last;
	input io_sinks_13_ready;
	output wire io_sinks_13_valid;
	output wire [31:0] io_sinks_13_bits_data;
	output wire [1:0] io_sinks_13_bits_resp;
	output wire io_sinks_13_bits_last;
	input io_sinks_14_ready;
	output wire io_sinks_14_valid;
	output wire [31:0] io_sinks_14_bits_data;
	output wire [1:0] io_sinks_14_bits_resp;
	output wire io_sinks_14_bits_last;
	input io_sinks_15_ready;
	output wire io_sinks_15_valid;
	output wire [31:0] io_sinks_15_bits_data;
	output wire [1:0] io_sinks_15_bits_resp;
	output wire io_sinks_15_bits_last;
	input io_sinks_16_ready;
	output wire io_sinks_16_valid;
	output wire [31:0] io_sinks_16_bits_data;
	output wire [1:0] io_sinks_16_bits_resp;
	output wire io_sinks_16_bits_last;
	input io_sinks_17_ready;
	output wire io_sinks_17_valid;
	output wire [31:0] io_sinks_17_bits_data;
	output wire [1:0] io_sinks_17_bits_resp;
	output wire io_sinks_17_bits_last;
	input io_sinks_18_ready;
	output wire io_sinks_18_valid;
	output wire [31:0] io_sinks_18_bits_data;
	output wire [1:0] io_sinks_18_bits_resp;
	output wire io_sinks_18_bits_last;
	input io_sinks_19_ready;
	output wire io_sinks_19_valid;
	output wire [31:0] io_sinks_19_bits_data;
	output wire [1:0] io_sinks_19_bits_resp;
	output wire io_sinks_19_bits_last;
	input io_sinks_20_ready;
	output wire io_sinks_20_valid;
	output wire [31:0] io_sinks_20_bits_data;
	output wire [1:0] io_sinks_20_bits_resp;
	output wire io_sinks_20_bits_last;
	input io_sinks_21_ready;
	output wire io_sinks_21_valid;
	output wire [31:0] io_sinks_21_bits_data;
	output wire [1:0] io_sinks_21_bits_resp;
	output wire io_sinks_21_bits_last;
	input io_sinks_22_ready;
	output wire io_sinks_22_valid;
	output wire [31:0] io_sinks_22_bits_data;
	output wire [1:0] io_sinks_22_bits_resp;
	output wire io_sinks_22_bits_last;
	input io_sinks_23_ready;
	output wire io_sinks_23_valid;
	output wire [31:0] io_sinks_23_bits_data;
	output wire [1:0] io_sinks_23_bits_resp;
	output wire io_sinks_23_bits_last;
	input io_sinks_24_ready;
	output wire io_sinks_24_valid;
	output wire [31:0] io_sinks_24_bits_data;
	output wire [1:0] io_sinks_24_bits_resp;
	output wire io_sinks_24_bits_last;
	input io_sinks_25_ready;
	output wire io_sinks_25_valid;
	output wire [31:0] io_sinks_25_bits_data;
	output wire [1:0] io_sinks_25_bits_resp;
	output wire io_sinks_25_bits_last;
	input io_sinks_26_ready;
	output wire io_sinks_26_valid;
	output wire [31:0] io_sinks_26_bits_data;
	output wire [1:0] io_sinks_26_bits_resp;
	output wire io_sinks_26_bits_last;
	input io_sinks_27_ready;
	output wire io_sinks_27_valid;
	output wire [31:0] io_sinks_27_bits_data;
	output wire [1:0] io_sinks_27_bits_resp;
	output wire io_sinks_27_bits_last;
	input io_sinks_28_ready;
	output wire io_sinks_28_valid;
	output wire [31:0] io_sinks_28_bits_data;
	output wire [1:0] io_sinks_28_bits_resp;
	output wire io_sinks_28_bits_last;
	input io_sinks_29_ready;
	output wire io_sinks_29_valid;
	output wire [31:0] io_sinks_29_bits_data;
	output wire [1:0] io_sinks_29_bits_resp;
	output wire io_sinks_29_bits_last;
	input io_sinks_30_ready;
	output wire io_sinks_30_valid;
	output wire [31:0] io_sinks_30_bits_data;
	output wire [1:0] io_sinks_30_bits_resp;
	output wire io_sinks_30_bits_last;
	input io_sinks_31_ready;
	output wire io_sinks_31_valid;
	output wire [31:0] io_sinks_31_bits_data;
	output wire [1:0] io_sinks_31_bits_resp;
	output wire io_sinks_31_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input [4:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [31:0] _GEN = {io_sinks_31_ready, io_sinks_30_ready, io_sinks_29_ready, io_sinks_28_ready, io_sinks_27_ready, io_sinks_26_ready, io_sinks_25_ready, io_sinks_24_ready, io_sinks_23_ready, io_sinks_22_ready, io_sinks_21_ready, io_sinks_20_ready, io_sinks_19_ready, io_sinks_18_ready, io_sinks_17_ready, io_sinks_16_ready, io_sinks_15_ready, io_sinks_14_ready, io_sinks_13_ready, io_sinks_12_ready, io_sinks_11_ready, io_sinks_10_ready, io_sinks_9_ready, io_sinks_8_ready, io_sinks_7_ready, io_sinks_6_ready, io_sinks_5_ready, io_sinks_4_ready, io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 5'h00);
	assign io_sinks_0_bits_data = io_source_bits_data;
	assign io_sinks_0_bits_resp = io_source_bits_resp;
	assign io_sinks_0_bits_last = io_source_bits_last;
	assign io_sinks_1_valid = valid & (io_select_bits == 5'h01);
	assign io_sinks_1_bits_data = io_source_bits_data;
	assign io_sinks_1_bits_resp = io_source_bits_resp;
	assign io_sinks_1_bits_last = io_source_bits_last;
	assign io_sinks_2_valid = valid & (io_select_bits == 5'h02);
	assign io_sinks_2_bits_data = io_source_bits_data;
	assign io_sinks_2_bits_resp = io_source_bits_resp;
	assign io_sinks_2_bits_last = io_source_bits_last;
	assign io_sinks_3_valid = valid & (io_select_bits == 5'h03);
	assign io_sinks_3_bits_data = io_source_bits_data;
	assign io_sinks_3_bits_resp = io_source_bits_resp;
	assign io_sinks_3_bits_last = io_source_bits_last;
	assign io_sinks_4_valid = valid & (io_select_bits == 5'h04);
	assign io_sinks_4_bits_data = io_source_bits_data;
	assign io_sinks_4_bits_resp = io_source_bits_resp;
	assign io_sinks_4_bits_last = io_source_bits_last;
	assign io_sinks_5_valid = valid & (io_select_bits == 5'h05);
	assign io_sinks_5_bits_data = io_source_bits_data;
	assign io_sinks_5_bits_resp = io_source_bits_resp;
	assign io_sinks_5_bits_last = io_source_bits_last;
	assign io_sinks_6_valid = valid & (io_select_bits == 5'h06);
	assign io_sinks_6_bits_data = io_source_bits_data;
	assign io_sinks_6_bits_resp = io_source_bits_resp;
	assign io_sinks_6_bits_last = io_source_bits_last;
	assign io_sinks_7_valid = valid & (io_select_bits == 5'h07);
	assign io_sinks_7_bits_data = io_source_bits_data;
	assign io_sinks_7_bits_resp = io_source_bits_resp;
	assign io_sinks_7_bits_last = io_source_bits_last;
	assign io_sinks_8_valid = valid & (io_select_bits == 5'h08);
	assign io_sinks_8_bits_data = io_source_bits_data;
	assign io_sinks_8_bits_resp = io_source_bits_resp;
	assign io_sinks_8_bits_last = io_source_bits_last;
	assign io_sinks_9_valid = valid & (io_select_bits == 5'h09);
	assign io_sinks_9_bits_data = io_source_bits_data;
	assign io_sinks_9_bits_resp = io_source_bits_resp;
	assign io_sinks_9_bits_last = io_source_bits_last;
	assign io_sinks_10_valid = valid & (io_select_bits == 5'h0a);
	assign io_sinks_10_bits_data = io_source_bits_data;
	assign io_sinks_10_bits_resp = io_source_bits_resp;
	assign io_sinks_10_bits_last = io_source_bits_last;
	assign io_sinks_11_valid = valid & (io_select_bits == 5'h0b);
	assign io_sinks_11_bits_data = io_source_bits_data;
	assign io_sinks_11_bits_resp = io_source_bits_resp;
	assign io_sinks_11_bits_last = io_source_bits_last;
	assign io_sinks_12_valid = valid & (io_select_bits == 5'h0c);
	assign io_sinks_12_bits_data = io_source_bits_data;
	assign io_sinks_12_bits_resp = io_source_bits_resp;
	assign io_sinks_12_bits_last = io_source_bits_last;
	assign io_sinks_13_valid = valid & (io_select_bits == 5'h0d);
	assign io_sinks_13_bits_data = io_source_bits_data;
	assign io_sinks_13_bits_resp = io_source_bits_resp;
	assign io_sinks_13_bits_last = io_source_bits_last;
	assign io_sinks_14_valid = valid & (io_select_bits == 5'h0e);
	assign io_sinks_14_bits_data = io_source_bits_data;
	assign io_sinks_14_bits_resp = io_source_bits_resp;
	assign io_sinks_14_bits_last = io_source_bits_last;
	assign io_sinks_15_valid = valid & (io_select_bits == 5'h0f);
	assign io_sinks_15_bits_data = io_source_bits_data;
	assign io_sinks_15_bits_resp = io_source_bits_resp;
	assign io_sinks_15_bits_last = io_source_bits_last;
	assign io_sinks_16_valid = valid & (io_select_bits == 5'h10);
	assign io_sinks_16_bits_data = io_source_bits_data;
	assign io_sinks_16_bits_resp = io_source_bits_resp;
	assign io_sinks_16_bits_last = io_source_bits_last;
	assign io_sinks_17_valid = valid & (io_select_bits == 5'h11);
	assign io_sinks_17_bits_data = io_source_bits_data;
	assign io_sinks_17_bits_resp = io_source_bits_resp;
	assign io_sinks_17_bits_last = io_source_bits_last;
	assign io_sinks_18_valid = valid & (io_select_bits == 5'h12);
	assign io_sinks_18_bits_data = io_source_bits_data;
	assign io_sinks_18_bits_resp = io_source_bits_resp;
	assign io_sinks_18_bits_last = io_source_bits_last;
	assign io_sinks_19_valid = valid & (io_select_bits == 5'h13);
	assign io_sinks_19_bits_data = io_source_bits_data;
	assign io_sinks_19_bits_resp = io_source_bits_resp;
	assign io_sinks_19_bits_last = io_source_bits_last;
	assign io_sinks_20_valid = valid & (io_select_bits == 5'h14);
	assign io_sinks_20_bits_data = io_source_bits_data;
	assign io_sinks_20_bits_resp = io_source_bits_resp;
	assign io_sinks_20_bits_last = io_source_bits_last;
	assign io_sinks_21_valid = valid & (io_select_bits == 5'h15);
	assign io_sinks_21_bits_data = io_source_bits_data;
	assign io_sinks_21_bits_resp = io_source_bits_resp;
	assign io_sinks_21_bits_last = io_source_bits_last;
	assign io_sinks_22_valid = valid & (io_select_bits == 5'h16);
	assign io_sinks_22_bits_data = io_source_bits_data;
	assign io_sinks_22_bits_resp = io_source_bits_resp;
	assign io_sinks_22_bits_last = io_source_bits_last;
	assign io_sinks_23_valid = valid & (io_select_bits == 5'h17);
	assign io_sinks_23_bits_data = io_source_bits_data;
	assign io_sinks_23_bits_resp = io_source_bits_resp;
	assign io_sinks_23_bits_last = io_source_bits_last;
	assign io_sinks_24_valid = valid & (io_select_bits == 5'h18);
	assign io_sinks_24_bits_data = io_source_bits_data;
	assign io_sinks_24_bits_resp = io_source_bits_resp;
	assign io_sinks_24_bits_last = io_source_bits_last;
	assign io_sinks_25_valid = valid & (io_select_bits == 5'h19);
	assign io_sinks_25_bits_data = io_source_bits_data;
	assign io_sinks_25_bits_resp = io_source_bits_resp;
	assign io_sinks_25_bits_last = io_source_bits_last;
	assign io_sinks_26_valid = valid & (io_select_bits == 5'h1a);
	assign io_sinks_26_bits_data = io_source_bits_data;
	assign io_sinks_26_bits_resp = io_source_bits_resp;
	assign io_sinks_26_bits_last = io_source_bits_last;
	assign io_sinks_27_valid = valid & (io_select_bits == 5'h1b);
	assign io_sinks_27_bits_data = io_source_bits_data;
	assign io_sinks_27_bits_resp = io_source_bits_resp;
	assign io_sinks_27_bits_last = io_source_bits_last;
	assign io_sinks_28_valid = valid & (io_select_bits == 5'h1c);
	assign io_sinks_28_bits_data = io_source_bits_data;
	assign io_sinks_28_bits_resp = io_source_bits_resp;
	assign io_sinks_28_bits_last = io_source_bits_last;
	assign io_sinks_29_valid = valid & (io_select_bits == 5'h1d);
	assign io_sinks_29_bits_data = io_source_bits_data;
	assign io_sinks_29_bits_resp = io_source_bits_resp;
	assign io_sinks_29_bits_last = io_source_bits_last;
	assign io_sinks_30_valid = valid & (io_select_bits == 5'h1e);
	assign io_sinks_30_bits_data = io_source_bits_data;
	assign io_sinks_30_bits_resp = io_source_bits_resp;
	assign io_sinks_30_bits_last = io_source_bits_last;
	assign io_sinks_31_valid = valid & (&io_select_bits);
	assign io_sinks_31_bits_data = io_source_bits_data;
	assign io_sinks_31_bits_resp = io_source_bits_resp;
	assign io_sinks_31_bits_last = io_source_bits_last;
	assign io_select_ready = fire;
endmodule
module ram_32x5 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [4:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [4:0] R0_data;
	input [4:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [4:0] W0_data;
	reg [4:0] Memory [0:31];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 5'bxxxxx);
endmodule
module Queue32_UInt5 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [4:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [4:0] io_deq_bits;
	wire io_enq_ready_0;
	wire [4:0] _ram_ext_R0_data;
	reg [4:0] enq_ptr_value;
	reg [4:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire io_deq_valid_0 = io_enq_valid | ~empty;
	wire do_deq = (~empty & io_deq_ready) & io_deq_valid_0;
	wire do_enq = (~(empty & io_deq_ready) & io_enq_ready_0) & io_enq_valid;
	assign io_enq_ready_0 = io_deq_ready | ~(ptr_match & maybe_full);
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 5'h00;
			deq_ptr_value <= 5'h00;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 5'h01;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 5'h01;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_32x5 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = io_enq_ready_0;
	assign io_deq_valid = io_deq_valid_0;
	assign io_deq_bits = (empty ? io_enq_bits : _ram_ext_R0_data);
endmodule
module elasticMux_5 (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_data,
	io_sources_0_bits_strb,
	io_sources_0_bits_last,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_data,
	io_sources_1_bits_strb,
	io_sources_1_bits_last,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_data,
	io_sources_2_bits_strb,
	io_sources_2_bits_last,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_data,
	io_sources_3_bits_strb,
	io_sources_3_bits_last,
	io_sources_4_ready,
	io_sources_4_valid,
	io_sources_4_bits_data,
	io_sources_4_bits_strb,
	io_sources_4_bits_last,
	io_sources_5_ready,
	io_sources_5_valid,
	io_sources_5_bits_data,
	io_sources_5_bits_strb,
	io_sources_5_bits_last,
	io_sources_6_ready,
	io_sources_6_valid,
	io_sources_6_bits_data,
	io_sources_6_bits_strb,
	io_sources_6_bits_last,
	io_sources_7_ready,
	io_sources_7_valid,
	io_sources_7_bits_data,
	io_sources_7_bits_strb,
	io_sources_7_bits_last,
	io_sources_8_ready,
	io_sources_8_valid,
	io_sources_8_bits_data,
	io_sources_8_bits_strb,
	io_sources_8_bits_last,
	io_sources_9_ready,
	io_sources_9_valid,
	io_sources_9_bits_data,
	io_sources_9_bits_strb,
	io_sources_9_bits_last,
	io_sources_10_ready,
	io_sources_10_valid,
	io_sources_10_bits_data,
	io_sources_10_bits_strb,
	io_sources_10_bits_last,
	io_sources_11_ready,
	io_sources_11_valid,
	io_sources_11_bits_data,
	io_sources_11_bits_strb,
	io_sources_11_bits_last,
	io_sources_12_ready,
	io_sources_12_valid,
	io_sources_12_bits_data,
	io_sources_12_bits_strb,
	io_sources_12_bits_last,
	io_sources_13_ready,
	io_sources_13_valid,
	io_sources_13_bits_data,
	io_sources_13_bits_strb,
	io_sources_13_bits_last,
	io_sources_14_ready,
	io_sources_14_valid,
	io_sources_14_bits_data,
	io_sources_14_bits_strb,
	io_sources_14_bits_last,
	io_sources_15_ready,
	io_sources_15_valid,
	io_sources_15_bits_data,
	io_sources_15_bits_strb,
	io_sources_15_bits_last,
	io_sources_16_ready,
	io_sources_16_valid,
	io_sources_16_bits_data,
	io_sources_16_bits_strb,
	io_sources_16_bits_last,
	io_sources_17_ready,
	io_sources_17_valid,
	io_sources_17_bits_data,
	io_sources_17_bits_strb,
	io_sources_17_bits_last,
	io_sources_18_ready,
	io_sources_18_valid,
	io_sources_18_bits_data,
	io_sources_18_bits_strb,
	io_sources_18_bits_last,
	io_sources_19_ready,
	io_sources_19_valid,
	io_sources_19_bits_data,
	io_sources_19_bits_strb,
	io_sources_19_bits_last,
	io_sources_20_ready,
	io_sources_20_valid,
	io_sources_20_bits_data,
	io_sources_20_bits_strb,
	io_sources_20_bits_last,
	io_sources_21_ready,
	io_sources_21_valid,
	io_sources_21_bits_data,
	io_sources_21_bits_strb,
	io_sources_21_bits_last,
	io_sources_22_ready,
	io_sources_22_valid,
	io_sources_22_bits_data,
	io_sources_22_bits_strb,
	io_sources_22_bits_last,
	io_sources_23_ready,
	io_sources_23_valid,
	io_sources_23_bits_data,
	io_sources_23_bits_strb,
	io_sources_23_bits_last,
	io_sources_24_ready,
	io_sources_24_valid,
	io_sources_24_bits_data,
	io_sources_24_bits_strb,
	io_sources_24_bits_last,
	io_sources_25_ready,
	io_sources_25_valid,
	io_sources_25_bits_data,
	io_sources_25_bits_strb,
	io_sources_25_bits_last,
	io_sources_26_ready,
	io_sources_26_valid,
	io_sources_26_bits_data,
	io_sources_26_bits_strb,
	io_sources_26_bits_last,
	io_sources_27_ready,
	io_sources_27_valid,
	io_sources_27_bits_data,
	io_sources_27_bits_strb,
	io_sources_27_bits_last,
	io_sources_28_ready,
	io_sources_28_valid,
	io_sources_28_bits_data,
	io_sources_28_bits_strb,
	io_sources_28_bits_last,
	io_sources_29_ready,
	io_sources_29_valid,
	io_sources_29_bits_data,
	io_sources_29_bits_strb,
	io_sources_29_bits_last,
	io_sources_30_ready,
	io_sources_30_valid,
	io_sources_30_bits_data,
	io_sources_30_bits_strb,
	io_sources_30_bits_last,
	io_sources_31_ready,
	io_sources_31_valid,
	io_sources_31_bits_data,
	io_sources_31_bits_strb,
	io_sources_31_bits_last,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_data,
	io_sink_bits_strb,
	io_sink_bits_last,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [31:0] io_sources_0_bits_data;
	input [3:0] io_sources_0_bits_strb;
	input io_sources_0_bits_last;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [31:0] io_sources_1_bits_data;
	input [3:0] io_sources_1_bits_strb;
	input io_sources_1_bits_last;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [31:0] io_sources_2_bits_data;
	input [3:0] io_sources_2_bits_strb;
	input io_sources_2_bits_last;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [31:0] io_sources_3_bits_data;
	input [3:0] io_sources_3_bits_strb;
	input io_sources_3_bits_last;
	output wire io_sources_4_ready;
	input io_sources_4_valid;
	input [31:0] io_sources_4_bits_data;
	input [3:0] io_sources_4_bits_strb;
	input io_sources_4_bits_last;
	output wire io_sources_5_ready;
	input io_sources_5_valid;
	input [31:0] io_sources_5_bits_data;
	input [3:0] io_sources_5_bits_strb;
	input io_sources_5_bits_last;
	output wire io_sources_6_ready;
	input io_sources_6_valid;
	input [31:0] io_sources_6_bits_data;
	input [3:0] io_sources_6_bits_strb;
	input io_sources_6_bits_last;
	output wire io_sources_7_ready;
	input io_sources_7_valid;
	input [31:0] io_sources_7_bits_data;
	input [3:0] io_sources_7_bits_strb;
	input io_sources_7_bits_last;
	output wire io_sources_8_ready;
	input io_sources_8_valid;
	input [31:0] io_sources_8_bits_data;
	input [3:0] io_sources_8_bits_strb;
	input io_sources_8_bits_last;
	output wire io_sources_9_ready;
	input io_sources_9_valid;
	input [31:0] io_sources_9_bits_data;
	input [3:0] io_sources_9_bits_strb;
	input io_sources_9_bits_last;
	output wire io_sources_10_ready;
	input io_sources_10_valid;
	input [31:0] io_sources_10_bits_data;
	input [3:0] io_sources_10_bits_strb;
	input io_sources_10_bits_last;
	output wire io_sources_11_ready;
	input io_sources_11_valid;
	input [31:0] io_sources_11_bits_data;
	input [3:0] io_sources_11_bits_strb;
	input io_sources_11_bits_last;
	output wire io_sources_12_ready;
	input io_sources_12_valid;
	input [31:0] io_sources_12_bits_data;
	input [3:0] io_sources_12_bits_strb;
	input io_sources_12_bits_last;
	output wire io_sources_13_ready;
	input io_sources_13_valid;
	input [31:0] io_sources_13_bits_data;
	input [3:0] io_sources_13_bits_strb;
	input io_sources_13_bits_last;
	output wire io_sources_14_ready;
	input io_sources_14_valid;
	input [31:0] io_sources_14_bits_data;
	input [3:0] io_sources_14_bits_strb;
	input io_sources_14_bits_last;
	output wire io_sources_15_ready;
	input io_sources_15_valid;
	input [31:0] io_sources_15_bits_data;
	input [3:0] io_sources_15_bits_strb;
	input io_sources_15_bits_last;
	output wire io_sources_16_ready;
	input io_sources_16_valid;
	input [31:0] io_sources_16_bits_data;
	input [3:0] io_sources_16_bits_strb;
	input io_sources_16_bits_last;
	output wire io_sources_17_ready;
	input io_sources_17_valid;
	input [31:0] io_sources_17_bits_data;
	input [3:0] io_sources_17_bits_strb;
	input io_sources_17_bits_last;
	output wire io_sources_18_ready;
	input io_sources_18_valid;
	input [31:0] io_sources_18_bits_data;
	input [3:0] io_sources_18_bits_strb;
	input io_sources_18_bits_last;
	output wire io_sources_19_ready;
	input io_sources_19_valid;
	input [31:0] io_sources_19_bits_data;
	input [3:0] io_sources_19_bits_strb;
	input io_sources_19_bits_last;
	output wire io_sources_20_ready;
	input io_sources_20_valid;
	input [31:0] io_sources_20_bits_data;
	input [3:0] io_sources_20_bits_strb;
	input io_sources_20_bits_last;
	output wire io_sources_21_ready;
	input io_sources_21_valid;
	input [31:0] io_sources_21_bits_data;
	input [3:0] io_sources_21_bits_strb;
	input io_sources_21_bits_last;
	output wire io_sources_22_ready;
	input io_sources_22_valid;
	input [31:0] io_sources_22_bits_data;
	input [3:0] io_sources_22_bits_strb;
	input io_sources_22_bits_last;
	output wire io_sources_23_ready;
	input io_sources_23_valid;
	input [31:0] io_sources_23_bits_data;
	input [3:0] io_sources_23_bits_strb;
	input io_sources_23_bits_last;
	output wire io_sources_24_ready;
	input io_sources_24_valid;
	input [31:0] io_sources_24_bits_data;
	input [3:0] io_sources_24_bits_strb;
	input io_sources_24_bits_last;
	output wire io_sources_25_ready;
	input io_sources_25_valid;
	input [31:0] io_sources_25_bits_data;
	input [3:0] io_sources_25_bits_strb;
	input io_sources_25_bits_last;
	output wire io_sources_26_ready;
	input io_sources_26_valid;
	input [31:0] io_sources_26_bits_data;
	input [3:0] io_sources_26_bits_strb;
	input io_sources_26_bits_last;
	output wire io_sources_27_ready;
	input io_sources_27_valid;
	input [31:0] io_sources_27_bits_data;
	input [3:0] io_sources_27_bits_strb;
	input io_sources_27_bits_last;
	output wire io_sources_28_ready;
	input io_sources_28_valid;
	input [31:0] io_sources_28_bits_data;
	input [3:0] io_sources_28_bits_strb;
	input io_sources_28_bits_last;
	output wire io_sources_29_ready;
	input io_sources_29_valid;
	input [31:0] io_sources_29_bits_data;
	input [3:0] io_sources_29_bits_strb;
	input io_sources_29_bits_last;
	output wire io_sources_30_ready;
	input io_sources_30_valid;
	input [31:0] io_sources_30_bits_data;
	input [3:0] io_sources_30_bits_strb;
	input io_sources_30_bits_last;
	output wire io_sources_31_ready;
	input io_sources_31_valid;
	input [31:0] io_sources_31_bits_data;
	input [3:0] io_sources_31_bits_strb;
	input io_sources_31_bits_last;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [31:0] io_sink_bits_data;
	output wire [3:0] io_sink_bits_strb;
	output wire io_sink_bits_last;
	output wire io_select_ready;
	input io_select_valid;
	input [4:0] io_select_bits;
	wire [31:0] _GEN = {io_sources_31_valid, io_sources_30_valid, io_sources_29_valid, io_sources_28_valid, io_sources_27_valid, io_sources_26_valid, io_sources_25_valid, io_sources_24_valid, io_sources_23_valid, io_sources_22_valid, io_sources_21_valid, io_sources_20_valid, io_sources_19_valid, io_sources_18_valid, io_sources_17_valid, io_sources_16_valid, io_sources_15_valid, io_sources_14_valid, io_sources_13_valid, io_sources_12_valid, io_sources_11_valid, io_sources_10_valid, io_sources_9_valid, io_sources_8_valid, io_sources_7_valid, io_sources_6_valid, io_sources_5_valid, io_sources_4_valid, io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [1023:0] _GEN_0 = {io_sources_31_bits_data, io_sources_30_bits_data, io_sources_29_bits_data, io_sources_28_bits_data, io_sources_27_bits_data, io_sources_26_bits_data, io_sources_25_bits_data, io_sources_24_bits_data, io_sources_23_bits_data, io_sources_22_bits_data, io_sources_21_bits_data, io_sources_20_bits_data, io_sources_19_bits_data, io_sources_18_bits_data, io_sources_17_bits_data, io_sources_16_bits_data, io_sources_15_bits_data, io_sources_14_bits_data, io_sources_13_bits_data, io_sources_12_bits_data, io_sources_11_bits_data, io_sources_10_bits_data, io_sources_9_bits_data, io_sources_8_bits_data, io_sources_7_bits_data, io_sources_6_bits_data, io_sources_5_bits_data, io_sources_4_bits_data, io_sources_3_bits_data, io_sources_2_bits_data, io_sources_1_bits_data, io_sources_0_bits_data};
	wire [127:0] _GEN_1 = {io_sources_31_bits_strb, io_sources_30_bits_strb, io_sources_29_bits_strb, io_sources_28_bits_strb, io_sources_27_bits_strb, io_sources_26_bits_strb, io_sources_25_bits_strb, io_sources_24_bits_strb, io_sources_23_bits_strb, io_sources_22_bits_strb, io_sources_21_bits_strb, io_sources_20_bits_strb, io_sources_19_bits_strb, io_sources_18_bits_strb, io_sources_17_bits_strb, io_sources_16_bits_strb, io_sources_15_bits_strb, io_sources_14_bits_strb, io_sources_13_bits_strb, io_sources_12_bits_strb, io_sources_11_bits_strb, io_sources_10_bits_strb, io_sources_9_bits_strb, io_sources_8_bits_strb, io_sources_7_bits_strb, io_sources_6_bits_strb, io_sources_5_bits_strb, io_sources_4_bits_strb, io_sources_3_bits_strb, io_sources_2_bits_strb, io_sources_1_bits_strb, io_sources_0_bits_strb};
	wire [31:0] _GEN_2 = {io_sources_31_bits_last, io_sources_30_bits_last, io_sources_29_bits_last, io_sources_28_bits_last, io_sources_27_bits_last, io_sources_26_bits_last, io_sources_25_bits_last, io_sources_24_bits_last, io_sources_23_bits_last, io_sources_22_bits_last, io_sources_21_bits_last, io_sources_20_bits_last, io_sources_19_bits_last, io_sources_18_bits_last, io_sources_17_bits_last, io_sources_16_bits_last, io_sources_15_bits_last, io_sources_14_bits_last, io_sources_13_bits_last, io_sources_12_bits_last, io_sources_11_bits_last, io_sources_10_bits_last, io_sources_9_bits_last, io_sources_8_bits_last, io_sources_7_bits_last, io_sources_6_bits_last, io_sources_5_bits_last, io_sources_4_bits_last, io_sources_3_bits_last, io_sources_2_bits_last, io_sources_1_bits_last, io_sources_0_bits_last};
	wire valid = io_select_valid & _GEN[io_select_bits];
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & (io_select_bits == 5'h00);
	assign io_sources_1_ready = fire & (io_select_bits == 5'h01);
	assign io_sources_2_ready = fire & (io_select_bits == 5'h02);
	assign io_sources_3_ready = fire & (io_select_bits == 5'h03);
	assign io_sources_4_ready = fire & (io_select_bits == 5'h04);
	assign io_sources_5_ready = fire & (io_select_bits == 5'h05);
	assign io_sources_6_ready = fire & (io_select_bits == 5'h06);
	assign io_sources_7_ready = fire & (io_select_bits == 5'h07);
	assign io_sources_8_ready = fire & (io_select_bits == 5'h08);
	assign io_sources_9_ready = fire & (io_select_bits == 5'h09);
	assign io_sources_10_ready = fire & (io_select_bits == 5'h0a);
	assign io_sources_11_ready = fire & (io_select_bits == 5'h0b);
	assign io_sources_12_ready = fire & (io_select_bits == 5'h0c);
	assign io_sources_13_ready = fire & (io_select_bits == 5'h0d);
	assign io_sources_14_ready = fire & (io_select_bits == 5'h0e);
	assign io_sources_15_ready = fire & (io_select_bits == 5'h0f);
	assign io_sources_16_ready = fire & (io_select_bits == 5'h10);
	assign io_sources_17_ready = fire & (io_select_bits == 5'h11);
	assign io_sources_18_ready = fire & (io_select_bits == 5'h12);
	assign io_sources_19_ready = fire & (io_select_bits == 5'h13);
	assign io_sources_20_ready = fire & (io_select_bits == 5'h14);
	assign io_sources_21_ready = fire & (io_select_bits == 5'h15);
	assign io_sources_22_ready = fire & (io_select_bits == 5'h16);
	assign io_sources_23_ready = fire & (io_select_bits == 5'h17);
	assign io_sources_24_ready = fire & (io_select_bits == 5'h18);
	assign io_sources_25_ready = fire & (io_select_bits == 5'h19);
	assign io_sources_26_ready = fire & (io_select_bits == 5'h1a);
	assign io_sources_27_ready = fire & (io_select_bits == 5'h1b);
	assign io_sources_28_ready = fire & (io_select_bits == 5'h1c);
	assign io_sources_29_ready = fire & (io_select_bits == 5'h1d);
	assign io_sources_30_ready = fire & (io_select_bits == 5'h1e);
	assign io_sources_31_ready = fire & (&io_select_bits);
	assign io_sink_valid = valid;
	assign io_sink_bits_data = _GEN_0[io_select_bits * 32+:32];
	assign io_sink_bits_strb = _GEN_1[io_select_bits * 4+:4];
	assign io_sink_bits_last = _GEN_2[io_select_bits];
	assign io_select_ready = fire & _GEN_2[io_select_bits];
endmodule
module elasticDemux_10 (
	io_source_ready,
	io_source_valid,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_4_ready,
	io_sinks_4_valid,
	io_sinks_5_ready,
	io_sinks_5_valid,
	io_sinks_6_ready,
	io_sinks_6_valid,
	io_sinks_7_ready,
	io_sinks_7_valid,
	io_sinks_8_ready,
	io_sinks_8_valid,
	io_sinks_9_ready,
	io_sinks_9_valid,
	io_sinks_10_ready,
	io_sinks_10_valid,
	io_sinks_11_ready,
	io_sinks_11_valid,
	io_sinks_12_ready,
	io_sinks_12_valid,
	io_sinks_13_ready,
	io_sinks_13_valid,
	io_sinks_14_ready,
	io_sinks_14_valid,
	io_sinks_15_ready,
	io_sinks_15_valid,
	io_sinks_16_ready,
	io_sinks_16_valid,
	io_sinks_17_ready,
	io_sinks_17_valid,
	io_sinks_18_ready,
	io_sinks_18_valid,
	io_sinks_19_ready,
	io_sinks_19_valid,
	io_sinks_20_ready,
	io_sinks_20_valid,
	io_sinks_21_ready,
	io_sinks_21_valid,
	io_sinks_22_ready,
	io_sinks_22_valid,
	io_sinks_23_ready,
	io_sinks_23_valid,
	io_sinks_24_ready,
	io_sinks_24_valid,
	io_sinks_25_ready,
	io_sinks_25_valid,
	io_sinks_26_ready,
	io_sinks_26_valid,
	io_sinks_27_ready,
	io_sinks_27_valid,
	io_sinks_28_ready,
	io_sinks_28_valid,
	io_sinks_29_ready,
	io_sinks_29_valid,
	io_sinks_30_ready,
	io_sinks_30_valid,
	io_sinks_31_ready,
	io_sinks_31_valid,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	input io_sinks_4_ready;
	output wire io_sinks_4_valid;
	input io_sinks_5_ready;
	output wire io_sinks_5_valid;
	input io_sinks_6_ready;
	output wire io_sinks_6_valid;
	input io_sinks_7_ready;
	output wire io_sinks_7_valid;
	input io_sinks_8_ready;
	output wire io_sinks_8_valid;
	input io_sinks_9_ready;
	output wire io_sinks_9_valid;
	input io_sinks_10_ready;
	output wire io_sinks_10_valid;
	input io_sinks_11_ready;
	output wire io_sinks_11_valid;
	input io_sinks_12_ready;
	output wire io_sinks_12_valid;
	input io_sinks_13_ready;
	output wire io_sinks_13_valid;
	input io_sinks_14_ready;
	output wire io_sinks_14_valid;
	input io_sinks_15_ready;
	output wire io_sinks_15_valid;
	input io_sinks_16_ready;
	output wire io_sinks_16_valid;
	input io_sinks_17_ready;
	output wire io_sinks_17_valid;
	input io_sinks_18_ready;
	output wire io_sinks_18_valid;
	input io_sinks_19_ready;
	output wire io_sinks_19_valid;
	input io_sinks_20_ready;
	output wire io_sinks_20_valid;
	input io_sinks_21_ready;
	output wire io_sinks_21_valid;
	input io_sinks_22_ready;
	output wire io_sinks_22_valid;
	input io_sinks_23_ready;
	output wire io_sinks_23_valid;
	input io_sinks_24_ready;
	output wire io_sinks_24_valid;
	input io_sinks_25_ready;
	output wire io_sinks_25_valid;
	input io_sinks_26_ready;
	output wire io_sinks_26_valid;
	input io_sinks_27_ready;
	output wire io_sinks_27_valid;
	input io_sinks_28_ready;
	output wire io_sinks_28_valid;
	input io_sinks_29_ready;
	output wire io_sinks_29_valid;
	input io_sinks_30_ready;
	output wire io_sinks_30_valid;
	input io_sinks_31_ready;
	output wire io_sinks_31_valid;
	output wire io_select_ready;
	input io_select_valid;
	input [4:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [31:0] _GEN = {io_sinks_31_ready, io_sinks_30_ready, io_sinks_29_ready, io_sinks_28_ready, io_sinks_27_ready, io_sinks_26_ready, io_sinks_25_ready, io_sinks_24_ready, io_sinks_23_ready, io_sinks_22_ready, io_sinks_21_ready, io_sinks_20_ready, io_sinks_19_ready, io_sinks_18_ready, io_sinks_17_ready, io_sinks_16_ready, io_sinks_15_ready, io_sinks_14_ready, io_sinks_13_ready, io_sinks_12_ready, io_sinks_11_ready, io_sinks_10_ready, io_sinks_9_ready, io_sinks_8_ready, io_sinks_7_ready, io_sinks_6_ready, io_sinks_5_ready, io_sinks_4_ready, io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 5'h00);
	assign io_sinks_1_valid = valid & (io_select_bits == 5'h01);
	assign io_sinks_2_valid = valid & (io_select_bits == 5'h02);
	assign io_sinks_3_valid = valid & (io_select_bits == 5'h03);
	assign io_sinks_4_valid = valid & (io_select_bits == 5'h04);
	assign io_sinks_5_valid = valid & (io_select_bits == 5'h05);
	assign io_sinks_6_valid = valid & (io_select_bits == 5'h06);
	assign io_sinks_7_valid = valid & (io_select_bits == 5'h07);
	assign io_sinks_8_valid = valid & (io_select_bits == 5'h08);
	assign io_sinks_9_valid = valid & (io_select_bits == 5'h09);
	assign io_sinks_10_valid = valid & (io_select_bits == 5'h0a);
	assign io_sinks_11_valid = valid & (io_select_bits == 5'h0b);
	assign io_sinks_12_valid = valid & (io_select_bits == 5'h0c);
	assign io_sinks_13_valid = valid & (io_select_bits == 5'h0d);
	assign io_sinks_14_valid = valid & (io_select_bits == 5'h0e);
	assign io_sinks_15_valid = valid & (io_select_bits == 5'h0f);
	assign io_sinks_16_valid = valid & (io_select_bits == 5'h10);
	assign io_sinks_17_valid = valid & (io_select_bits == 5'h11);
	assign io_sinks_18_valid = valid & (io_select_bits == 5'h12);
	assign io_sinks_19_valid = valid & (io_select_bits == 5'h13);
	assign io_sinks_20_valid = valid & (io_select_bits == 5'h14);
	assign io_sinks_21_valid = valid & (io_select_bits == 5'h15);
	assign io_sinks_22_valid = valid & (io_select_bits == 5'h16);
	assign io_sinks_23_valid = valid & (io_select_bits == 5'h17);
	assign io_sinks_24_valid = valid & (io_select_bits == 5'h18);
	assign io_sinks_25_valid = valid & (io_select_bits == 5'h19);
	assign io_sinks_26_valid = valid & (io_select_bits == 5'h1a);
	assign io_sinks_27_valid = valid & (io_select_bits == 5'h1b);
	assign io_sinks_28_valid = valid & (io_select_bits == 5'h1c);
	assign io_sinks_29_valid = valid & (io_select_bits == 5'h1d);
	assign io_sinks_30_valid = valid & (io_select_bits == 5'h1e);
	assign io_sinks_31_valid = valid & (&io_select_bits);
	assign io_select_ready = fire;
endmodule
module axi4FullMux_3 (
	clock,
	reset,
	s_axi_0_ar_ready,
	s_axi_0_ar_valid,
	s_axi_0_ar_bits_addr,
	s_axi_0_r_ready,
	s_axi_0_r_valid,
	s_axi_0_r_bits_data,
	s_axi_0_aw_ready,
	s_axi_0_aw_valid,
	s_axi_0_aw_bits_addr,
	s_axi_0_w_ready,
	s_axi_0_w_valid,
	s_axi_0_w_bits_data,
	s_axi_0_b_valid,
	s_axi_1_ar_ready,
	s_axi_1_ar_valid,
	s_axi_1_ar_bits_addr,
	s_axi_1_r_ready,
	s_axi_1_r_valid,
	s_axi_1_r_bits_data,
	s_axi_1_aw_ready,
	s_axi_1_aw_valid,
	s_axi_1_aw_bits_addr,
	s_axi_1_w_ready,
	s_axi_1_w_valid,
	s_axi_1_w_bits_data,
	s_axi_1_b_valid,
	s_axi_2_ar_ready,
	s_axi_2_ar_valid,
	s_axi_2_ar_bits_addr,
	s_axi_2_r_ready,
	s_axi_2_r_valid,
	s_axi_2_r_bits_data,
	s_axi_2_aw_ready,
	s_axi_2_aw_valid,
	s_axi_2_aw_bits_addr,
	s_axi_2_w_ready,
	s_axi_2_w_valid,
	s_axi_2_w_bits_data,
	s_axi_2_b_valid,
	s_axi_3_ar_ready,
	s_axi_3_ar_valid,
	s_axi_3_ar_bits_addr,
	s_axi_3_r_ready,
	s_axi_3_r_valid,
	s_axi_3_r_bits_data,
	s_axi_3_aw_ready,
	s_axi_3_aw_valid,
	s_axi_3_aw_bits_addr,
	s_axi_3_w_ready,
	s_axi_3_w_valid,
	s_axi_3_w_bits_data,
	s_axi_3_b_valid,
	s_axi_4_ar_ready,
	s_axi_4_ar_valid,
	s_axi_4_ar_bits_addr,
	s_axi_4_r_ready,
	s_axi_4_r_valid,
	s_axi_4_r_bits_data,
	s_axi_4_aw_ready,
	s_axi_4_aw_valid,
	s_axi_4_aw_bits_addr,
	s_axi_4_w_ready,
	s_axi_4_w_valid,
	s_axi_4_w_bits_data,
	s_axi_4_b_valid,
	s_axi_5_ar_ready,
	s_axi_5_ar_valid,
	s_axi_5_ar_bits_addr,
	s_axi_5_r_ready,
	s_axi_5_r_valid,
	s_axi_5_r_bits_data,
	s_axi_5_aw_ready,
	s_axi_5_aw_valid,
	s_axi_5_aw_bits_addr,
	s_axi_5_w_ready,
	s_axi_5_w_valid,
	s_axi_5_w_bits_data,
	s_axi_5_b_valid,
	s_axi_6_ar_ready,
	s_axi_6_ar_valid,
	s_axi_6_ar_bits_addr,
	s_axi_6_r_ready,
	s_axi_6_r_valid,
	s_axi_6_r_bits_data,
	s_axi_6_aw_ready,
	s_axi_6_aw_valid,
	s_axi_6_aw_bits_addr,
	s_axi_6_w_ready,
	s_axi_6_w_valid,
	s_axi_6_w_bits_data,
	s_axi_6_b_valid,
	s_axi_7_ar_ready,
	s_axi_7_ar_valid,
	s_axi_7_ar_bits_addr,
	s_axi_7_r_ready,
	s_axi_7_r_valid,
	s_axi_7_r_bits_data,
	s_axi_7_aw_ready,
	s_axi_7_aw_valid,
	s_axi_7_aw_bits_addr,
	s_axi_7_w_ready,
	s_axi_7_w_valid,
	s_axi_7_w_bits_data,
	s_axi_7_b_valid,
	s_axi_8_ar_ready,
	s_axi_8_ar_valid,
	s_axi_8_ar_bits_addr,
	s_axi_8_r_ready,
	s_axi_8_r_valid,
	s_axi_8_r_bits_data,
	s_axi_8_aw_ready,
	s_axi_8_aw_valid,
	s_axi_8_aw_bits_addr,
	s_axi_8_w_ready,
	s_axi_8_w_valid,
	s_axi_8_w_bits_data,
	s_axi_8_b_valid,
	s_axi_9_ar_ready,
	s_axi_9_ar_valid,
	s_axi_9_ar_bits_addr,
	s_axi_9_r_ready,
	s_axi_9_r_valid,
	s_axi_9_r_bits_data,
	s_axi_9_aw_ready,
	s_axi_9_aw_valid,
	s_axi_9_aw_bits_addr,
	s_axi_9_w_ready,
	s_axi_9_w_valid,
	s_axi_9_w_bits_data,
	s_axi_9_b_valid,
	s_axi_10_ar_ready,
	s_axi_10_ar_valid,
	s_axi_10_ar_bits_addr,
	s_axi_10_r_ready,
	s_axi_10_r_valid,
	s_axi_10_r_bits_data,
	s_axi_10_aw_ready,
	s_axi_10_aw_valid,
	s_axi_10_aw_bits_addr,
	s_axi_10_w_ready,
	s_axi_10_w_valid,
	s_axi_10_w_bits_data,
	s_axi_10_b_valid,
	s_axi_11_ar_ready,
	s_axi_11_ar_valid,
	s_axi_11_ar_bits_addr,
	s_axi_11_r_ready,
	s_axi_11_r_valid,
	s_axi_11_r_bits_data,
	s_axi_11_aw_ready,
	s_axi_11_aw_valid,
	s_axi_11_aw_bits_addr,
	s_axi_11_w_ready,
	s_axi_11_w_valid,
	s_axi_11_w_bits_data,
	s_axi_11_b_valid,
	s_axi_12_ar_ready,
	s_axi_12_ar_valid,
	s_axi_12_ar_bits_addr,
	s_axi_12_r_ready,
	s_axi_12_r_valid,
	s_axi_12_r_bits_data,
	s_axi_12_aw_ready,
	s_axi_12_aw_valid,
	s_axi_12_aw_bits_addr,
	s_axi_12_w_ready,
	s_axi_12_w_valid,
	s_axi_12_w_bits_data,
	s_axi_12_b_valid,
	s_axi_13_ar_ready,
	s_axi_13_ar_valid,
	s_axi_13_ar_bits_addr,
	s_axi_13_r_ready,
	s_axi_13_r_valid,
	s_axi_13_r_bits_data,
	s_axi_13_aw_ready,
	s_axi_13_aw_valid,
	s_axi_13_aw_bits_addr,
	s_axi_13_w_ready,
	s_axi_13_w_valid,
	s_axi_13_w_bits_data,
	s_axi_13_b_valid,
	s_axi_14_ar_ready,
	s_axi_14_ar_valid,
	s_axi_14_ar_bits_addr,
	s_axi_14_r_ready,
	s_axi_14_r_valid,
	s_axi_14_r_bits_data,
	s_axi_14_aw_ready,
	s_axi_14_aw_valid,
	s_axi_14_aw_bits_addr,
	s_axi_14_w_ready,
	s_axi_14_w_valid,
	s_axi_14_w_bits_data,
	s_axi_14_b_valid,
	s_axi_15_ar_ready,
	s_axi_15_ar_valid,
	s_axi_15_ar_bits_addr,
	s_axi_15_r_ready,
	s_axi_15_r_valid,
	s_axi_15_r_bits_data,
	s_axi_15_aw_ready,
	s_axi_15_aw_valid,
	s_axi_15_aw_bits_addr,
	s_axi_15_w_ready,
	s_axi_15_w_valid,
	s_axi_15_w_bits_data,
	s_axi_15_b_valid,
	s_axi_16_ar_ready,
	s_axi_16_ar_valid,
	s_axi_16_ar_bits_addr,
	s_axi_16_r_ready,
	s_axi_16_r_valid,
	s_axi_16_r_bits_data,
	s_axi_17_ar_ready,
	s_axi_17_ar_valid,
	s_axi_17_ar_bits_addr,
	s_axi_17_r_ready,
	s_axi_17_r_valid,
	s_axi_17_r_bits_data,
	s_axi_18_ar_ready,
	s_axi_18_ar_valid,
	s_axi_18_ar_bits_addr,
	s_axi_18_r_ready,
	s_axi_18_r_valid,
	s_axi_18_r_bits_data,
	s_axi_19_ar_ready,
	s_axi_19_ar_valid,
	s_axi_19_ar_bits_addr,
	s_axi_19_r_ready,
	s_axi_19_r_valid,
	s_axi_19_r_bits_data,
	s_axi_20_ar_ready,
	s_axi_20_ar_valid,
	s_axi_20_ar_bits_addr,
	s_axi_20_r_ready,
	s_axi_20_r_valid,
	s_axi_20_r_bits_data,
	s_axi_21_ar_ready,
	s_axi_21_ar_valid,
	s_axi_21_ar_bits_addr,
	s_axi_21_r_ready,
	s_axi_21_r_valid,
	s_axi_21_r_bits_data,
	s_axi_22_ar_ready,
	s_axi_22_ar_valid,
	s_axi_22_ar_bits_addr,
	s_axi_22_r_ready,
	s_axi_22_r_valid,
	s_axi_22_r_bits_data,
	s_axi_23_ar_ready,
	s_axi_23_ar_valid,
	s_axi_23_ar_bits_addr,
	s_axi_23_r_ready,
	s_axi_23_r_valid,
	s_axi_23_r_bits_data,
	s_axi_24_ar_ready,
	s_axi_24_ar_valid,
	s_axi_24_ar_bits_addr,
	s_axi_24_r_ready,
	s_axi_24_r_valid,
	s_axi_24_r_bits_data,
	s_axi_25_ar_ready,
	s_axi_25_ar_valid,
	s_axi_25_ar_bits_addr,
	s_axi_25_r_ready,
	s_axi_25_r_valid,
	s_axi_25_r_bits_data,
	s_axi_26_ar_ready,
	s_axi_26_ar_valid,
	s_axi_26_ar_bits_addr,
	s_axi_26_r_ready,
	s_axi_26_r_valid,
	s_axi_26_r_bits_data,
	s_axi_27_ar_ready,
	s_axi_27_ar_valid,
	s_axi_27_ar_bits_addr,
	s_axi_27_r_ready,
	s_axi_27_r_valid,
	s_axi_27_r_bits_data,
	s_axi_28_ar_ready,
	s_axi_28_ar_valid,
	s_axi_28_ar_bits_addr,
	s_axi_28_r_ready,
	s_axi_28_r_valid,
	s_axi_28_r_bits_data,
	s_axi_29_ar_ready,
	s_axi_29_ar_valid,
	s_axi_29_ar_bits_addr,
	s_axi_29_r_ready,
	s_axi_29_r_valid,
	s_axi_29_r_bits_data,
	s_axi_30_ar_ready,
	s_axi_30_ar_valid,
	s_axi_30_ar_bits_addr,
	s_axi_30_r_ready,
	s_axi_30_r_valid,
	s_axi_30_r_bits_data,
	s_axi_31_ar_ready,
	s_axi_31_ar_valid,
	s_axi_31_ar_bits_addr,
	s_axi_31_r_ready,
	s_axi_31_r_valid,
	s_axi_31_r_bits_data,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_id,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_id,
	m_axi_r_bits_data,
	m_axi_r_bits_resp,
	m_axi_r_bits_last,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_id,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_strb,
	m_axi_w_bits_last,
	m_axi_b_ready,
	m_axi_b_valid,
	m_axi_b_bits_id,
	m_axi_b_bits_resp
);
	input clock;
	input reset;
	output wire s_axi_0_ar_ready;
	input s_axi_0_ar_valid;
	input [63:0] s_axi_0_ar_bits_addr;
	input s_axi_0_r_ready;
	output wire s_axi_0_r_valid;
	output wire [31:0] s_axi_0_r_bits_data;
	output wire s_axi_0_aw_ready;
	input s_axi_0_aw_valid;
	input [63:0] s_axi_0_aw_bits_addr;
	output wire s_axi_0_w_ready;
	input s_axi_0_w_valid;
	input [31:0] s_axi_0_w_bits_data;
	output wire s_axi_0_b_valid;
	output wire s_axi_1_ar_ready;
	input s_axi_1_ar_valid;
	input [63:0] s_axi_1_ar_bits_addr;
	input s_axi_1_r_ready;
	output wire s_axi_1_r_valid;
	output wire [31:0] s_axi_1_r_bits_data;
	output wire s_axi_1_aw_ready;
	input s_axi_1_aw_valid;
	input [63:0] s_axi_1_aw_bits_addr;
	output wire s_axi_1_w_ready;
	input s_axi_1_w_valid;
	input [31:0] s_axi_1_w_bits_data;
	output wire s_axi_1_b_valid;
	output wire s_axi_2_ar_ready;
	input s_axi_2_ar_valid;
	input [63:0] s_axi_2_ar_bits_addr;
	input s_axi_2_r_ready;
	output wire s_axi_2_r_valid;
	output wire [31:0] s_axi_2_r_bits_data;
	output wire s_axi_2_aw_ready;
	input s_axi_2_aw_valid;
	input [63:0] s_axi_2_aw_bits_addr;
	output wire s_axi_2_w_ready;
	input s_axi_2_w_valid;
	input [31:0] s_axi_2_w_bits_data;
	output wire s_axi_2_b_valid;
	output wire s_axi_3_ar_ready;
	input s_axi_3_ar_valid;
	input [63:0] s_axi_3_ar_bits_addr;
	input s_axi_3_r_ready;
	output wire s_axi_3_r_valid;
	output wire [31:0] s_axi_3_r_bits_data;
	output wire s_axi_3_aw_ready;
	input s_axi_3_aw_valid;
	input [63:0] s_axi_3_aw_bits_addr;
	output wire s_axi_3_w_ready;
	input s_axi_3_w_valid;
	input [31:0] s_axi_3_w_bits_data;
	output wire s_axi_3_b_valid;
	output wire s_axi_4_ar_ready;
	input s_axi_4_ar_valid;
	input [63:0] s_axi_4_ar_bits_addr;
	input s_axi_4_r_ready;
	output wire s_axi_4_r_valid;
	output wire [31:0] s_axi_4_r_bits_data;
	output wire s_axi_4_aw_ready;
	input s_axi_4_aw_valid;
	input [63:0] s_axi_4_aw_bits_addr;
	output wire s_axi_4_w_ready;
	input s_axi_4_w_valid;
	input [31:0] s_axi_4_w_bits_data;
	output wire s_axi_4_b_valid;
	output wire s_axi_5_ar_ready;
	input s_axi_5_ar_valid;
	input [63:0] s_axi_5_ar_bits_addr;
	input s_axi_5_r_ready;
	output wire s_axi_5_r_valid;
	output wire [31:0] s_axi_5_r_bits_data;
	output wire s_axi_5_aw_ready;
	input s_axi_5_aw_valid;
	input [63:0] s_axi_5_aw_bits_addr;
	output wire s_axi_5_w_ready;
	input s_axi_5_w_valid;
	input [31:0] s_axi_5_w_bits_data;
	output wire s_axi_5_b_valid;
	output wire s_axi_6_ar_ready;
	input s_axi_6_ar_valid;
	input [63:0] s_axi_6_ar_bits_addr;
	input s_axi_6_r_ready;
	output wire s_axi_6_r_valid;
	output wire [31:0] s_axi_6_r_bits_data;
	output wire s_axi_6_aw_ready;
	input s_axi_6_aw_valid;
	input [63:0] s_axi_6_aw_bits_addr;
	output wire s_axi_6_w_ready;
	input s_axi_6_w_valid;
	input [31:0] s_axi_6_w_bits_data;
	output wire s_axi_6_b_valid;
	output wire s_axi_7_ar_ready;
	input s_axi_7_ar_valid;
	input [63:0] s_axi_7_ar_bits_addr;
	input s_axi_7_r_ready;
	output wire s_axi_7_r_valid;
	output wire [31:0] s_axi_7_r_bits_data;
	output wire s_axi_7_aw_ready;
	input s_axi_7_aw_valid;
	input [63:0] s_axi_7_aw_bits_addr;
	output wire s_axi_7_w_ready;
	input s_axi_7_w_valid;
	input [31:0] s_axi_7_w_bits_data;
	output wire s_axi_7_b_valid;
	output wire s_axi_8_ar_ready;
	input s_axi_8_ar_valid;
	input [63:0] s_axi_8_ar_bits_addr;
	input s_axi_8_r_ready;
	output wire s_axi_8_r_valid;
	output wire [31:0] s_axi_8_r_bits_data;
	output wire s_axi_8_aw_ready;
	input s_axi_8_aw_valid;
	input [63:0] s_axi_8_aw_bits_addr;
	output wire s_axi_8_w_ready;
	input s_axi_8_w_valid;
	input [31:0] s_axi_8_w_bits_data;
	output wire s_axi_8_b_valid;
	output wire s_axi_9_ar_ready;
	input s_axi_9_ar_valid;
	input [63:0] s_axi_9_ar_bits_addr;
	input s_axi_9_r_ready;
	output wire s_axi_9_r_valid;
	output wire [31:0] s_axi_9_r_bits_data;
	output wire s_axi_9_aw_ready;
	input s_axi_9_aw_valid;
	input [63:0] s_axi_9_aw_bits_addr;
	output wire s_axi_9_w_ready;
	input s_axi_9_w_valid;
	input [31:0] s_axi_9_w_bits_data;
	output wire s_axi_9_b_valid;
	output wire s_axi_10_ar_ready;
	input s_axi_10_ar_valid;
	input [63:0] s_axi_10_ar_bits_addr;
	input s_axi_10_r_ready;
	output wire s_axi_10_r_valid;
	output wire [31:0] s_axi_10_r_bits_data;
	output wire s_axi_10_aw_ready;
	input s_axi_10_aw_valid;
	input [63:0] s_axi_10_aw_bits_addr;
	output wire s_axi_10_w_ready;
	input s_axi_10_w_valid;
	input [31:0] s_axi_10_w_bits_data;
	output wire s_axi_10_b_valid;
	output wire s_axi_11_ar_ready;
	input s_axi_11_ar_valid;
	input [63:0] s_axi_11_ar_bits_addr;
	input s_axi_11_r_ready;
	output wire s_axi_11_r_valid;
	output wire [31:0] s_axi_11_r_bits_data;
	output wire s_axi_11_aw_ready;
	input s_axi_11_aw_valid;
	input [63:0] s_axi_11_aw_bits_addr;
	output wire s_axi_11_w_ready;
	input s_axi_11_w_valid;
	input [31:0] s_axi_11_w_bits_data;
	output wire s_axi_11_b_valid;
	output wire s_axi_12_ar_ready;
	input s_axi_12_ar_valid;
	input [63:0] s_axi_12_ar_bits_addr;
	input s_axi_12_r_ready;
	output wire s_axi_12_r_valid;
	output wire [31:0] s_axi_12_r_bits_data;
	output wire s_axi_12_aw_ready;
	input s_axi_12_aw_valid;
	input [63:0] s_axi_12_aw_bits_addr;
	output wire s_axi_12_w_ready;
	input s_axi_12_w_valid;
	input [31:0] s_axi_12_w_bits_data;
	output wire s_axi_12_b_valid;
	output wire s_axi_13_ar_ready;
	input s_axi_13_ar_valid;
	input [63:0] s_axi_13_ar_bits_addr;
	input s_axi_13_r_ready;
	output wire s_axi_13_r_valid;
	output wire [31:0] s_axi_13_r_bits_data;
	output wire s_axi_13_aw_ready;
	input s_axi_13_aw_valid;
	input [63:0] s_axi_13_aw_bits_addr;
	output wire s_axi_13_w_ready;
	input s_axi_13_w_valid;
	input [31:0] s_axi_13_w_bits_data;
	output wire s_axi_13_b_valid;
	output wire s_axi_14_ar_ready;
	input s_axi_14_ar_valid;
	input [63:0] s_axi_14_ar_bits_addr;
	input s_axi_14_r_ready;
	output wire s_axi_14_r_valid;
	output wire [31:0] s_axi_14_r_bits_data;
	output wire s_axi_14_aw_ready;
	input s_axi_14_aw_valid;
	input [63:0] s_axi_14_aw_bits_addr;
	output wire s_axi_14_w_ready;
	input s_axi_14_w_valid;
	input [31:0] s_axi_14_w_bits_data;
	output wire s_axi_14_b_valid;
	output wire s_axi_15_ar_ready;
	input s_axi_15_ar_valid;
	input [63:0] s_axi_15_ar_bits_addr;
	input s_axi_15_r_ready;
	output wire s_axi_15_r_valid;
	output wire [31:0] s_axi_15_r_bits_data;
	output wire s_axi_15_aw_ready;
	input s_axi_15_aw_valid;
	input [63:0] s_axi_15_aw_bits_addr;
	output wire s_axi_15_w_ready;
	input s_axi_15_w_valid;
	input [31:0] s_axi_15_w_bits_data;
	output wire s_axi_15_b_valid;
	output wire s_axi_16_ar_ready;
	input s_axi_16_ar_valid;
	input [63:0] s_axi_16_ar_bits_addr;
	input s_axi_16_r_ready;
	output wire s_axi_16_r_valid;
	output wire [31:0] s_axi_16_r_bits_data;
	output wire s_axi_17_ar_ready;
	input s_axi_17_ar_valid;
	input [63:0] s_axi_17_ar_bits_addr;
	input s_axi_17_r_ready;
	output wire s_axi_17_r_valid;
	output wire [31:0] s_axi_17_r_bits_data;
	output wire s_axi_18_ar_ready;
	input s_axi_18_ar_valid;
	input [63:0] s_axi_18_ar_bits_addr;
	input s_axi_18_r_ready;
	output wire s_axi_18_r_valid;
	output wire [31:0] s_axi_18_r_bits_data;
	output wire s_axi_19_ar_ready;
	input s_axi_19_ar_valid;
	input [63:0] s_axi_19_ar_bits_addr;
	input s_axi_19_r_ready;
	output wire s_axi_19_r_valid;
	output wire [31:0] s_axi_19_r_bits_data;
	output wire s_axi_20_ar_ready;
	input s_axi_20_ar_valid;
	input [63:0] s_axi_20_ar_bits_addr;
	input s_axi_20_r_ready;
	output wire s_axi_20_r_valid;
	output wire [31:0] s_axi_20_r_bits_data;
	output wire s_axi_21_ar_ready;
	input s_axi_21_ar_valid;
	input [63:0] s_axi_21_ar_bits_addr;
	input s_axi_21_r_ready;
	output wire s_axi_21_r_valid;
	output wire [31:0] s_axi_21_r_bits_data;
	output wire s_axi_22_ar_ready;
	input s_axi_22_ar_valid;
	input [63:0] s_axi_22_ar_bits_addr;
	input s_axi_22_r_ready;
	output wire s_axi_22_r_valid;
	output wire [31:0] s_axi_22_r_bits_data;
	output wire s_axi_23_ar_ready;
	input s_axi_23_ar_valid;
	input [63:0] s_axi_23_ar_bits_addr;
	input s_axi_23_r_ready;
	output wire s_axi_23_r_valid;
	output wire [31:0] s_axi_23_r_bits_data;
	output wire s_axi_24_ar_ready;
	input s_axi_24_ar_valid;
	input [63:0] s_axi_24_ar_bits_addr;
	input s_axi_24_r_ready;
	output wire s_axi_24_r_valid;
	output wire [31:0] s_axi_24_r_bits_data;
	output wire s_axi_25_ar_ready;
	input s_axi_25_ar_valid;
	input [63:0] s_axi_25_ar_bits_addr;
	input s_axi_25_r_ready;
	output wire s_axi_25_r_valid;
	output wire [31:0] s_axi_25_r_bits_data;
	output wire s_axi_26_ar_ready;
	input s_axi_26_ar_valid;
	input [63:0] s_axi_26_ar_bits_addr;
	input s_axi_26_r_ready;
	output wire s_axi_26_r_valid;
	output wire [31:0] s_axi_26_r_bits_data;
	output wire s_axi_27_ar_ready;
	input s_axi_27_ar_valid;
	input [63:0] s_axi_27_ar_bits_addr;
	input s_axi_27_r_ready;
	output wire s_axi_27_r_valid;
	output wire [31:0] s_axi_27_r_bits_data;
	output wire s_axi_28_ar_ready;
	input s_axi_28_ar_valid;
	input [63:0] s_axi_28_ar_bits_addr;
	input s_axi_28_r_ready;
	output wire s_axi_28_r_valid;
	output wire [31:0] s_axi_28_r_bits_data;
	output wire s_axi_29_ar_ready;
	input s_axi_29_ar_valid;
	input [63:0] s_axi_29_ar_bits_addr;
	input s_axi_29_r_ready;
	output wire s_axi_29_r_valid;
	output wire [31:0] s_axi_29_r_bits_data;
	output wire s_axi_30_ar_ready;
	input s_axi_30_ar_valid;
	input [63:0] s_axi_30_ar_bits_addr;
	input s_axi_30_r_ready;
	output wire s_axi_30_r_valid;
	output wire [31:0] s_axi_30_r_bits_data;
	output wire s_axi_31_ar_ready;
	input s_axi_31_ar_valid;
	input [63:0] s_axi_31_ar_bits_addr;
	input s_axi_31_r_ready;
	output wire s_axi_31_r_valid;
	output wire [31:0] s_axi_31_r_bits_data;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [4:0] m_axi_ar_bits_id;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [4:0] m_axi_r_bits_id;
	input [31:0] m_axi_r_bits_data;
	input [1:0] m_axi_r_bits_resp;
	input m_axi_r_bits_last;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [4:0] m_axi_aw_bits_id;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [31:0] m_axi_w_bits_data;
	output wire [3:0] m_axi_w_bits_strb;
	output wire m_axi_w_bits_last;
	output wire m_axi_b_ready;
	input m_axi_b_valid;
	input [4:0] m_axi_b_bits_id;
	input [1:0] m_axi_b_bits_resp;
	wire _write_demux_io_source_ready;
	wire _write_demux_io_sinks_0_valid;
	wire _write_demux_io_sinks_1_valid;
	wire _write_demux_io_sinks_2_valid;
	wire _write_demux_io_sinks_3_valid;
	wire _write_demux_io_sinks_4_valid;
	wire _write_demux_io_sinks_5_valid;
	wire _write_demux_io_sinks_6_valid;
	wire _write_demux_io_sinks_7_valid;
	wire _write_demux_io_sinks_8_valid;
	wire _write_demux_io_sinks_9_valid;
	wire _write_demux_io_sinks_10_valid;
	wire _write_demux_io_sinks_11_valid;
	wire _write_demux_io_sinks_12_valid;
	wire _write_demux_io_sinks_13_valid;
	wire _write_demux_io_sinks_14_valid;
	wire _write_demux_io_sinks_15_valid;
	wire _write_demux_io_sinks_16_valid;
	wire _write_demux_io_sinks_17_valid;
	wire _write_demux_io_sinks_18_valid;
	wire _write_demux_io_sinks_19_valid;
	wire _write_demux_io_sinks_20_valid;
	wire _write_demux_io_sinks_21_valid;
	wire _write_demux_io_sinks_22_valid;
	wire _write_demux_io_sinks_23_valid;
	wire _write_demux_io_sinks_24_valid;
	wire _write_demux_io_sinks_25_valid;
	wire _write_demux_io_sinks_26_valid;
	wire _write_demux_io_sinks_27_valid;
	wire _write_demux_io_sinks_28_valid;
	wire _write_demux_io_sinks_29_valid;
	wire _write_demux_io_sinks_30_valid;
	wire _write_demux_io_sinks_31_valid;
	wire _write_demux_io_select_ready;
	wire _write_mux_io_sources_0_ready;
	wire _write_mux_io_sources_1_ready;
	wire _write_mux_io_sources_2_ready;
	wire _write_mux_io_sources_3_ready;
	wire _write_mux_io_sources_4_ready;
	wire _write_mux_io_sources_5_ready;
	wire _write_mux_io_sources_6_ready;
	wire _write_mux_io_sources_7_ready;
	wire _write_mux_io_sources_8_ready;
	wire _write_mux_io_sources_9_ready;
	wire _write_mux_io_sources_10_ready;
	wire _write_mux_io_sources_11_ready;
	wire _write_mux_io_sources_12_ready;
	wire _write_mux_io_sources_13_ready;
	wire _write_mux_io_sources_14_ready;
	wire _write_mux_io_sources_15_ready;
	wire _write_mux_io_sources_16_ready;
	wire _write_mux_io_sources_17_ready;
	wire _write_mux_io_sources_18_ready;
	wire _write_mux_io_sources_19_ready;
	wire _write_mux_io_sources_20_ready;
	wire _write_mux_io_sources_21_ready;
	wire _write_mux_io_sources_22_ready;
	wire _write_mux_io_sources_23_ready;
	wire _write_mux_io_sources_24_ready;
	wire _write_mux_io_sources_25_ready;
	wire _write_mux_io_sources_26_ready;
	wire _write_mux_io_sources_27_ready;
	wire _write_mux_io_sources_28_ready;
	wire _write_mux_io_sources_29_ready;
	wire _write_mux_io_sources_30_ready;
	wire _write_mux_io_sources_31_ready;
	wire _write_mux_io_sink_valid;
	wire [31:0] _write_mux_io_sink_bits_data;
	wire [3:0] _write_mux_io_sink_bits_strb;
	wire _write_mux_io_sink_bits_last;
	wire _write_mux_io_select_ready;
	wire _write_arbiter_io_sources_0_ready;
	wire _write_arbiter_io_sources_1_ready;
	wire _write_arbiter_io_sources_2_ready;
	wire _write_arbiter_io_sources_3_ready;
	wire _write_arbiter_io_sources_4_ready;
	wire _write_arbiter_io_sources_5_ready;
	wire _write_arbiter_io_sources_6_ready;
	wire _write_arbiter_io_sources_7_ready;
	wire _write_arbiter_io_sources_8_ready;
	wire _write_arbiter_io_sources_9_ready;
	wire _write_arbiter_io_sources_10_ready;
	wire _write_arbiter_io_sources_11_ready;
	wire _write_arbiter_io_sources_12_ready;
	wire _write_arbiter_io_sources_13_ready;
	wire _write_arbiter_io_sources_14_ready;
	wire _write_arbiter_io_sources_15_ready;
	wire _write_arbiter_io_sources_16_ready;
	wire _write_arbiter_io_sources_17_ready;
	wire _write_arbiter_io_sources_18_ready;
	wire _write_arbiter_io_sources_19_ready;
	wire _write_arbiter_io_sources_20_ready;
	wire _write_arbiter_io_sources_21_ready;
	wire _write_arbiter_io_sources_22_ready;
	wire _write_arbiter_io_sources_23_ready;
	wire _write_arbiter_io_sources_24_ready;
	wire _write_arbiter_io_sources_25_ready;
	wire _write_arbiter_io_sources_26_ready;
	wire _write_arbiter_io_sources_27_ready;
	wire _write_arbiter_io_sources_28_ready;
	wire _write_arbiter_io_sources_29_ready;
	wire _write_arbiter_io_sources_30_ready;
	wire _write_arbiter_io_sources_31_ready;
	wire _write_arbiter_io_sink_valid;
	wire [4:0] _write_arbiter_io_sink_bits_id;
	wire [63:0] _write_arbiter_io_sink_bits_addr;
	wire [7:0] _write_arbiter_io_sink_bits_len;
	wire [2:0] _write_arbiter_io_sink_bits_size;
	wire [1:0] _write_arbiter_io_sink_bits_burst;
	wire _write_arbiter_io_sink_bits_lock;
	wire [3:0] _write_arbiter_io_sink_bits_cache;
	wire [2:0] _write_arbiter_io_sink_bits_prot;
	wire [3:0] _write_arbiter_io_sink_bits_qos;
	wire [3:0] _write_arbiter_io_sink_bits_region;
	wire _write_arbiter_io_select_valid;
	wire [4:0] _write_arbiter_io_select_bits;
	wire _write_portQueue_io_enq_ready;
	wire _write_portQueue_io_deq_valid;
	wire [4:0] _write_portQueue_io_deq_bits;
	wire _read_demux_io_source_ready;
	wire _read_demux_io_sinks_0_valid;
	wire [31:0] _read_demux_io_sinks_0_bits_data;
	wire [1:0] _read_demux_io_sinks_0_bits_resp;
	wire _read_demux_io_sinks_0_bits_last;
	wire _read_demux_io_sinks_1_valid;
	wire [31:0] _read_demux_io_sinks_1_bits_data;
	wire [1:0] _read_demux_io_sinks_1_bits_resp;
	wire _read_demux_io_sinks_1_bits_last;
	wire _read_demux_io_sinks_2_valid;
	wire [31:0] _read_demux_io_sinks_2_bits_data;
	wire [1:0] _read_demux_io_sinks_2_bits_resp;
	wire _read_demux_io_sinks_2_bits_last;
	wire _read_demux_io_sinks_3_valid;
	wire [31:0] _read_demux_io_sinks_3_bits_data;
	wire [1:0] _read_demux_io_sinks_3_bits_resp;
	wire _read_demux_io_sinks_3_bits_last;
	wire _read_demux_io_sinks_4_valid;
	wire [31:0] _read_demux_io_sinks_4_bits_data;
	wire [1:0] _read_demux_io_sinks_4_bits_resp;
	wire _read_demux_io_sinks_4_bits_last;
	wire _read_demux_io_sinks_5_valid;
	wire [31:0] _read_demux_io_sinks_5_bits_data;
	wire [1:0] _read_demux_io_sinks_5_bits_resp;
	wire _read_demux_io_sinks_5_bits_last;
	wire _read_demux_io_sinks_6_valid;
	wire [31:0] _read_demux_io_sinks_6_bits_data;
	wire [1:0] _read_demux_io_sinks_6_bits_resp;
	wire _read_demux_io_sinks_6_bits_last;
	wire _read_demux_io_sinks_7_valid;
	wire [31:0] _read_demux_io_sinks_7_bits_data;
	wire [1:0] _read_demux_io_sinks_7_bits_resp;
	wire _read_demux_io_sinks_7_bits_last;
	wire _read_demux_io_sinks_8_valid;
	wire [31:0] _read_demux_io_sinks_8_bits_data;
	wire [1:0] _read_demux_io_sinks_8_bits_resp;
	wire _read_demux_io_sinks_8_bits_last;
	wire _read_demux_io_sinks_9_valid;
	wire [31:0] _read_demux_io_sinks_9_bits_data;
	wire [1:0] _read_demux_io_sinks_9_bits_resp;
	wire _read_demux_io_sinks_9_bits_last;
	wire _read_demux_io_sinks_10_valid;
	wire [31:0] _read_demux_io_sinks_10_bits_data;
	wire [1:0] _read_demux_io_sinks_10_bits_resp;
	wire _read_demux_io_sinks_10_bits_last;
	wire _read_demux_io_sinks_11_valid;
	wire [31:0] _read_demux_io_sinks_11_bits_data;
	wire [1:0] _read_demux_io_sinks_11_bits_resp;
	wire _read_demux_io_sinks_11_bits_last;
	wire _read_demux_io_sinks_12_valid;
	wire [31:0] _read_demux_io_sinks_12_bits_data;
	wire [1:0] _read_demux_io_sinks_12_bits_resp;
	wire _read_demux_io_sinks_12_bits_last;
	wire _read_demux_io_sinks_13_valid;
	wire [31:0] _read_demux_io_sinks_13_bits_data;
	wire [1:0] _read_demux_io_sinks_13_bits_resp;
	wire _read_demux_io_sinks_13_bits_last;
	wire _read_demux_io_sinks_14_valid;
	wire [31:0] _read_demux_io_sinks_14_bits_data;
	wire [1:0] _read_demux_io_sinks_14_bits_resp;
	wire _read_demux_io_sinks_14_bits_last;
	wire _read_demux_io_sinks_15_valid;
	wire [31:0] _read_demux_io_sinks_15_bits_data;
	wire [1:0] _read_demux_io_sinks_15_bits_resp;
	wire _read_demux_io_sinks_15_bits_last;
	wire _read_demux_io_sinks_16_valid;
	wire [31:0] _read_demux_io_sinks_16_bits_data;
	wire [1:0] _read_demux_io_sinks_16_bits_resp;
	wire _read_demux_io_sinks_16_bits_last;
	wire _read_demux_io_sinks_17_valid;
	wire [31:0] _read_demux_io_sinks_17_bits_data;
	wire [1:0] _read_demux_io_sinks_17_bits_resp;
	wire _read_demux_io_sinks_17_bits_last;
	wire _read_demux_io_sinks_18_valid;
	wire [31:0] _read_demux_io_sinks_18_bits_data;
	wire [1:0] _read_demux_io_sinks_18_bits_resp;
	wire _read_demux_io_sinks_18_bits_last;
	wire _read_demux_io_sinks_19_valid;
	wire [31:0] _read_demux_io_sinks_19_bits_data;
	wire [1:0] _read_demux_io_sinks_19_bits_resp;
	wire _read_demux_io_sinks_19_bits_last;
	wire _read_demux_io_sinks_20_valid;
	wire [31:0] _read_demux_io_sinks_20_bits_data;
	wire [1:0] _read_demux_io_sinks_20_bits_resp;
	wire _read_demux_io_sinks_20_bits_last;
	wire _read_demux_io_sinks_21_valid;
	wire [31:0] _read_demux_io_sinks_21_bits_data;
	wire [1:0] _read_demux_io_sinks_21_bits_resp;
	wire _read_demux_io_sinks_21_bits_last;
	wire _read_demux_io_sinks_22_valid;
	wire [31:0] _read_demux_io_sinks_22_bits_data;
	wire [1:0] _read_demux_io_sinks_22_bits_resp;
	wire _read_demux_io_sinks_22_bits_last;
	wire _read_demux_io_sinks_23_valid;
	wire [31:0] _read_demux_io_sinks_23_bits_data;
	wire [1:0] _read_demux_io_sinks_23_bits_resp;
	wire _read_demux_io_sinks_23_bits_last;
	wire _read_demux_io_sinks_24_valid;
	wire [31:0] _read_demux_io_sinks_24_bits_data;
	wire [1:0] _read_demux_io_sinks_24_bits_resp;
	wire _read_demux_io_sinks_24_bits_last;
	wire _read_demux_io_sinks_25_valid;
	wire [31:0] _read_demux_io_sinks_25_bits_data;
	wire [1:0] _read_demux_io_sinks_25_bits_resp;
	wire _read_demux_io_sinks_25_bits_last;
	wire _read_demux_io_sinks_26_valid;
	wire [31:0] _read_demux_io_sinks_26_bits_data;
	wire [1:0] _read_demux_io_sinks_26_bits_resp;
	wire _read_demux_io_sinks_26_bits_last;
	wire _read_demux_io_sinks_27_valid;
	wire [31:0] _read_demux_io_sinks_27_bits_data;
	wire [1:0] _read_demux_io_sinks_27_bits_resp;
	wire _read_demux_io_sinks_27_bits_last;
	wire _read_demux_io_sinks_28_valid;
	wire [31:0] _read_demux_io_sinks_28_bits_data;
	wire [1:0] _read_demux_io_sinks_28_bits_resp;
	wire _read_demux_io_sinks_28_bits_last;
	wire _read_demux_io_sinks_29_valid;
	wire [31:0] _read_demux_io_sinks_29_bits_data;
	wire [1:0] _read_demux_io_sinks_29_bits_resp;
	wire _read_demux_io_sinks_29_bits_last;
	wire _read_demux_io_sinks_30_valid;
	wire [31:0] _read_demux_io_sinks_30_bits_data;
	wire [1:0] _read_demux_io_sinks_30_bits_resp;
	wire _read_demux_io_sinks_30_bits_last;
	wire _read_demux_io_sinks_31_valid;
	wire [31:0] _read_demux_io_sinks_31_bits_data;
	wire [1:0] _read_demux_io_sinks_31_bits_resp;
	wire _read_demux_io_sinks_31_bits_last;
	wire _read_demux_io_select_ready;
	wire _read_arbiter_io_sources_0_ready;
	wire _read_arbiter_io_sources_1_ready;
	wire _read_arbiter_io_sources_2_ready;
	wire _read_arbiter_io_sources_3_ready;
	wire _read_arbiter_io_sources_4_ready;
	wire _read_arbiter_io_sources_5_ready;
	wire _read_arbiter_io_sources_6_ready;
	wire _read_arbiter_io_sources_7_ready;
	wire _read_arbiter_io_sources_8_ready;
	wire _read_arbiter_io_sources_9_ready;
	wire _read_arbiter_io_sources_10_ready;
	wire _read_arbiter_io_sources_11_ready;
	wire _read_arbiter_io_sources_12_ready;
	wire _read_arbiter_io_sources_13_ready;
	wire _read_arbiter_io_sources_14_ready;
	wire _read_arbiter_io_sources_15_ready;
	wire _read_arbiter_io_sources_16_ready;
	wire _read_arbiter_io_sources_17_ready;
	wire _read_arbiter_io_sources_18_ready;
	wire _read_arbiter_io_sources_19_ready;
	wire _read_arbiter_io_sources_20_ready;
	wire _read_arbiter_io_sources_21_ready;
	wire _read_arbiter_io_sources_22_ready;
	wire _read_arbiter_io_sources_23_ready;
	wire _read_arbiter_io_sources_24_ready;
	wire _read_arbiter_io_sources_25_ready;
	wire _read_arbiter_io_sources_26_ready;
	wire _read_arbiter_io_sources_27_ready;
	wire _read_arbiter_io_sources_28_ready;
	wire _read_arbiter_io_sources_29_ready;
	wire _read_arbiter_io_sources_30_ready;
	wire _read_arbiter_io_sources_31_ready;
	wire _read_arbiter_io_sink_valid;
	wire [4:0] _read_arbiter_io_sink_bits_id;
	wire [63:0] _read_arbiter_io_sink_bits_addr;
	wire [7:0] _read_arbiter_io_sink_bits_len;
	wire [2:0] _read_arbiter_io_sink_bits_size;
	wire [1:0] _read_arbiter_io_sink_bits_burst;
	wire _read_arbiter_io_sink_bits_lock;
	wire [3:0] _read_arbiter_io_sink_bits_cache;
	wire [2:0] _read_arbiter_io_sink_bits_prot;
	wire [3:0] _read_arbiter_io_sink_bits_qos;
	wire [3:0] _read_arbiter_io_sink_bits_region;
	wire _m_axi__sinkBuffer_1_io_deq_valid;
	wire [4:0] _m_axi__sinkBuffer_1_io_deq_bits_id;
	wire _m_axi__sourceBuffer_2_io_enq_ready;
	wire _m_axi__sourceBuffer_1_io_enq_ready;
	wire _m_axi__sinkBuffer_io_deq_valid;
	wire [4:0] _m_axi__sinkBuffer_io_deq_bits_id;
	wire [31:0] _m_axi__sinkBuffer_io_deq_bits_data;
	wire [1:0] _m_axi__sinkBuffer_io_deq_bits_resp;
	wire _m_axi__sinkBuffer_io_deq_bits_last;
	wire _m_axi__sourceBuffer_io_enq_ready;
	wire _s_axi__buffered_sinkBuffer_63_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_95_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_95_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_95_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_95_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_94_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_94_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_94_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_62_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_93_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_93_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_93_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_61_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_92_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_92_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_92_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_92_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_91_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_91_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_91_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_60_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_90_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_90_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_90_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_59_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_89_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_89_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_89_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_89_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_88_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_88_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_88_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_58_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_87_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_87_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_87_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_57_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_86_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_86_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_86_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_86_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_85_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_85_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_85_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_56_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_84_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_84_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_84_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_55_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_83_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_83_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_83_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_83_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_82_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_82_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_82_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_54_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_81_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_81_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_81_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_53_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_80_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_80_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_80_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_80_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_79_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_79_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_79_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_52_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_78_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_78_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_78_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_51_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_77_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_77_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_77_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_77_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_76_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_76_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_76_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_50_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_75_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_75_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_75_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_49_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_74_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_74_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_74_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_74_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_73_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_73_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_73_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_48_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_72_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_72_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_72_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_47_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_71_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_71_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_71_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_71_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_70_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_70_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_70_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_46_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_69_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_69_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_69_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_45_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_68_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_68_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_68_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_68_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_67_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_67_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_67_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_44_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_66_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_66_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_66_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_43_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_65_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_65_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_65_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_65_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_64_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_64_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_64_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_42_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_63_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_63_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_63_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_41_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_62_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_62_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_62_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_62_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_61_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_61_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_61_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_40_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_60_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_60_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_60_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_39_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_59_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_59_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_59_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_59_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_58_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_58_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_58_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_38_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_57_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_57_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_57_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_37_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_56_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_56_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_56_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_56_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_55_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_55_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_55_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_36_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_54_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_54_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_54_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_35_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_53_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_53_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_53_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_53_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_52_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_52_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_52_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_34_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_51_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_51_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_51_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_33_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_50_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_50_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_50_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_50_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_49_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_49_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_49_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_32_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_48_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_48_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_48_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_31_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_47_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_47_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_47_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_47_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_46_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_46_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_46_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_30_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_45_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_45_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_45_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_29_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_44_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_44_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_44_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_44_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_43_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_43_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_43_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_28_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_42_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_42_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_42_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_27_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_41_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_41_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_41_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_41_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_40_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_40_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_40_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_26_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_39_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_39_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_39_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_25_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_38_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_38_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_38_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_38_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_37_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_37_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_37_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_24_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_36_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_36_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_36_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_23_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_35_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_35_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_35_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_35_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_34_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_34_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_34_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_22_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_33_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_33_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_33_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_21_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_32_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_32_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_32_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_32_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_31_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_31_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_31_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_20_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_30_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_30_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_30_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_19_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_29_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_29_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_29_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_29_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_28_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_28_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_28_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_18_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_27_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_27_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_27_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_17_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_26_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_26_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_26_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_26_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_25_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_25_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_25_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_16_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_24_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_24_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_24_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_15_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_23_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_23_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_23_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_23_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_22_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_22_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_22_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_14_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_21_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_21_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_21_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_13_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_20_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_20_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_20_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_20_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_19_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_19_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_19_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_12_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_18_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_18_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_18_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_11_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_17_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_17_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_17_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_17_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_16_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_16_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_16_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_10_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_15_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_15_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_15_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_9_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_14_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_14_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_14_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_14_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_13_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_13_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_13_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_8_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_12_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_12_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_12_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_7_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_11_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_11_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_11_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_11_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_10_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_10_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_10_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_6_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_9_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_9_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_9_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_5_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_8_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_8_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_8_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_8_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_7_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_7_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_7_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_4_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_6_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_6_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_6_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_3_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_5_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_5_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_4_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_4_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_2_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_3_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_3_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_1_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_valid;
	wire [31:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_data;
	wire [3:0] _s_axi__buffered_sourceBuffer_2_io_deq_bits_strb;
	wire _s_axi__buffered_sourceBuffer_2_io_deq_bits_last;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_1_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_1_io_deq_bits_region;
	wire _s_axi__buffered_sinkBuffer_io_enq_ready;
	wire _s_axi__buffered_sourceBuffer_io_deq_valid;
	wire [63:0] _s_axi__buffered_sourceBuffer_io_deq_bits_addr;
	wire [7:0] _s_axi__buffered_sourceBuffer_io_deq_bits_len;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_size;
	wire [1:0] _s_axi__buffered_sourceBuffer_io_deq_bits_burst;
	wire _s_axi__buffered_sourceBuffer_io_deq_bits_lock;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_cache;
	wire [2:0] _s_axi__buffered_sourceBuffer_io_deq_bits_prot;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_qos;
	wire [3:0] _s_axi__buffered_sourceBuffer_io_deq_bits_region;
	reg read_eagerFork_regs_0;
	reg read_eagerFork_regs_1;
	wire read_eagerFork_m_axi__r_ready_qual1_0 = _read_demux_io_source_ready | read_eagerFork_regs_0;
	wire read_eagerFork_m_axi__r_ready_qual1_1 = _read_demux_io_select_ready | read_eagerFork_regs_1;
	wire m_axi__r_ready = read_eagerFork_m_axi__r_ready_qual1_0 & read_eagerFork_m_axi__r_ready_qual1_1;
	reg write_eagerFork_regs_0;
	reg write_eagerFork_regs_1;
	wire write_eagerFork_m_axi__b_ready_qual1_0 = _write_demux_io_source_ready | write_eagerFork_regs_0;
	wire write_eagerFork_m_axi__b_ready_qual1_1 = _write_demux_io_select_ready | write_eagerFork_regs_1;
	wire m_axi__b_ready = write_eagerFork_m_axi__b_ready_qual1_0 & write_eagerFork_m_axi__b_ready_qual1_1;
	always @(posedge clock)
		if (reset) begin
			read_eagerFork_regs_0 <= 1'h0;
			read_eagerFork_regs_1 <= 1'h0;
			write_eagerFork_regs_0 <= 1'h0;
			write_eagerFork_regs_1 <= 1'h0;
		end
		else begin
			read_eagerFork_regs_0 <= (read_eagerFork_m_axi__r_ready_qual1_0 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			read_eagerFork_regs_1 <= (read_eagerFork_m_axi__r_ready_qual1_1 & _m_axi__sinkBuffer_io_deq_valid) & ~m_axi__r_ready;
			write_eagerFork_regs_0 <= (write_eagerFork_m_axi__b_ready_qual1_0 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
			write_eagerFork_regs_1 <= (write_eagerFork_m_axi__b_ready_qual1_1 & _m_axi__sinkBuffer_1_io_deq_valid) & ~m_axi__b_ready;
		end
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_ar_ready),
		.io_enq_valid(s_axi_0_ar_valid),
		.io_enq_bits_addr(s_axi_0_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_0_valid),
		.io_enq_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_deq_ready(s_axi_0_r_ready),
		.io_deq_valid(s_axi_0_r_valid),
		.io_deq_bits_data(s_axi_0_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_aw_ready),
		.io_enq_valid(s_axi_0_aw_valid),
		.io_enq_bits_addr(s_axi_0_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_0_w_ready),
		.io_enq_valid(s_axi_0_w_valid),
		.io_enq_bits_data(s_axi_0_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_0_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_0_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_0_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_ar_ready),
		.io_enq_valid(s_axi_1_ar_valid),
		.io_enq_bits_addr(s_axi_1_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_1_valid),
		.io_enq_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_deq_ready(s_axi_1_r_ready),
		.io_deq_valid(s_axi_1_r_valid),
		.io_deq_bits_data(s_axi_1_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_4(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_aw_ready),
		.io_enq_valid(s_axi_1_aw_valid),
		.io_enq_bits_addr(s_axi_1_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_1_w_ready),
		.io_enq_valid(s_axi_1_w_valid),
		.io_enq_bits_data(s_axi_1_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_1_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_1_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_1_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_6(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_2_ar_ready),
		.io_enq_valid(s_axi_2_ar_valid),
		.io_enq_bits_addr(s_axi_2_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_2_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_6_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_6_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_6_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_6_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_6_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_6_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_6_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_6_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_6_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_6_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_4(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_4_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_2_valid),
		.io_enq_bits_data(_read_demux_io_sinks_2_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_2_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_2_bits_last),
		.io_deq_ready(s_axi_2_r_ready),
		.io_deq_valid(s_axi_2_r_valid),
		.io_deq_bits_data(s_axi_2_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_7(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_2_aw_ready),
		.io_enq_valid(s_axi_2_aw_valid),
		.io_enq_bits_addr(s_axi_2_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_2_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_7_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_7_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_7_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_7_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_7_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_7_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_7_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_7_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_7_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_7_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_8(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_2_w_ready),
		.io_enq_valid(s_axi_2_w_valid),
		.io_enq_bits_data(s_axi_2_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_2_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_8_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_8_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_8_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_8_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_5_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_2_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_2_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_9(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_3_ar_ready),
		.io_enq_valid(s_axi_3_ar_valid),
		.io_enq_bits_addr(s_axi_3_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_3_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_9_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_9_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_9_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_9_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_9_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_9_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_9_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_9_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_9_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_9_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_6(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_6_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_3_valid),
		.io_enq_bits_data(_read_demux_io_sinks_3_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_3_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_3_bits_last),
		.io_deq_ready(s_axi_3_r_ready),
		.io_deq_valid(s_axi_3_r_valid),
		.io_deq_bits_data(s_axi_3_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_10(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_3_aw_ready),
		.io_enq_valid(s_axi_3_aw_valid),
		.io_enq_bits_addr(s_axi_3_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_3_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_10_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_10_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_10_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_10_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_10_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_10_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_10_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_10_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_10_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_10_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_11(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_3_w_ready),
		.io_enq_valid(s_axi_3_w_valid),
		.io_enq_bits_data(s_axi_3_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_3_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_11_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_11_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_11_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_11_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_7(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_7_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_3_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_3_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_12(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_4_ar_ready),
		.io_enq_valid(s_axi_4_ar_valid),
		.io_enq_bits_addr(s_axi_4_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_4_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_12_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_12_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_12_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_12_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_12_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_12_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_12_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_12_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_12_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_12_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_8(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_8_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_4_valid),
		.io_enq_bits_data(_read_demux_io_sinks_4_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_4_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_4_bits_last),
		.io_deq_ready(s_axi_4_r_ready),
		.io_deq_valid(s_axi_4_r_valid),
		.io_deq_bits_data(s_axi_4_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_13(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_4_aw_ready),
		.io_enq_valid(s_axi_4_aw_valid),
		.io_enq_bits_addr(s_axi_4_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_4_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_13_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_13_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_13_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_13_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_13_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_13_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_13_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_13_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_13_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_13_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_14(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_4_w_ready),
		.io_enq_valid(s_axi_4_w_valid),
		.io_enq_bits_data(s_axi_4_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_4_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_14_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_14_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_14_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_14_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_9(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_9_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_4_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_4_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_15(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_5_ar_ready),
		.io_enq_valid(s_axi_5_ar_valid),
		.io_enq_bits_addr(s_axi_5_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_5_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_15_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_15_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_15_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_15_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_15_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_15_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_15_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_15_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_15_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_15_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_10(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_10_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_5_valid),
		.io_enq_bits_data(_read_demux_io_sinks_5_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_5_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_5_bits_last),
		.io_deq_ready(s_axi_5_r_ready),
		.io_deq_valid(s_axi_5_r_valid),
		.io_deq_bits_data(s_axi_5_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_16(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_5_aw_ready),
		.io_enq_valid(s_axi_5_aw_valid),
		.io_enq_bits_addr(s_axi_5_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_5_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_16_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_16_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_16_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_16_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_16_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_16_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_16_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_16_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_16_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_16_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_17(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_5_w_ready),
		.io_enq_valid(s_axi_5_w_valid),
		.io_enq_bits_data(s_axi_5_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_5_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_17_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_17_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_17_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_17_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_11(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_11_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_5_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_5_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_18(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_6_ar_ready),
		.io_enq_valid(s_axi_6_ar_valid),
		.io_enq_bits_addr(s_axi_6_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_6_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_18_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_18_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_18_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_18_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_18_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_18_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_18_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_18_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_18_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_18_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_12(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_12_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_6_valid),
		.io_enq_bits_data(_read_demux_io_sinks_6_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_6_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_6_bits_last),
		.io_deq_ready(s_axi_6_r_ready),
		.io_deq_valid(s_axi_6_r_valid),
		.io_deq_bits_data(s_axi_6_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_19(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_6_aw_ready),
		.io_enq_valid(s_axi_6_aw_valid),
		.io_enq_bits_addr(s_axi_6_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_6_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_19_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_19_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_19_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_19_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_19_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_19_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_19_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_19_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_19_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_19_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_20(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_6_w_ready),
		.io_enq_valid(s_axi_6_w_valid),
		.io_enq_bits_data(s_axi_6_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_6_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_20_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_20_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_20_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_20_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_13(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_13_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_6_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_6_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_21(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_7_ar_ready),
		.io_enq_valid(s_axi_7_ar_valid),
		.io_enq_bits_addr(s_axi_7_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_7_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_21_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_21_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_21_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_21_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_21_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_21_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_21_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_21_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_21_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_21_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_14(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_14_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_7_valid),
		.io_enq_bits_data(_read_demux_io_sinks_7_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_7_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_7_bits_last),
		.io_deq_ready(s_axi_7_r_ready),
		.io_deq_valid(s_axi_7_r_valid),
		.io_deq_bits_data(s_axi_7_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_22(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_7_aw_ready),
		.io_enq_valid(s_axi_7_aw_valid),
		.io_enq_bits_addr(s_axi_7_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_7_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_22_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_22_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_22_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_22_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_22_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_22_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_22_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_22_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_22_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_22_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_23(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_7_w_ready),
		.io_enq_valid(s_axi_7_w_valid),
		.io_enq_bits_data(s_axi_7_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_7_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_23_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_23_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_23_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_23_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_15(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_15_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_7_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_7_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_24(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_8_ar_ready),
		.io_enq_valid(s_axi_8_ar_valid),
		.io_enq_bits_addr(s_axi_8_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_8_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_24_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_24_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_24_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_24_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_24_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_24_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_24_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_24_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_24_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_24_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_16(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_16_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_8_valid),
		.io_enq_bits_data(_read_demux_io_sinks_8_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_8_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_8_bits_last),
		.io_deq_ready(s_axi_8_r_ready),
		.io_deq_valid(s_axi_8_r_valid),
		.io_deq_bits_data(s_axi_8_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_25(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_8_aw_ready),
		.io_enq_valid(s_axi_8_aw_valid),
		.io_enq_bits_addr(s_axi_8_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_8_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_25_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_25_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_25_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_25_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_25_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_25_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_25_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_25_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_25_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_25_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_26(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_8_w_ready),
		.io_enq_valid(s_axi_8_w_valid),
		.io_enq_bits_data(s_axi_8_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_8_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_26_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_26_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_26_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_26_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_17(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_17_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_8_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_8_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_27(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_9_ar_ready),
		.io_enq_valid(s_axi_9_ar_valid),
		.io_enq_bits_addr(s_axi_9_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_9_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_27_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_27_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_27_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_27_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_27_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_27_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_27_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_27_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_27_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_27_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_18(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_18_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_9_valid),
		.io_enq_bits_data(_read_demux_io_sinks_9_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_9_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_9_bits_last),
		.io_deq_ready(s_axi_9_r_ready),
		.io_deq_valid(s_axi_9_r_valid),
		.io_deq_bits_data(s_axi_9_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_28(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_9_aw_ready),
		.io_enq_valid(s_axi_9_aw_valid),
		.io_enq_bits_addr(s_axi_9_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_9_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_28_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_28_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_28_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_28_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_28_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_28_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_28_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_28_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_28_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_28_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_29(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_9_w_ready),
		.io_enq_valid(s_axi_9_w_valid),
		.io_enq_bits_data(s_axi_9_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_9_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_29_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_29_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_29_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_29_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_19(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_19_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_9_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_9_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_30(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_10_ar_ready),
		.io_enq_valid(s_axi_10_ar_valid),
		.io_enq_bits_addr(s_axi_10_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_10_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_30_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_30_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_30_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_30_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_30_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_30_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_30_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_30_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_30_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_30_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_20(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_20_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_10_valid),
		.io_enq_bits_data(_read_demux_io_sinks_10_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_10_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_10_bits_last),
		.io_deq_ready(s_axi_10_r_ready),
		.io_deq_valid(s_axi_10_r_valid),
		.io_deq_bits_data(s_axi_10_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_31(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_10_aw_ready),
		.io_enq_valid(s_axi_10_aw_valid),
		.io_enq_bits_addr(s_axi_10_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_10_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_31_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_31_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_31_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_31_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_31_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_31_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_31_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_31_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_31_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_31_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_32(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_10_w_ready),
		.io_enq_valid(s_axi_10_w_valid),
		.io_enq_bits_data(s_axi_10_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_10_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_32_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_32_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_32_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_32_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_21(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_21_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_10_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_10_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_33(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_11_ar_ready),
		.io_enq_valid(s_axi_11_ar_valid),
		.io_enq_bits_addr(s_axi_11_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_11_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_33_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_33_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_33_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_33_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_33_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_33_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_33_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_33_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_33_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_33_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_22(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_22_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_11_valid),
		.io_enq_bits_data(_read_demux_io_sinks_11_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_11_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_11_bits_last),
		.io_deq_ready(s_axi_11_r_ready),
		.io_deq_valid(s_axi_11_r_valid),
		.io_deq_bits_data(s_axi_11_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_34(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_11_aw_ready),
		.io_enq_valid(s_axi_11_aw_valid),
		.io_enq_bits_addr(s_axi_11_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_11_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_34_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_34_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_34_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_34_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_34_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_34_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_34_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_34_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_34_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_34_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_35(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_11_w_ready),
		.io_enq_valid(s_axi_11_w_valid),
		.io_enq_bits_data(s_axi_11_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_11_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_35_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_35_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_35_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_35_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_23(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_23_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_11_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_11_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_36(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_12_ar_ready),
		.io_enq_valid(s_axi_12_ar_valid),
		.io_enq_bits_addr(s_axi_12_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_12_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_36_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_36_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_36_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_36_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_36_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_36_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_36_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_36_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_36_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_36_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_24(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_24_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_12_valid),
		.io_enq_bits_data(_read_demux_io_sinks_12_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_12_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_12_bits_last),
		.io_deq_ready(s_axi_12_r_ready),
		.io_deq_valid(s_axi_12_r_valid),
		.io_deq_bits_data(s_axi_12_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_37(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_12_aw_ready),
		.io_enq_valid(s_axi_12_aw_valid),
		.io_enq_bits_addr(s_axi_12_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_12_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_37_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_37_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_37_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_37_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_37_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_37_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_37_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_37_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_37_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_37_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_38(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_12_w_ready),
		.io_enq_valid(s_axi_12_w_valid),
		.io_enq_bits_data(s_axi_12_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_12_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_38_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_38_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_38_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_38_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_25(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_25_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_12_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_12_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_39(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_13_ar_ready),
		.io_enq_valid(s_axi_13_ar_valid),
		.io_enq_bits_addr(s_axi_13_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_13_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_39_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_39_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_39_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_39_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_39_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_39_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_39_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_39_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_39_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_39_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_26(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_26_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_13_valid),
		.io_enq_bits_data(_read_demux_io_sinks_13_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_13_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_13_bits_last),
		.io_deq_ready(s_axi_13_r_ready),
		.io_deq_valid(s_axi_13_r_valid),
		.io_deq_bits_data(s_axi_13_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_40(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_13_aw_ready),
		.io_enq_valid(s_axi_13_aw_valid),
		.io_enq_bits_addr(s_axi_13_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_13_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_40_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_40_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_40_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_40_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_40_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_40_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_40_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_40_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_40_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_40_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_41(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_13_w_ready),
		.io_enq_valid(s_axi_13_w_valid),
		.io_enq_bits_data(s_axi_13_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_13_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_41_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_41_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_41_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_41_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_27(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_27_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_13_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_13_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_42(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_14_ar_ready),
		.io_enq_valid(s_axi_14_ar_valid),
		.io_enq_bits_addr(s_axi_14_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_14_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_42_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_42_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_42_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_42_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_42_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_42_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_42_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_42_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_42_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_42_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_28(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_28_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_14_valid),
		.io_enq_bits_data(_read_demux_io_sinks_14_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_14_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_14_bits_last),
		.io_deq_ready(s_axi_14_r_ready),
		.io_deq_valid(s_axi_14_r_valid),
		.io_deq_bits_data(s_axi_14_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_43(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_14_aw_ready),
		.io_enq_valid(s_axi_14_aw_valid),
		.io_enq_bits_addr(s_axi_14_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_14_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_43_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_43_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_43_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_43_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_43_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_43_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_43_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_43_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_43_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_43_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_44(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_14_w_ready),
		.io_enq_valid(s_axi_14_w_valid),
		.io_enq_bits_data(s_axi_14_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_14_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_44_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_44_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_44_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_44_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_29(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_29_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_14_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_14_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_45(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_15_ar_ready),
		.io_enq_valid(s_axi_15_ar_valid),
		.io_enq_bits_addr(s_axi_15_ar_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_15_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_45_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_45_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_45_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_45_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_45_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_45_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_45_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_45_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_45_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_45_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_30(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_30_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_15_valid),
		.io_enq_bits_data(_read_demux_io_sinks_15_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_15_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_15_bits_last),
		.io_deq_ready(s_axi_15_r_ready),
		.io_deq_valid(s_axi_15_r_valid),
		.io_deq_bits_data(s_axi_15_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_46(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_15_aw_ready),
		.io_enq_valid(s_axi_15_aw_valid),
		.io_enq_bits_addr(s_axi_15_aw_bits_addr),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h2),
		.io_enq_bits_burst(2'h1),
		.io_deq_ready(_write_arbiter_io_sources_15_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_46_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_46_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_46_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_46_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_46_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_46_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_46_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_46_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_46_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_46_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_47(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_15_w_ready),
		.io_enq_valid(s_axi_15_w_valid),
		.io_enq_bits_data(s_axi_15_w_bits_data),
		.io_enq_bits_strb(4'hf),
		.io_enq_bits_last(1'h1),
		.io_deq_ready(_write_mux_io_sources_15_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_47_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_47_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_47_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_47_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_31(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_31_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_15_valid),
		.io_deq_ready(1'h1),
		.io_deq_valid(s_axi_15_b_valid)
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_48(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_16_ar_ready),
		.io_enq_valid(s_axi_16_ar_valid),
		.io_enq_bits_addr(s_axi_16_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_16_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_48_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_48_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_48_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_48_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_48_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_48_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_48_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_48_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_48_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_48_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_32(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_32_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_16_valid),
		.io_enq_bits_data(_read_demux_io_sinks_16_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_16_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_16_bits_last),
		.io_deq_ready(s_axi_16_r_ready),
		.io_deq_valid(s_axi_16_r_valid),
		.io_deq_bits_data(s_axi_16_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_49(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_16_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_49_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_49_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_49_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_49_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_49_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_49_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_49_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_49_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_49_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_49_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_50(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_16_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_50_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_50_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_50_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_50_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_33(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_33_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_16_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_51(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_17_ar_ready),
		.io_enq_valid(s_axi_17_ar_valid),
		.io_enq_bits_addr(s_axi_17_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_17_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_51_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_51_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_51_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_51_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_51_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_51_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_51_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_51_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_51_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_51_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_34(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_34_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_17_valid),
		.io_enq_bits_data(_read_demux_io_sinks_17_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_17_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_17_bits_last),
		.io_deq_ready(s_axi_17_r_ready),
		.io_deq_valid(s_axi_17_r_valid),
		.io_deq_bits_data(s_axi_17_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_52(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_17_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_52_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_52_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_52_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_52_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_52_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_52_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_52_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_52_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_52_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_52_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_53(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_17_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_53_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_53_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_53_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_53_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_35(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_35_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_17_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_54(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_18_ar_ready),
		.io_enq_valid(s_axi_18_ar_valid),
		.io_enq_bits_addr(s_axi_18_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_18_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_54_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_54_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_54_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_54_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_54_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_54_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_54_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_54_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_54_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_54_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_36(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_36_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_18_valid),
		.io_enq_bits_data(_read_demux_io_sinks_18_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_18_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_18_bits_last),
		.io_deq_ready(s_axi_18_r_ready),
		.io_deq_valid(s_axi_18_r_valid),
		.io_deq_bits_data(s_axi_18_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_55(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_18_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_55_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_55_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_55_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_55_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_55_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_55_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_55_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_55_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_55_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_55_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_56(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_18_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_56_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_56_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_56_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_56_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_37(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_37_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_18_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_57(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_19_ar_ready),
		.io_enq_valid(s_axi_19_ar_valid),
		.io_enq_bits_addr(s_axi_19_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_19_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_57_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_57_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_57_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_57_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_57_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_57_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_57_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_57_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_57_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_57_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_38(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_38_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_19_valid),
		.io_enq_bits_data(_read_demux_io_sinks_19_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_19_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_19_bits_last),
		.io_deq_ready(s_axi_19_r_ready),
		.io_deq_valid(s_axi_19_r_valid),
		.io_deq_bits_data(s_axi_19_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_58(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_19_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_58_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_58_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_58_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_58_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_58_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_58_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_58_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_58_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_58_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_58_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_59(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_19_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_59_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_59_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_59_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_59_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_39(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_39_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_19_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_60(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_20_ar_ready),
		.io_enq_valid(s_axi_20_ar_valid),
		.io_enq_bits_addr(s_axi_20_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_20_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_60_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_60_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_60_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_60_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_60_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_60_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_60_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_60_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_60_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_60_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_40(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_40_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_20_valid),
		.io_enq_bits_data(_read_demux_io_sinks_20_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_20_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_20_bits_last),
		.io_deq_ready(s_axi_20_r_ready),
		.io_deq_valid(s_axi_20_r_valid),
		.io_deq_bits_data(s_axi_20_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_61(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_20_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_61_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_61_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_61_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_61_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_61_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_61_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_61_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_61_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_61_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_61_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_62(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_20_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_62_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_62_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_62_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_62_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_41(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_41_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_20_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_63(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_21_ar_ready),
		.io_enq_valid(s_axi_21_ar_valid),
		.io_enq_bits_addr(s_axi_21_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_21_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_63_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_63_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_63_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_63_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_63_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_63_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_63_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_63_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_63_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_63_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_42(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_42_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_21_valid),
		.io_enq_bits_data(_read_demux_io_sinks_21_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_21_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_21_bits_last),
		.io_deq_ready(s_axi_21_r_ready),
		.io_deq_valid(s_axi_21_r_valid),
		.io_deq_bits_data(s_axi_21_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_64(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_21_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_64_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_64_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_64_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_64_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_64_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_64_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_64_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_64_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_64_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_64_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_65(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_21_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_65_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_65_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_65_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_65_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_43(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_43_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_21_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_66(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_22_ar_ready),
		.io_enq_valid(s_axi_22_ar_valid),
		.io_enq_bits_addr(s_axi_22_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_22_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_66_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_66_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_66_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_66_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_66_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_66_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_66_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_66_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_66_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_66_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_44(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_44_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_22_valid),
		.io_enq_bits_data(_read_demux_io_sinks_22_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_22_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_22_bits_last),
		.io_deq_ready(s_axi_22_r_ready),
		.io_deq_valid(s_axi_22_r_valid),
		.io_deq_bits_data(s_axi_22_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_67(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_22_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_67_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_67_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_67_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_67_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_67_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_67_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_67_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_67_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_67_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_67_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_68(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_22_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_68_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_68_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_68_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_68_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_45(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_45_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_22_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_69(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_23_ar_ready),
		.io_enq_valid(s_axi_23_ar_valid),
		.io_enq_bits_addr(s_axi_23_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_23_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_69_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_69_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_69_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_69_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_69_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_69_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_69_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_69_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_69_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_69_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_46(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_46_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_23_valid),
		.io_enq_bits_data(_read_demux_io_sinks_23_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_23_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_23_bits_last),
		.io_deq_ready(s_axi_23_r_ready),
		.io_deq_valid(s_axi_23_r_valid),
		.io_deq_bits_data(s_axi_23_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_70(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_23_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_70_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_70_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_70_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_70_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_70_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_70_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_70_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_70_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_70_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_70_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_71(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_23_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_71_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_71_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_71_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_71_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_47(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_47_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_23_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_72(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_24_ar_ready),
		.io_enq_valid(s_axi_24_ar_valid),
		.io_enq_bits_addr(s_axi_24_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_24_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_72_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_72_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_72_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_72_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_72_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_72_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_72_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_72_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_72_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_72_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_48(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_48_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_24_valid),
		.io_enq_bits_data(_read_demux_io_sinks_24_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_24_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_24_bits_last),
		.io_deq_ready(s_axi_24_r_ready),
		.io_deq_valid(s_axi_24_r_valid),
		.io_deq_bits_data(s_axi_24_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_73(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_24_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_73_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_73_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_73_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_73_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_73_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_73_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_73_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_73_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_73_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_73_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_74(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_24_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_74_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_74_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_74_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_74_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_49(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_49_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_24_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_75(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_25_ar_ready),
		.io_enq_valid(s_axi_25_ar_valid),
		.io_enq_bits_addr(s_axi_25_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_25_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_75_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_75_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_75_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_75_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_75_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_75_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_75_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_75_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_75_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_75_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_50(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_50_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_25_valid),
		.io_enq_bits_data(_read_demux_io_sinks_25_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_25_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_25_bits_last),
		.io_deq_ready(s_axi_25_r_ready),
		.io_deq_valid(s_axi_25_r_valid),
		.io_deq_bits_data(s_axi_25_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_76(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_25_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_76_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_76_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_76_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_76_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_76_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_76_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_76_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_76_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_76_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_76_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_77(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_25_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_77_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_77_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_77_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_77_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_51(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_51_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_25_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_78(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_26_ar_ready),
		.io_enq_valid(s_axi_26_ar_valid),
		.io_enq_bits_addr(s_axi_26_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_26_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_78_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_78_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_78_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_78_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_78_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_78_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_78_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_78_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_78_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_78_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_52(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_52_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_26_valid),
		.io_enq_bits_data(_read_demux_io_sinks_26_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_26_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_26_bits_last),
		.io_deq_ready(s_axi_26_r_ready),
		.io_deq_valid(s_axi_26_r_valid),
		.io_deq_bits_data(s_axi_26_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_79(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_26_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_79_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_79_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_79_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_79_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_79_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_79_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_79_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_79_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_79_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_79_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_80(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_26_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_80_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_80_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_80_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_80_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_53(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_53_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_26_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_81(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_27_ar_ready),
		.io_enq_valid(s_axi_27_ar_valid),
		.io_enq_bits_addr(s_axi_27_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_27_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_81_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_81_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_81_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_81_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_81_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_81_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_81_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_81_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_81_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_81_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_54(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_54_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_27_valid),
		.io_enq_bits_data(_read_demux_io_sinks_27_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_27_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_27_bits_last),
		.io_deq_ready(s_axi_27_r_ready),
		.io_deq_valid(s_axi_27_r_valid),
		.io_deq_bits_data(s_axi_27_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_82(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_27_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_82_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_82_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_82_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_82_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_82_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_82_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_82_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_82_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_82_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_82_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_83(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_27_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_83_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_83_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_83_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_83_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_55(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_55_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_27_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_84(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_28_ar_ready),
		.io_enq_valid(s_axi_28_ar_valid),
		.io_enq_bits_addr(s_axi_28_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_28_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_84_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_84_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_84_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_84_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_84_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_84_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_84_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_84_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_84_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_84_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_56(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_56_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_28_valid),
		.io_enq_bits_data(_read_demux_io_sinks_28_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_28_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_28_bits_last),
		.io_deq_ready(s_axi_28_r_ready),
		.io_deq_valid(s_axi_28_r_valid),
		.io_deq_bits_data(s_axi_28_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_85(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_28_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_85_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_85_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_85_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_85_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_85_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_85_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_85_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_85_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_85_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_85_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_86(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_28_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_86_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_86_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_86_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_86_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_57(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_57_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_28_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_87(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_29_ar_ready),
		.io_enq_valid(s_axi_29_ar_valid),
		.io_enq_bits_addr(s_axi_29_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_29_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_87_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_87_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_87_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_87_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_87_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_87_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_87_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_87_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_87_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_87_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_58(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_58_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_29_valid),
		.io_enq_bits_data(_read_demux_io_sinks_29_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_29_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_29_bits_last),
		.io_deq_ready(s_axi_29_r_ready),
		.io_deq_valid(s_axi_29_r_valid),
		.io_deq_bits_data(s_axi_29_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_88(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_29_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_88_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_88_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_88_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_88_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_88_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_88_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_88_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_88_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_88_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_88_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_89(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_29_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_89_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_89_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_89_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_89_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_59(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_59_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_29_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_90(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_30_ar_ready),
		.io_enq_valid(s_axi_30_ar_valid),
		.io_enq_bits_addr(s_axi_30_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_30_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_90_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_90_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_90_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_90_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_90_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_90_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_90_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_90_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_90_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_90_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_60(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_60_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_30_valid),
		.io_enq_bits_data(_read_demux_io_sinks_30_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_30_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_30_bits_last),
		.io_deq_ready(s_axi_30_r_ready),
		.io_deq_valid(s_axi_30_r_valid),
		.io_deq_bits_data(s_axi_30_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_91(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_30_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_91_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_91_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_91_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_91_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_91_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_91_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_91_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_91_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_91_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_91_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_92(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_30_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_92_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_92_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_92_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_92_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_61(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_61_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_30_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_1 s_axi__buffered_sourceBuffer_93(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axi_31_ar_ready),
		.io_enq_valid(s_axi_31_ar_valid),
		.io_enq_bits_addr(s_axi_31_ar_bits_addr),
		.io_enq_bits_len(8'h06),
		.io_enq_bits_size(3'h2),
		.io_deq_ready(_read_arbiter_io_sources_31_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_93_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_93_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_93_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_93_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_93_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_93_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_93_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_93_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_93_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_93_io_deq_bits_region)
	);
	Queue2_ReadDataChannel_16 s_axi__buffered_sinkBuffer_62(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_62_io_enq_ready),
		.io_enq_valid(_read_demux_io_sinks_31_valid),
		.io_enq_bits_data(_read_demux_io_sinks_31_bits_data),
		.io_enq_bits_resp(_read_demux_io_sinks_31_bits_resp),
		.io_enq_bits_last(_read_demux_io_sinks_31_bits_last),
		.io_deq_ready(s_axi_31_r_ready),
		.io_deq_valid(s_axi_31_r_valid),
		.io_deq_bits_data(s_axi_31_r_bits_data)
	);
	Queue2_WriteAddressChannel_1 s_axi__buffered_sourceBuffer_94(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_addr(64'h0000000000000000),
		.io_enq_bits_len(8'h00),
		.io_enq_bits_size(3'h0),
		.io_enq_bits_burst(2'h0),
		.io_deq_ready(_write_arbiter_io_sources_31_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_94_io_deq_valid),
		.io_deq_bits_addr(_s_axi__buffered_sourceBuffer_94_io_deq_bits_addr),
		.io_deq_bits_len(_s_axi__buffered_sourceBuffer_94_io_deq_bits_len),
		.io_deq_bits_size(_s_axi__buffered_sourceBuffer_94_io_deq_bits_size),
		.io_deq_bits_burst(_s_axi__buffered_sourceBuffer_94_io_deq_bits_burst),
		.io_deq_bits_lock(_s_axi__buffered_sourceBuffer_94_io_deq_bits_lock),
		.io_deq_bits_cache(_s_axi__buffered_sourceBuffer_94_io_deq_bits_cache),
		.io_deq_bits_prot(_s_axi__buffered_sourceBuffer_94_io_deq_bits_prot),
		.io_deq_bits_qos(_s_axi__buffered_sourceBuffer_94_io_deq_bits_qos),
		.io_deq_bits_region(_s_axi__buffered_sourceBuffer_94_io_deq_bits_region)
	);
	Queue2_WriteDataChannel_16 s_axi__buffered_sourceBuffer_95(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(),
		.io_enq_valid(1'h0),
		.io_enq_bits_data(32'h00000000),
		.io_enq_bits_strb(4'h0),
		.io_enq_bits_last(1'h0),
		.io_deq_ready(_write_mux_io_sources_31_ready),
		.io_deq_valid(_s_axi__buffered_sourceBuffer_95_io_deq_valid),
		.io_deq_bits_data(_s_axi__buffered_sourceBuffer_95_io_deq_bits_data),
		.io_deq_bits_strb(_s_axi__buffered_sourceBuffer_95_io_deq_bits_strb),
		.io_deq_bits_last(_s_axi__buffered_sourceBuffer_95_io_deq_bits_last)
	);
	Queue2_WriteResponseChannel_16 s_axi__buffered_sinkBuffer_63(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axi__buffered_sinkBuffer_63_io_enq_ready),
		.io_enq_valid(_write_demux_io_sinks_31_valid),
		.io_deq_ready(1'h0),
		.io_deq_valid()
	);
	Queue2_ReadAddressChannel_43 m_axi__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_enq_valid(_read_arbiter_io_sink_valid),
		.io_enq_bits_id(_read_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_read_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_read_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_read_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_id(m_axi_ar_bits_id),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	Queue2_ReadDataChannel_48 m_axi__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_r_ready),
		.io_enq_valid(m_axi_r_valid),
		.io_enq_bits_id(m_axi_r_bits_id),
		.io_enq_bits_data(m_axi_r_bits_data),
		.io_enq_bits_resp(m_axi_r_bits_resp),
		.io_enq_bits_last(m_axi_r_bits_last),
		.io_deq_ready(m_axi__r_ready),
		.io_deq_valid(_m_axi__sinkBuffer_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_io_deq_bits_id),
		.io_deq_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_deq_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_deq_bits_last(_m_axi__sinkBuffer_io_deq_bits_last)
	);
	Queue2_WriteAddressChannel_43 m_axi__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_sink_valid),
		.io_enq_bits_id(_write_arbiter_io_sink_bits_id),
		.io_enq_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_enq_bits_len(_write_arbiter_io_sink_bits_len),
		.io_enq_bits_size(_write_arbiter_io_sink_bits_size),
		.io_enq_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_enq_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_enq_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_enq_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_enq_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_enq_bits_region(_write_arbiter_io_sink_bits_region),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_id(m_axi_aw_bits_id),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_WriteDataChannel_16 m_axi__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_enq_valid(_write_mux_io_sink_valid),
		.io_enq_bits_data(_write_mux_io_sink_bits_data),
		.io_enq_bits_strb(_write_mux_io_sink_bits_strb),
		.io_enq_bits_last(_write_mux_io_sink_bits_last),
		.io_deq_ready(m_axi_w_ready),
		.io_deq_valid(m_axi_w_valid),
		.io_deq_bits_data(m_axi_w_bits_data),
		.io_deq_bits_strb(m_axi_w_bits_strb),
		.io_deq_bits_last(m_axi_w_bits_last)
	);
	Queue2_WriteResponseChannel_48 m_axi__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(m_axi_b_ready),
		.io_enq_valid(m_axi_b_valid),
		.io_enq_bits_id(m_axi_b_bits_id),
		.io_enq_bits_resp(m_axi_b_bits_resp),
		.io_deq_ready(m_axi__b_ready),
		.io_deq_valid(_m_axi__sinkBuffer_1_io_deq_valid),
		.io_deq_bits_id(_m_axi__sinkBuffer_1_io_deq_bits_id)
	);
	elasticArbiter_6 read_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_read_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_io_deq_valid),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_io_deq_bits_region),
		.io_sources_1_ready(_read_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_3_io_deq_valid),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_3_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_3_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_3_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_3_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_3_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_3_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_3_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_3_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_3_io_deq_bits_region),
		.io_sources_2_ready(_read_arbiter_io_sources_2_ready),
		.io_sources_2_valid(_s_axi__buffered_sourceBuffer_6_io_deq_valid),
		.io_sources_2_bits_addr(_s_axi__buffered_sourceBuffer_6_io_deq_bits_addr),
		.io_sources_2_bits_len(_s_axi__buffered_sourceBuffer_6_io_deq_bits_len),
		.io_sources_2_bits_size(_s_axi__buffered_sourceBuffer_6_io_deq_bits_size),
		.io_sources_2_bits_burst(_s_axi__buffered_sourceBuffer_6_io_deq_bits_burst),
		.io_sources_2_bits_lock(_s_axi__buffered_sourceBuffer_6_io_deq_bits_lock),
		.io_sources_2_bits_cache(_s_axi__buffered_sourceBuffer_6_io_deq_bits_cache),
		.io_sources_2_bits_prot(_s_axi__buffered_sourceBuffer_6_io_deq_bits_prot),
		.io_sources_2_bits_qos(_s_axi__buffered_sourceBuffer_6_io_deq_bits_qos),
		.io_sources_2_bits_region(_s_axi__buffered_sourceBuffer_6_io_deq_bits_region),
		.io_sources_3_ready(_read_arbiter_io_sources_3_ready),
		.io_sources_3_valid(_s_axi__buffered_sourceBuffer_9_io_deq_valid),
		.io_sources_3_bits_addr(_s_axi__buffered_sourceBuffer_9_io_deq_bits_addr),
		.io_sources_3_bits_len(_s_axi__buffered_sourceBuffer_9_io_deq_bits_len),
		.io_sources_3_bits_size(_s_axi__buffered_sourceBuffer_9_io_deq_bits_size),
		.io_sources_3_bits_burst(_s_axi__buffered_sourceBuffer_9_io_deq_bits_burst),
		.io_sources_3_bits_lock(_s_axi__buffered_sourceBuffer_9_io_deq_bits_lock),
		.io_sources_3_bits_cache(_s_axi__buffered_sourceBuffer_9_io_deq_bits_cache),
		.io_sources_3_bits_prot(_s_axi__buffered_sourceBuffer_9_io_deq_bits_prot),
		.io_sources_3_bits_qos(_s_axi__buffered_sourceBuffer_9_io_deq_bits_qos),
		.io_sources_3_bits_region(_s_axi__buffered_sourceBuffer_9_io_deq_bits_region),
		.io_sources_4_ready(_read_arbiter_io_sources_4_ready),
		.io_sources_4_valid(_s_axi__buffered_sourceBuffer_12_io_deq_valid),
		.io_sources_4_bits_addr(_s_axi__buffered_sourceBuffer_12_io_deq_bits_addr),
		.io_sources_4_bits_len(_s_axi__buffered_sourceBuffer_12_io_deq_bits_len),
		.io_sources_4_bits_size(_s_axi__buffered_sourceBuffer_12_io_deq_bits_size),
		.io_sources_4_bits_burst(_s_axi__buffered_sourceBuffer_12_io_deq_bits_burst),
		.io_sources_4_bits_lock(_s_axi__buffered_sourceBuffer_12_io_deq_bits_lock),
		.io_sources_4_bits_cache(_s_axi__buffered_sourceBuffer_12_io_deq_bits_cache),
		.io_sources_4_bits_prot(_s_axi__buffered_sourceBuffer_12_io_deq_bits_prot),
		.io_sources_4_bits_qos(_s_axi__buffered_sourceBuffer_12_io_deq_bits_qos),
		.io_sources_4_bits_region(_s_axi__buffered_sourceBuffer_12_io_deq_bits_region),
		.io_sources_5_ready(_read_arbiter_io_sources_5_ready),
		.io_sources_5_valid(_s_axi__buffered_sourceBuffer_15_io_deq_valid),
		.io_sources_5_bits_addr(_s_axi__buffered_sourceBuffer_15_io_deq_bits_addr),
		.io_sources_5_bits_len(_s_axi__buffered_sourceBuffer_15_io_deq_bits_len),
		.io_sources_5_bits_size(_s_axi__buffered_sourceBuffer_15_io_deq_bits_size),
		.io_sources_5_bits_burst(_s_axi__buffered_sourceBuffer_15_io_deq_bits_burst),
		.io_sources_5_bits_lock(_s_axi__buffered_sourceBuffer_15_io_deq_bits_lock),
		.io_sources_5_bits_cache(_s_axi__buffered_sourceBuffer_15_io_deq_bits_cache),
		.io_sources_5_bits_prot(_s_axi__buffered_sourceBuffer_15_io_deq_bits_prot),
		.io_sources_5_bits_qos(_s_axi__buffered_sourceBuffer_15_io_deq_bits_qos),
		.io_sources_5_bits_region(_s_axi__buffered_sourceBuffer_15_io_deq_bits_region),
		.io_sources_6_ready(_read_arbiter_io_sources_6_ready),
		.io_sources_6_valid(_s_axi__buffered_sourceBuffer_18_io_deq_valid),
		.io_sources_6_bits_addr(_s_axi__buffered_sourceBuffer_18_io_deq_bits_addr),
		.io_sources_6_bits_len(_s_axi__buffered_sourceBuffer_18_io_deq_bits_len),
		.io_sources_6_bits_size(_s_axi__buffered_sourceBuffer_18_io_deq_bits_size),
		.io_sources_6_bits_burst(_s_axi__buffered_sourceBuffer_18_io_deq_bits_burst),
		.io_sources_6_bits_lock(_s_axi__buffered_sourceBuffer_18_io_deq_bits_lock),
		.io_sources_6_bits_cache(_s_axi__buffered_sourceBuffer_18_io_deq_bits_cache),
		.io_sources_6_bits_prot(_s_axi__buffered_sourceBuffer_18_io_deq_bits_prot),
		.io_sources_6_bits_qos(_s_axi__buffered_sourceBuffer_18_io_deq_bits_qos),
		.io_sources_6_bits_region(_s_axi__buffered_sourceBuffer_18_io_deq_bits_region),
		.io_sources_7_ready(_read_arbiter_io_sources_7_ready),
		.io_sources_7_valid(_s_axi__buffered_sourceBuffer_21_io_deq_valid),
		.io_sources_7_bits_addr(_s_axi__buffered_sourceBuffer_21_io_deq_bits_addr),
		.io_sources_7_bits_len(_s_axi__buffered_sourceBuffer_21_io_deq_bits_len),
		.io_sources_7_bits_size(_s_axi__buffered_sourceBuffer_21_io_deq_bits_size),
		.io_sources_7_bits_burst(_s_axi__buffered_sourceBuffer_21_io_deq_bits_burst),
		.io_sources_7_bits_lock(_s_axi__buffered_sourceBuffer_21_io_deq_bits_lock),
		.io_sources_7_bits_cache(_s_axi__buffered_sourceBuffer_21_io_deq_bits_cache),
		.io_sources_7_bits_prot(_s_axi__buffered_sourceBuffer_21_io_deq_bits_prot),
		.io_sources_7_bits_qos(_s_axi__buffered_sourceBuffer_21_io_deq_bits_qos),
		.io_sources_7_bits_region(_s_axi__buffered_sourceBuffer_21_io_deq_bits_region),
		.io_sources_8_ready(_read_arbiter_io_sources_8_ready),
		.io_sources_8_valid(_s_axi__buffered_sourceBuffer_24_io_deq_valid),
		.io_sources_8_bits_addr(_s_axi__buffered_sourceBuffer_24_io_deq_bits_addr),
		.io_sources_8_bits_len(_s_axi__buffered_sourceBuffer_24_io_deq_bits_len),
		.io_sources_8_bits_size(_s_axi__buffered_sourceBuffer_24_io_deq_bits_size),
		.io_sources_8_bits_burst(_s_axi__buffered_sourceBuffer_24_io_deq_bits_burst),
		.io_sources_8_bits_lock(_s_axi__buffered_sourceBuffer_24_io_deq_bits_lock),
		.io_sources_8_bits_cache(_s_axi__buffered_sourceBuffer_24_io_deq_bits_cache),
		.io_sources_8_bits_prot(_s_axi__buffered_sourceBuffer_24_io_deq_bits_prot),
		.io_sources_8_bits_qos(_s_axi__buffered_sourceBuffer_24_io_deq_bits_qos),
		.io_sources_8_bits_region(_s_axi__buffered_sourceBuffer_24_io_deq_bits_region),
		.io_sources_9_ready(_read_arbiter_io_sources_9_ready),
		.io_sources_9_valid(_s_axi__buffered_sourceBuffer_27_io_deq_valid),
		.io_sources_9_bits_addr(_s_axi__buffered_sourceBuffer_27_io_deq_bits_addr),
		.io_sources_9_bits_len(_s_axi__buffered_sourceBuffer_27_io_deq_bits_len),
		.io_sources_9_bits_size(_s_axi__buffered_sourceBuffer_27_io_deq_bits_size),
		.io_sources_9_bits_burst(_s_axi__buffered_sourceBuffer_27_io_deq_bits_burst),
		.io_sources_9_bits_lock(_s_axi__buffered_sourceBuffer_27_io_deq_bits_lock),
		.io_sources_9_bits_cache(_s_axi__buffered_sourceBuffer_27_io_deq_bits_cache),
		.io_sources_9_bits_prot(_s_axi__buffered_sourceBuffer_27_io_deq_bits_prot),
		.io_sources_9_bits_qos(_s_axi__buffered_sourceBuffer_27_io_deq_bits_qos),
		.io_sources_9_bits_region(_s_axi__buffered_sourceBuffer_27_io_deq_bits_region),
		.io_sources_10_ready(_read_arbiter_io_sources_10_ready),
		.io_sources_10_valid(_s_axi__buffered_sourceBuffer_30_io_deq_valid),
		.io_sources_10_bits_addr(_s_axi__buffered_sourceBuffer_30_io_deq_bits_addr),
		.io_sources_10_bits_len(_s_axi__buffered_sourceBuffer_30_io_deq_bits_len),
		.io_sources_10_bits_size(_s_axi__buffered_sourceBuffer_30_io_deq_bits_size),
		.io_sources_10_bits_burst(_s_axi__buffered_sourceBuffer_30_io_deq_bits_burst),
		.io_sources_10_bits_lock(_s_axi__buffered_sourceBuffer_30_io_deq_bits_lock),
		.io_sources_10_bits_cache(_s_axi__buffered_sourceBuffer_30_io_deq_bits_cache),
		.io_sources_10_bits_prot(_s_axi__buffered_sourceBuffer_30_io_deq_bits_prot),
		.io_sources_10_bits_qos(_s_axi__buffered_sourceBuffer_30_io_deq_bits_qos),
		.io_sources_10_bits_region(_s_axi__buffered_sourceBuffer_30_io_deq_bits_region),
		.io_sources_11_ready(_read_arbiter_io_sources_11_ready),
		.io_sources_11_valid(_s_axi__buffered_sourceBuffer_33_io_deq_valid),
		.io_sources_11_bits_addr(_s_axi__buffered_sourceBuffer_33_io_deq_bits_addr),
		.io_sources_11_bits_len(_s_axi__buffered_sourceBuffer_33_io_deq_bits_len),
		.io_sources_11_bits_size(_s_axi__buffered_sourceBuffer_33_io_deq_bits_size),
		.io_sources_11_bits_burst(_s_axi__buffered_sourceBuffer_33_io_deq_bits_burst),
		.io_sources_11_bits_lock(_s_axi__buffered_sourceBuffer_33_io_deq_bits_lock),
		.io_sources_11_bits_cache(_s_axi__buffered_sourceBuffer_33_io_deq_bits_cache),
		.io_sources_11_bits_prot(_s_axi__buffered_sourceBuffer_33_io_deq_bits_prot),
		.io_sources_11_bits_qos(_s_axi__buffered_sourceBuffer_33_io_deq_bits_qos),
		.io_sources_11_bits_region(_s_axi__buffered_sourceBuffer_33_io_deq_bits_region),
		.io_sources_12_ready(_read_arbiter_io_sources_12_ready),
		.io_sources_12_valid(_s_axi__buffered_sourceBuffer_36_io_deq_valid),
		.io_sources_12_bits_addr(_s_axi__buffered_sourceBuffer_36_io_deq_bits_addr),
		.io_sources_12_bits_len(_s_axi__buffered_sourceBuffer_36_io_deq_bits_len),
		.io_sources_12_bits_size(_s_axi__buffered_sourceBuffer_36_io_deq_bits_size),
		.io_sources_12_bits_burst(_s_axi__buffered_sourceBuffer_36_io_deq_bits_burst),
		.io_sources_12_bits_lock(_s_axi__buffered_sourceBuffer_36_io_deq_bits_lock),
		.io_sources_12_bits_cache(_s_axi__buffered_sourceBuffer_36_io_deq_bits_cache),
		.io_sources_12_bits_prot(_s_axi__buffered_sourceBuffer_36_io_deq_bits_prot),
		.io_sources_12_bits_qos(_s_axi__buffered_sourceBuffer_36_io_deq_bits_qos),
		.io_sources_12_bits_region(_s_axi__buffered_sourceBuffer_36_io_deq_bits_region),
		.io_sources_13_ready(_read_arbiter_io_sources_13_ready),
		.io_sources_13_valid(_s_axi__buffered_sourceBuffer_39_io_deq_valid),
		.io_sources_13_bits_addr(_s_axi__buffered_sourceBuffer_39_io_deq_bits_addr),
		.io_sources_13_bits_len(_s_axi__buffered_sourceBuffer_39_io_deq_bits_len),
		.io_sources_13_bits_size(_s_axi__buffered_sourceBuffer_39_io_deq_bits_size),
		.io_sources_13_bits_burst(_s_axi__buffered_sourceBuffer_39_io_deq_bits_burst),
		.io_sources_13_bits_lock(_s_axi__buffered_sourceBuffer_39_io_deq_bits_lock),
		.io_sources_13_bits_cache(_s_axi__buffered_sourceBuffer_39_io_deq_bits_cache),
		.io_sources_13_bits_prot(_s_axi__buffered_sourceBuffer_39_io_deq_bits_prot),
		.io_sources_13_bits_qos(_s_axi__buffered_sourceBuffer_39_io_deq_bits_qos),
		.io_sources_13_bits_region(_s_axi__buffered_sourceBuffer_39_io_deq_bits_region),
		.io_sources_14_ready(_read_arbiter_io_sources_14_ready),
		.io_sources_14_valid(_s_axi__buffered_sourceBuffer_42_io_deq_valid),
		.io_sources_14_bits_addr(_s_axi__buffered_sourceBuffer_42_io_deq_bits_addr),
		.io_sources_14_bits_len(_s_axi__buffered_sourceBuffer_42_io_deq_bits_len),
		.io_sources_14_bits_size(_s_axi__buffered_sourceBuffer_42_io_deq_bits_size),
		.io_sources_14_bits_burst(_s_axi__buffered_sourceBuffer_42_io_deq_bits_burst),
		.io_sources_14_bits_lock(_s_axi__buffered_sourceBuffer_42_io_deq_bits_lock),
		.io_sources_14_bits_cache(_s_axi__buffered_sourceBuffer_42_io_deq_bits_cache),
		.io_sources_14_bits_prot(_s_axi__buffered_sourceBuffer_42_io_deq_bits_prot),
		.io_sources_14_bits_qos(_s_axi__buffered_sourceBuffer_42_io_deq_bits_qos),
		.io_sources_14_bits_region(_s_axi__buffered_sourceBuffer_42_io_deq_bits_region),
		.io_sources_15_ready(_read_arbiter_io_sources_15_ready),
		.io_sources_15_valid(_s_axi__buffered_sourceBuffer_45_io_deq_valid),
		.io_sources_15_bits_addr(_s_axi__buffered_sourceBuffer_45_io_deq_bits_addr),
		.io_sources_15_bits_len(_s_axi__buffered_sourceBuffer_45_io_deq_bits_len),
		.io_sources_15_bits_size(_s_axi__buffered_sourceBuffer_45_io_deq_bits_size),
		.io_sources_15_bits_burst(_s_axi__buffered_sourceBuffer_45_io_deq_bits_burst),
		.io_sources_15_bits_lock(_s_axi__buffered_sourceBuffer_45_io_deq_bits_lock),
		.io_sources_15_bits_cache(_s_axi__buffered_sourceBuffer_45_io_deq_bits_cache),
		.io_sources_15_bits_prot(_s_axi__buffered_sourceBuffer_45_io_deq_bits_prot),
		.io_sources_15_bits_qos(_s_axi__buffered_sourceBuffer_45_io_deq_bits_qos),
		.io_sources_15_bits_region(_s_axi__buffered_sourceBuffer_45_io_deq_bits_region),
		.io_sources_16_ready(_read_arbiter_io_sources_16_ready),
		.io_sources_16_valid(_s_axi__buffered_sourceBuffer_48_io_deq_valid),
		.io_sources_16_bits_addr(_s_axi__buffered_sourceBuffer_48_io_deq_bits_addr),
		.io_sources_16_bits_len(_s_axi__buffered_sourceBuffer_48_io_deq_bits_len),
		.io_sources_16_bits_size(_s_axi__buffered_sourceBuffer_48_io_deq_bits_size),
		.io_sources_16_bits_burst(_s_axi__buffered_sourceBuffer_48_io_deq_bits_burst),
		.io_sources_16_bits_lock(_s_axi__buffered_sourceBuffer_48_io_deq_bits_lock),
		.io_sources_16_bits_cache(_s_axi__buffered_sourceBuffer_48_io_deq_bits_cache),
		.io_sources_16_bits_prot(_s_axi__buffered_sourceBuffer_48_io_deq_bits_prot),
		.io_sources_16_bits_qos(_s_axi__buffered_sourceBuffer_48_io_deq_bits_qos),
		.io_sources_16_bits_region(_s_axi__buffered_sourceBuffer_48_io_deq_bits_region),
		.io_sources_17_ready(_read_arbiter_io_sources_17_ready),
		.io_sources_17_valid(_s_axi__buffered_sourceBuffer_51_io_deq_valid),
		.io_sources_17_bits_addr(_s_axi__buffered_sourceBuffer_51_io_deq_bits_addr),
		.io_sources_17_bits_len(_s_axi__buffered_sourceBuffer_51_io_deq_bits_len),
		.io_sources_17_bits_size(_s_axi__buffered_sourceBuffer_51_io_deq_bits_size),
		.io_sources_17_bits_burst(_s_axi__buffered_sourceBuffer_51_io_deq_bits_burst),
		.io_sources_17_bits_lock(_s_axi__buffered_sourceBuffer_51_io_deq_bits_lock),
		.io_sources_17_bits_cache(_s_axi__buffered_sourceBuffer_51_io_deq_bits_cache),
		.io_sources_17_bits_prot(_s_axi__buffered_sourceBuffer_51_io_deq_bits_prot),
		.io_sources_17_bits_qos(_s_axi__buffered_sourceBuffer_51_io_deq_bits_qos),
		.io_sources_17_bits_region(_s_axi__buffered_sourceBuffer_51_io_deq_bits_region),
		.io_sources_18_ready(_read_arbiter_io_sources_18_ready),
		.io_sources_18_valid(_s_axi__buffered_sourceBuffer_54_io_deq_valid),
		.io_sources_18_bits_addr(_s_axi__buffered_sourceBuffer_54_io_deq_bits_addr),
		.io_sources_18_bits_len(_s_axi__buffered_sourceBuffer_54_io_deq_bits_len),
		.io_sources_18_bits_size(_s_axi__buffered_sourceBuffer_54_io_deq_bits_size),
		.io_sources_18_bits_burst(_s_axi__buffered_sourceBuffer_54_io_deq_bits_burst),
		.io_sources_18_bits_lock(_s_axi__buffered_sourceBuffer_54_io_deq_bits_lock),
		.io_sources_18_bits_cache(_s_axi__buffered_sourceBuffer_54_io_deq_bits_cache),
		.io_sources_18_bits_prot(_s_axi__buffered_sourceBuffer_54_io_deq_bits_prot),
		.io_sources_18_bits_qos(_s_axi__buffered_sourceBuffer_54_io_deq_bits_qos),
		.io_sources_18_bits_region(_s_axi__buffered_sourceBuffer_54_io_deq_bits_region),
		.io_sources_19_ready(_read_arbiter_io_sources_19_ready),
		.io_sources_19_valid(_s_axi__buffered_sourceBuffer_57_io_deq_valid),
		.io_sources_19_bits_addr(_s_axi__buffered_sourceBuffer_57_io_deq_bits_addr),
		.io_sources_19_bits_len(_s_axi__buffered_sourceBuffer_57_io_deq_bits_len),
		.io_sources_19_bits_size(_s_axi__buffered_sourceBuffer_57_io_deq_bits_size),
		.io_sources_19_bits_burst(_s_axi__buffered_sourceBuffer_57_io_deq_bits_burst),
		.io_sources_19_bits_lock(_s_axi__buffered_sourceBuffer_57_io_deq_bits_lock),
		.io_sources_19_bits_cache(_s_axi__buffered_sourceBuffer_57_io_deq_bits_cache),
		.io_sources_19_bits_prot(_s_axi__buffered_sourceBuffer_57_io_deq_bits_prot),
		.io_sources_19_bits_qos(_s_axi__buffered_sourceBuffer_57_io_deq_bits_qos),
		.io_sources_19_bits_region(_s_axi__buffered_sourceBuffer_57_io_deq_bits_region),
		.io_sources_20_ready(_read_arbiter_io_sources_20_ready),
		.io_sources_20_valid(_s_axi__buffered_sourceBuffer_60_io_deq_valid),
		.io_sources_20_bits_addr(_s_axi__buffered_sourceBuffer_60_io_deq_bits_addr),
		.io_sources_20_bits_len(_s_axi__buffered_sourceBuffer_60_io_deq_bits_len),
		.io_sources_20_bits_size(_s_axi__buffered_sourceBuffer_60_io_deq_bits_size),
		.io_sources_20_bits_burst(_s_axi__buffered_sourceBuffer_60_io_deq_bits_burst),
		.io_sources_20_bits_lock(_s_axi__buffered_sourceBuffer_60_io_deq_bits_lock),
		.io_sources_20_bits_cache(_s_axi__buffered_sourceBuffer_60_io_deq_bits_cache),
		.io_sources_20_bits_prot(_s_axi__buffered_sourceBuffer_60_io_deq_bits_prot),
		.io_sources_20_bits_qos(_s_axi__buffered_sourceBuffer_60_io_deq_bits_qos),
		.io_sources_20_bits_region(_s_axi__buffered_sourceBuffer_60_io_deq_bits_region),
		.io_sources_21_ready(_read_arbiter_io_sources_21_ready),
		.io_sources_21_valid(_s_axi__buffered_sourceBuffer_63_io_deq_valid),
		.io_sources_21_bits_addr(_s_axi__buffered_sourceBuffer_63_io_deq_bits_addr),
		.io_sources_21_bits_len(_s_axi__buffered_sourceBuffer_63_io_deq_bits_len),
		.io_sources_21_bits_size(_s_axi__buffered_sourceBuffer_63_io_deq_bits_size),
		.io_sources_21_bits_burst(_s_axi__buffered_sourceBuffer_63_io_deq_bits_burst),
		.io_sources_21_bits_lock(_s_axi__buffered_sourceBuffer_63_io_deq_bits_lock),
		.io_sources_21_bits_cache(_s_axi__buffered_sourceBuffer_63_io_deq_bits_cache),
		.io_sources_21_bits_prot(_s_axi__buffered_sourceBuffer_63_io_deq_bits_prot),
		.io_sources_21_bits_qos(_s_axi__buffered_sourceBuffer_63_io_deq_bits_qos),
		.io_sources_21_bits_region(_s_axi__buffered_sourceBuffer_63_io_deq_bits_region),
		.io_sources_22_ready(_read_arbiter_io_sources_22_ready),
		.io_sources_22_valid(_s_axi__buffered_sourceBuffer_66_io_deq_valid),
		.io_sources_22_bits_addr(_s_axi__buffered_sourceBuffer_66_io_deq_bits_addr),
		.io_sources_22_bits_len(_s_axi__buffered_sourceBuffer_66_io_deq_bits_len),
		.io_sources_22_bits_size(_s_axi__buffered_sourceBuffer_66_io_deq_bits_size),
		.io_sources_22_bits_burst(_s_axi__buffered_sourceBuffer_66_io_deq_bits_burst),
		.io_sources_22_bits_lock(_s_axi__buffered_sourceBuffer_66_io_deq_bits_lock),
		.io_sources_22_bits_cache(_s_axi__buffered_sourceBuffer_66_io_deq_bits_cache),
		.io_sources_22_bits_prot(_s_axi__buffered_sourceBuffer_66_io_deq_bits_prot),
		.io_sources_22_bits_qos(_s_axi__buffered_sourceBuffer_66_io_deq_bits_qos),
		.io_sources_22_bits_region(_s_axi__buffered_sourceBuffer_66_io_deq_bits_region),
		.io_sources_23_ready(_read_arbiter_io_sources_23_ready),
		.io_sources_23_valid(_s_axi__buffered_sourceBuffer_69_io_deq_valid),
		.io_sources_23_bits_addr(_s_axi__buffered_sourceBuffer_69_io_deq_bits_addr),
		.io_sources_23_bits_len(_s_axi__buffered_sourceBuffer_69_io_deq_bits_len),
		.io_sources_23_bits_size(_s_axi__buffered_sourceBuffer_69_io_deq_bits_size),
		.io_sources_23_bits_burst(_s_axi__buffered_sourceBuffer_69_io_deq_bits_burst),
		.io_sources_23_bits_lock(_s_axi__buffered_sourceBuffer_69_io_deq_bits_lock),
		.io_sources_23_bits_cache(_s_axi__buffered_sourceBuffer_69_io_deq_bits_cache),
		.io_sources_23_bits_prot(_s_axi__buffered_sourceBuffer_69_io_deq_bits_prot),
		.io_sources_23_bits_qos(_s_axi__buffered_sourceBuffer_69_io_deq_bits_qos),
		.io_sources_23_bits_region(_s_axi__buffered_sourceBuffer_69_io_deq_bits_region),
		.io_sources_24_ready(_read_arbiter_io_sources_24_ready),
		.io_sources_24_valid(_s_axi__buffered_sourceBuffer_72_io_deq_valid),
		.io_sources_24_bits_addr(_s_axi__buffered_sourceBuffer_72_io_deq_bits_addr),
		.io_sources_24_bits_len(_s_axi__buffered_sourceBuffer_72_io_deq_bits_len),
		.io_sources_24_bits_size(_s_axi__buffered_sourceBuffer_72_io_deq_bits_size),
		.io_sources_24_bits_burst(_s_axi__buffered_sourceBuffer_72_io_deq_bits_burst),
		.io_sources_24_bits_lock(_s_axi__buffered_sourceBuffer_72_io_deq_bits_lock),
		.io_sources_24_bits_cache(_s_axi__buffered_sourceBuffer_72_io_deq_bits_cache),
		.io_sources_24_bits_prot(_s_axi__buffered_sourceBuffer_72_io_deq_bits_prot),
		.io_sources_24_bits_qos(_s_axi__buffered_sourceBuffer_72_io_deq_bits_qos),
		.io_sources_24_bits_region(_s_axi__buffered_sourceBuffer_72_io_deq_bits_region),
		.io_sources_25_ready(_read_arbiter_io_sources_25_ready),
		.io_sources_25_valid(_s_axi__buffered_sourceBuffer_75_io_deq_valid),
		.io_sources_25_bits_addr(_s_axi__buffered_sourceBuffer_75_io_deq_bits_addr),
		.io_sources_25_bits_len(_s_axi__buffered_sourceBuffer_75_io_deq_bits_len),
		.io_sources_25_bits_size(_s_axi__buffered_sourceBuffer_75_io_deq_bits_size),
		.io_sources_25_bits_burst(_s_axi__buffered_sourceBuffer_75_io_deq_bits_burst),
		.io_sources_25_bits_lock(_s_axi__buffered_sourceBuffer_75_io_deq_bits_lock),
		.io_sources_25_bits_cache(_s_axi__buffered_sourceBuffer_75_io_deq_bits_cache),
		.io_sources_25_bits_prot(_s_axi__buffered_sourceBuffer_75_io_deq_bits_prot),
		.io_sources_25_bits_qos(_s_axi__buffered_sourceBuffer_75_io_deq_bits_qos),
		.io_sources_25_bits_region(_s_axi__buffered_sourceBuffer_75_io_deq_bits_region),
		.io_sources_26_ready(_read_arbiter_io_sources_26_ready),
		.io_sources_26_valid(_s_axi__buffered_sourceBuffer_78_io_deq_valid),
		.io_sources_26_bits_addr(_s_axi__buffered_sourceBuffer_78_io_deq_bits_addr),
		.io_sources_26_bits_len(_s_axi__buffered_sourceBuffer_78_io_deq_bits_len),
		.io_sources_26_bits_size(_s_axi__buffered_sourceBuffer_78_io_deq_bits_size),
		.io_sources_26_bits_burst(_s_axi__buffered_sourceBuffer_78_io_deq_bits_burst),
		.io_sources_26_bits_lock(_s_axi__buffered_sourceBuffer_78_io_deq_bits_lock),
		.io_sources_26_bits_cache(_s_axi__buffered_sourceBuffer_78_io_deq_bits_cache),
		.io_sources_26_bits_prot(_s_axi__buffered_sourceBuffer_78_io_deq_bits_prot),
		.io_sources_26_bits_qos(_s_axi__buffered_sourceBuffer_78_io_deq_bits_qos),
		.io_sources_26_bits_region(_s_axi__buffered_sourceBuffer_78_io_deq_bits_region),
		.io_sources_27_ready(_read_arbiter_io_sources_27_ready),
		.io_sources_27_valid(_s_axi__buffered_sourceBuffer_81_io_deq_valid),
		.io_sources_27_bits_addr(_s_axi__buffered_sourceBuffer_81_io_deq_bits_addr),
		.io_sources_27_bits_len(_s_axi__buffered_sourceBuffer_81_io_deq_bits_len),
		.io_sources_27_bits_size(_s_axi__buffered_sourceBuffer_81_io_deq_bits_size),
		.io_sources_27_bits_burst(_s_axi__buffered_sourceBuffer_81_io_deq_bits_burst),
		.io_sources_27_bits_lock(_s_axi__buffered_sourceBuffer_81_io_deq_bits_lock),
		.io_sources_27_bits_cache(_s_axi__buffered_sourceBuffer_81_io_deq_bits_cache),
		.io_sources_27_bits_prot(_s_axi__buffered_sourceBuffer_81_io_deq_bits_prot),
		.io_sources_27_bits_qos(_s_axi__buffered_sourceBuffer_81_io_deq_bits_qos),
		.io_sources_27_bits_region(_s_axi__buffered_sourceBuffer_81_io_deq_bits_region),
		.io_sources_28_ready(_read_arbiter_io_sources_28_ready),
		.io_sources_28_valid(_s_axi__buffered_sourceBuffer_84_io_deq_valid),
		.io_sources_28_bits_addr(_s_axi__buffered_sourceBuffer_84_io_deq_bits_addr),
		.io_sources_28_bits_len(_s_axi__buffered_sourceBuffer_84_io_deq_bits_len),
		.io_sources_28_bits_size(_s_axi__buffered_sourceBuffer_84_io_deq_bits_size),
		.io_sources_28_bits_burst(_s_axi__buffered_sourceBuffer_84_io_deq_bits_burst),
		.io_sources_28_bits_lock(_s_axi__buffered_sourceBuffer_84_io_deq_bits_lock),
		.io_sources_28_bits_cache(_s_axi__buffered_sourceBuffer_84_io_deq_bits_cache),
		.io_sources_28_bits_prot(_s_axi__buffered_sourceBuffer_84_io_deq_bits_prot),
		.io_sources_28_bits_qos(_s_axi__buffered_sourceBuffer_84_io_deq_bits_qos),
		.io_sources_28_bits_region(_s_axi__buffered_sourceBuffer_84_io_deq_bits_region),
		.io_sources_29_ready(_read_arbiter_io_sources_29_ready),
		.io_sources_29_valid(_s_axi__buffered_sourceBuffer_87_io_deq_valid),
		.io_sources_29_bits_addr(_s_axi__buffered_sourceBuffer_87_io_deq_bits_addr),
		.io_sources_29_bits_len(_s_axi__buffered_sourceBuffer_87_io_deq_bits_len),
		.io_sources_29_bits_size(_s_axi__buffered_sourceBuffer_87_io_deq_bits_size),
		.io_sources_29_bits_burst(_s_axi__buffered_sourceBuffer_87_io_deq_bits_burst),
		.io_sources_29_bits_lock(_s_axi__buffered_sourceBuffer_87_io_deq_bits_lock),
		.io_sources_29_bits_cache(_s_axi__buffered_sourceBuffer_87_io_deq_bits_cache),
		.io_sources_29_bits_prot(_s_axi__buffered_sourceBuffer_87_io_deq_bits_prot),
		.io_sources_29_bits_qos(_s_axi__buffered_sourceBuffer_87_io_deq_bits_qos),
		.io_sources_29_bits_region(_s_axi__buffered_sourceBuffer_87_io_deq_bits_region),
		.io_sources_30_ready(_read_arbiter_io_sources_30_ready),
		.io_sources_30_valid(_s_axi__buffered_sourceBuffer_90_io_deq_valid),
		.io_sources_30_bits_addr(_s_axi__buffered_sourceBuffer_90_io_deq_bits_addr),
		.io_sources_30_bits_len(_s_axi__buffered_sourceBuffer_90_io_deq_bits_len),
		.io_sources_30_bits_size(_s_axi__buffered_sourceBuffer_90_io_deq_bits_size),
		.io_sources_30_bits_burst(_s_axi__buffered_sourceBuffer_90_io_deq_bits_burst),
		.io_sources_30_bits_lock(_s_axi__buffered_sourceBuffer_90_io_deq_bits_lock),
		.io_sources_30_bits_cache(_s_axi__buffered_sourceBuffer_90_io_deq_bits_cache),
		.io_sources_30_bits_prot(_s_axi__buffered_sourceBuffer_90_io_deq_bits_prot),
		.io_sources_30_bits_qos(_s_axi__buffered_sourceBuffer_90_io_deq_bits_qos),
		.io_sources_30_bits_region(_s_axi__buffered_sourceBuffer_90_io_deq_bits_region),
		.io_sources_31_ready(_read_arbiter_io_sources_31_ready),
		.io_sources_31_valid(_s_axi__buffered_sourceBuffer_93_io_deq_valid),
		.io_sources_31_bits_addr(_s_axi__buffered_sourceBuffer_93_io_deq_bits_addr),
		.io_sources_31_bits_len(_s_axi__buffered_sourceBuffer_93_io_deq_bits_len),
		.io_sources_31_bits_size(_s_axi__buffered_sourceBuffer_93_io_deq_bits_size),
		.io_sources_31_bits_burst(_s_axi__buffered_sourceBuffer_93_io_deq_bits_burst),
		.io_sources_31_bits_lock(_s_axi__buffered_sourceBuffer_93_io_deq_bits_lock),
		.io_sources_31_bits_cache(_s_axi__buffered_sourceBuffer_93_io_deq_bits_cache),
		.io_sources_31_bits_prot(_s_axi__buffered_sourceBuffer_93_io_deq_bits_prot),
		.io_sources_31_bits_qos(_s_axi__buffered_sourceBuffer_93_io_deq_bits_qos),
		.io_sources_31_bits_region(_s_axi__buffered_sourceBuffer_93_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_io_enq_ready),
		.io_sink_valid(_read_arbiter_io_sink_valid),
		.io_sink_bits_id(_read_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_read_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_read_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_read_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_read_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_read_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_read_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_read_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_read_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_read_arbiter_io_sink_bits_region),
		.io_select_ready(1'h1),
		.io_select_valid(),
		.io_select_bits()
	);
	elasticDemux_9 read_demux(
		.io_source_ready(_read_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_0),
		.io_source_bits_data(_m_axi__sinkBuffer_io_deq_bits_data),
		.io_source_bits_resp(_m_axi__sinkBuffer_io_deq_bits_resp),
		.io_source_bits_last(_m_axi__sinkBuffer_io_deq_bits_last),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_io_enq_ready),
		.io_sinks_0_valid(_read_demux_io_sinks_0_valid),
		.io_sinks_0_bits_data(_read_demux_io_sinks_0_bits_data),
		.io_sinks_0_bits_resp(_read_demux_io_sinks_0_bits_resp),
		.io_sinks_0_bits_last(_read_demux_io_sinks_0_bits_last),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_2_io_enq_ready),
		.io_sinks_1_valid(_read_demux_io_sinks_1_valid),
		.io_sinks_1_bits_data(_read_demux_io_sinks_1_bits_data),
		.io_sinks_1_bits_resp(_read_demux_io_sinks_1_bits_resp),
		.io_sinks_1_bits_last(_read_demux_io_sinks_1_bits_last),
		.io_sinks_2_ready(_s_axi__buffered_sinkBuffer_4_io_enq_ready),
		.io_sinks_2_valid(_read_demux_io_sinks_2_valid),
		.io_sinks_2_bits_data(_read_demux_io_sinks_2_bits_data),
		.io_sinks_2_bits_resp(_read_demux_io_sinks_2_bits_resp),
		.io_sinks_2_bits_last(_read_demux_io_sinks_2_bits_last),
		.io_sinks_3_ready(_s_axi__buffered_sinkBuffer_6_io_enq_ready),
		.io_sinks_3_valid(_read_demux_io_sinks_3_valid),
		.io_sinks_3_bits_data(_read_demux_io_sinks_3_bits_data),
		.io_sinks_3_bits_resp(_read_demux_io_sinks_3_bits_resp),
		.io_sinks_3_bits_last(_read_demux_io_sinks_3_bits_last),
		.io_sinks_4_ready(_s_axi__buffered_sinkBuffer_8_io_enq_ready),
		.io_sinks_4_valid(_read_demux_io_sinks_4_valid),
		.io_sinks_4_bits_data(_read_demux_io_sinks_4_bits_data),
		.io_sinks_4_bits_resp(_read_demux_io_sinks_4_bits_resp),
		.io_sinks_4_bits_last(_read_demux_io_sinks_4_bits_last),
		.io_sinks_5_ready(_s_axi__buffered_sinkBuffer_10_io_enq_ready),
		.io_sinks_5_valid(_read_demux_io_sinks_5_valid),
		.io_sinks_5_bits_data(_read_demux_io_sinks_5_bits_data),
		.io_sinks_5_bits_resp(_read_demux_io_sinks_5_bits_resp),
		.io_sinks_5_bits_last(_read_demux_io_sinks_5_bits_last),
		.io_sinks_6_ready(_s_axi__buffered_sinkBuffer_12_io_enq_ready),
		.io_sinks_6_valid(_read_demux_io_sinks_6_valid),
		.io_sinks_6_bits_data(_read_demux_io_sinks_6_bits_data),
		.io_sinks_6_bits_resp(_read_demux_io_sinks_6_bits_resp),
		.io_sinks_6_bits_last(_read_demux_io_sinks_6_bits_last),
		.io_sinks_7_ready(_s_axi__buffered_sinkBuffer_14_io_enq_ready),
		.io_sinks_7_valid(_read_demux_io_sinks_7_valid),
		.io_sinks_7_bits_data(_read_demux_io_sinks_7_bits_data),
		.io_sinks_7_bits_resp(_read_demux_io_sinks_7_bits_resp),
		.io_sinks_7_bits_last(_read_demux_io_sinks_7_bits_last),
		.io_sinks_8_ready(_s_axi__buffered_sinkBuffer_16_io_enq_ready),
		.io_sinks_8_valid(_read_demux_io_sinks_8_valid),
		.io_sinks_8_bits_data(_read_demux_io_sinks_8_bits_data),
		.io_sinks_8_bits_resp(_read_demux_io_sinks_8_bits_resp),
		.io_sinks_8_bits_last(_read_demux_io_sinks_8_bits_last),
		.io_sinks_9_ready(_s_axi__buffered_sinkBuffer_18_io_enq_ready),
		.io_sinks_9_valid(_read_demux_io_sinks_9_valid),
		.io_sinks_9_bits_data(_read_demux_io_sinks_9_bits_data),
		.io_sinks_9_bits_resp(_read_demux_io_sinks_9_bits_resp),
		.io_sinks_9_bits_last(_read_demux_io_sinks_9_bits_last),
		.io_sinks_10_ready(_s_axi__buffered_sinkBuffer_20_io_enq_ready),
		.io_sinks_10_valid(_read_demux_io_sinks_10_valid),
		.io_sinks_10_bits_data(_read_demux_io_sinks_10_bits_data),
		.io_sinks_10_bits_resp(_read_demux_io_sinks_10_bits_resp),
		.io_sinks_10_bits_last(_read_demux_io_sinks_10_bits_last),
		.io_sinks_11_ready(_s_axi__buffered_sinkBuffer_22_io_enq_ready),
		.io_sinks_11_valid(_read_demux_io_sinks_11_valid),
		.io_sinks_11_bits_data(_read_demux_io_sinks_11_bits_data),
		.io_sinks_11_bits_resp(_read_demux_io_sinks_11_bits_resp),
		.io_sinks_11_bits_last(_read_demux_io_sinks_11_bits_last),
		.io_sinks_12_ready(_s_axi__buffered_sinkBuffer_24_io_enq_ready),
		.io_sinks_12_valid(_read_demux_io_sinks_12_valid),
		.io_sinks_12_bits_data(_read_demux_io_sinks_12_bits_data),
		.io_sinks_12_bits_resp(_read_demux_io_sinks_12_bits_resp),
		.io_sinks_12_bits_last(_read_demux_io_sinks_12_bits_last),
		.io_sinks_13_ready(_s_axi__buffered_sinkBuffer_26_io_enq_ready),
		.io_sinks_13_valid(_read_demux_io_sinks_13_valid),
		.io_sinks_13_bits_data(_read_demux_io_sinks_13_bits_data),
		.io_sinks_13_bits_resp(_read_demux_io_sinks_13_bits_resp),
		.io_sinks_13_bits_last(_read_demux_io_sinks_13_bits_last),
		.io_sinks_14_ready(_s_axi__buffered_sinkBuffer_28_io_enq_ready),
		.io_sinks_14_valid(_read_demux_io_sinks_14_valid),
		.io_sinks_14_bits_data(_read_demux_io_sinks_14_bits_data),
		.io_sinks_14_bits_resp(_read_demux_io_sinks_14_bits_resp),
		.io_sinks_14_bits_last(_read_demux_io_sinks_14_bits_last),
		.io_sinks_15_ready(_s_axi__buffered_sinkBuffer_30_io_enq_ready),
		.io_sinks_15_valid(_read_demux_io_sinks_15_valid),
		.io_sinks_15_bits_data(_read_demux_io_sinks_15_bits_data),
		.io_sinks_15_bits_resp(_read_demux_io_sinks_15_bits_resp),
		.io_sinks_15_bits_last(_read_demux_io_sinks_15_bits_last),
		.io_sinks_16_ready(_s_axi__buffered_sinkBuffer_32_io_enq_ready),
		.io_sinks_16_valid(_read_demux_io_sinks_16_valid),
		.io_sinks_16_bits_data(_read_demux_io_sinks_16_bits_data),
		.io_sinks_16_bits_resp(_read_demux_io_sinks_16_bits_resp),
		.io_sinks_16_bits_last(_read_demux_io_sinks_16_bits_last),
		.io_sinks_17_ready(_s_axi__buffered_sinkBuffer_34_io_enq_ready),
		.io_sinks_17_valid(_read_demux_io_sinks_17_valid),
		.io_sinks_17_bits_data(_read_demux_io_sinks_17_bits_data),
		.io_sinks_17_bits_resp(_read_demux_io_sinks_17_bits_resp),
		.io_sinks_17_bits_last(_read_demux_io_sinks_17_bits_last),
		.io_sinks_18_ready(_s_axi__buffered_sinkBuffer_36_io_enq_ready),
		.io_sinks_18_valid(_read_demux_io_sinks_18_valid),
		.io_sinks_18_bits_data(_read_demux_io_sinks_18_bits_data),
		.io_sinks_18_bits_resp(_read_demux_io_sinks_18_bits_resp),
		.io_sinks_18_bits_last(_read_demux_io_sinks_18_bits_last),
		.io_sinks_19_ready(_s_axi__buffered_sinkBuffer_38_io_enq_ready),
		.io_sinks_19_valid(_read_demux_io_sinks_19_valid),
		.io_sinks_19_bits_data(_read_demux_io_sinks_19_bits_data),
		.io_sinks_19_bits_resp(_read_demux_io_sinks_19_bits_resp),
		.io_sinks_19_bits_last(_read_demux_io_sinks_19_bits_last),
		.io_sinks_20_ready(_s_axi__buffered_sinkBuffer_40_io_enq_ready),
		.io_sinks_20_valid(_read_demux_io_sinks_20_valid),
		.io_sinks_20_bits_data(_read_demux_io_sinks_20_bits_data),
		.io_sinks_20_bits_resp(_read_demux_io_sinks_20_bits_resp),
		.io_sinks_20_bits_last(_read_demux_io_sinks_20_bits_last),
		.io_sinks_21_ready(_s_axi__buffered_sinkBuffer_42_io_enq_ready),
		.io_sinks_21_valid(_read_demux_io_sinks_21_valid),
		.io_sinks_21_bits_data(_read_demux_io_sinks_21_bits_data),
		.io_sinks_21_bits_resp(_read_demux_io_sinks_21_bits_resp),
		.io_sinks_21_bits_last(_read_demux_io_sinks_21_bits_last),
		.io_sinks_22_ready(_s_axi__buffered_sinkBuffer_44_io_enq_ready),
		.io_sinks_22_valid(_read_demux_io_sinks_22_valid),
		.io_sinks_22_bits_data(_read_demux_io_sinks_22_bits_data),
		.io_sinks_22_bits_resp(_read_demux_io_sinks_22_bits_resp),
		.io_sinks_22_bits_last(_read_demux_io_sinks_22_bits_last),
		.io_sinks_23_ready(_s_axi__buffered_sinkBuffer_46_io_enq_ready),
		.io_sinks_23_valid(_read_demux_io_sinks_23_valid),
		.io_sinks_23_bits_data(_read_demux_io_sinks_23_bits_data),
		.io_sinks_23_bits_resp(_read_demux_io_sinks_23_bits_resp),
		.io_sinks_23_bits_last(_read_demux_io_sinks_23_bits_last),
		.io_sinks_24_ready(_s_axi__buffered_sinkBuffer_48_io_enq_ready),
		.io_sinks_24_valid(_read_demux_io_sinks_24_valid),
		.io_sinks_24_bits_data(_read_demux_io_sinks_24_bits_data),
		.io_sinks_24_bits_resp(_read_demux_io_sinks_24_bits_resp),
		.io_sinks_24_bits_last(_read_demux_io_sinks_24_bits_last),
		.io_sinks_25_ready(_s_axi__buffered_sinkBuffer_50_io_enq_ready),
		.io_sinks_25_valid(_read_demux_io_sinks_25_valid),
		.io_sinks_25_bits_data(_read_demux_io_sinks_25_bits_data),
		.io_sinks_25_bits_resp(_read_demux_io_sinks_25_bits_resp),
		.io_sinks_25_bits_last(_read_demux_io_sinks_25_bits_last),
		.io_sinks_26_ready(_s_axi__buffered_sinkBuffer_52_io_enq_ready),
		.io_sinks_26_valid(_read_demux_io_sinks_26_valid),
		.io_sinks_26_bits_data(_read_demux_io_sinks_26_bits_data),
		.io_sinks_26_bits_resp(_read_demux_io_sinks_26_bits_resp),
		.io_sinks_26_bits_last(_read_demux_io_sinks_26_bits_last),
		.io_sinks_27_ready(_s_axi__buffered_sinkBuffer_54_io_enq_ready),
		.io_sinks_27_valid(_read_demux_io_sinks_27_valid),
		.io_sinks_27_bits_data(_read_demux_io_sinks_27_bits_data),
		.io_sinks_27_bits_resp(_read_demux_io_sinks_27_bits_resp),
		.io_sinks_27_bits_last(_read_demux_io_sinks_27_bits_last),
		.io_sinks_28_ready(_s_axi__buffered_sinkBuffer_56_io_enq_ready),
		.io_sinks_28_valid(_read_demux_io_sinks_28_valid),
		.io_sinks_28_bits_data(_read_demux_io_sinks_28_bits_data),
		.io_sinks_28_bits_resp(_read_demux_io_sinks_28_bits_resp),
		.io_sinks_28_bits_last(_read_demux_io_sinks_28_bits_last),
		.io_sinks_29_ready(_s_axi__buffered_sinkBuffer_58_io_enq_ready),
		.io_sinks_29_valid(_read_demux_io_sinks_29_valid),
		.io_sinks_29_bits_data(_read_demux_io_sinks_29_bits_data),
		.io_sinks_29_bits_resp(_read_demux_io_sinks_29_bits_resp),
		.io_sinks_29_bits_last(_read_demux_io_sinks_29_bits_last),
		.io_sinks_30_ready(_s_axi__buffered_sinkBuffer_60_io_enq_ready),
		.io_sinks_30_valid(_read_demux_io_sinks_30_valid),
		.io_sinks_30_bits_data(_read_demux_io_sinks_30_bits_data),
		.io_sinks_30_bits_resp(_read_demux_io_sinks_30_bits_resp),
		.io_sinks_30_bits_last(_read_demux_io_sinks_30_bits_last),
		.io_sinks_31_ready(_s_axi__buffered_sinkBuffer_62_io_enq_ready),
		.io_sinks_31_valid(_read_demux_io_sinks_31_valid),
		.io_sinks_31_bits_data(_read_demux_io_sinks_31_bits_data),
		.io_sinks_31_bits_resp(_read_demux_io_sinks_31_bits_resp),
		.io_sinks_31_bits_last(_read_demux_io_sinks_31_bits_last),
		.io_select_ready(_read_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_io_deq_valid & ~read_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_io_deq_bits_id)
	);
	Queue32_UInt5 write_portQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueue_io_enq_ready),
		.io_enq_valid(_write_arbiter_io_select_valid),
		.io_enq_bits(_write_arbiter_io_select_bits),
		.io_deq_ready(_write_mux_io_select_ready),
		.io_deq_valid(_write_portQueue_io_deq_valid),
		.io_deq_bits(_write_portQueue_io_deq_bits)
	);
	elasticArbiter_6 write_arbiter(
		.clock(clock),
		.reset(reset),
		.io_sources_0_ready(_write_arbiter_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_1_io_deq_valid),
		.io_sources_0_bits_addr(_s_axi__buffered_sourceBuffer_1_io_deq_bits_addr),
		.io_sources_0_bits_len(_s_axi__buffered_sourceBuffer_1_io_deq_bits_len),
		.io_sources_0_bits_size(_s_axi__buffered_sourceBuffer_1_io_deq_bits_size),
		.io_sources_0_bits_burst(_s_axi__buffered_sourceBuffer_1_io_deq_bits_burst),
		.io_sources_0_bits_lock(_s_axi__buffered_sourceBuffer_1_io_deq_bits_lock),
		.io_sources_0_bits_cache(_s_axi__buffered_sourceBuffer_1_io_deq_bits_cache),
		.io_sources_0_bits_prot(_s_axi__buffered_sourceBuffer_1_io_deq_bits_prot),
		.io_sources_0_bits_qos(_s_axi__buffered_sourceBuffer_1_io_deq_bits_qos),
		.io_sources_0_bits_region(_s_axi__buffered_sourceBuffer_1_io_deq_bits_region),
		.io_sources_1_ready(_write_arbiter_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_4_io_deq_valid),
		.io_sources_1_bits_addr(_s_axi__buffered_sourceBuffer_4_io_deq_bits_addr),
		.io_sources_1_bits_len(_s_axi__buffered_sourceBuffer_4_io_deq_bits_len),
		.io_sources_1_bits_size(_s_axi__buffered_sourceBuffer_4_io_deq_bits_size),
		.io_sources_1_bits_burst(_s_axi__buffered_sourceBuffer_4_io_deq_bits_burst),
		.io_sources_1_bits_lock(_s_axi__buffered_sourceBuffer_4_io_deq_bits_lock),
		.io_sources_1_bits_cache(_s_axi__buffered_sourceBuffer_4_io_deq_bits_cache),
		.io_sources_1_bits_prot(_s_axi__buffered_sourceBuffer_4_io_deq_bits_prot),
		.io_sources_1_bits_qos(_s_axi__buffered_sourceBuffer_4_io_deq_bits_qos),
		.io_sources_1_bits_region(_s_axi__buffered_sourceBuffer_4_io_deq_bits_region),
		.io_sources_2_ready(_write_arbiter_io_sources_2_ready),
		.io_sources_2_valid(_s_axi__buffered_sourceBuffer_7_io_deq_valid),
		.io_sources_2_bits_addr(_s_axi__buffered_sourceBuffer_7_io_deq_bits_addr),
		.io_sources_2_bits_len(_s_axi__buffered_sourceBuffer_7_io_deq_bits_len),
		.io_sources_2_bits_size(_s_axi__buffered_sourceBuffer_7_io_deq_bits_size),
		.io_sources_2_bits_burst(_s_axi__buffered_sourceBuffer_7_io_deq_bits_burst),
		.io_sources_2_bits_lock(_s_axi__buffered_sourceBuffer_7_io_deq_bits_lock),
		.io_sources_2_bits_cache(_s_axi__buffered_sourceBuffer_7_io_deq_bits_cache),
		.io_sources_2_bits_prot(_s_axi__buffered_sourceBuffer_7_io_deq_bits_prot),
		.io_sources_2_bits_qos(_s_axi__buffered_sourceBuffer_7_io_deq_bits_qos),
		.io_sources_2_bits_region(_s_axi__buffered_sourceBuffer_7_io_deq_bits_region),
		.io_sources_3_ready(_write_arbiter_io_sources_3_ready),
		.io_sources_3_valid(_s_axi__buffered_sourceBuffer_10_io_deq_valid),
		.io_sources_3_bits_addr(_s_axi__buffered_sourceBuffer_10_io_deq_bits_addr),
		.io_sources_3_bits_len(_s_axi__buffered_sourceBuffer_10_io_deq_bits_len),
		.io_sources_3_bits_size(_s_axi__buffered_sourceBuffer_10_io_deq_bits_size),
		.io_sources_3_bits_burst(_s_axi__buffered_sourceBuffer_10_io_deq_bits_burst),
		.io_sources_3_bits_lock(_s_axi__buffered_sourceBuffer_10_io_deq_bits_lock),
		.io_sources_3_bits_cache(_s_axi__buffered_sourceBuffer_10_io_deq_bits_cache),
		.io_sources_3_bits_prot(_s_axi__buffered_sourceBuffer_10_io_deq_bits_prot),
		.io_sources_3_bits_qos(_s_axi__buffered_sourceBuffer_10_io_deq_bits_qos),
		.io_sources_3_bits_region(_s_axi__buffered_sourceBuffer_10_io_deq_bits_region),
		.io_sources_4_ready(_write_arbiter_io_sources_4_ready),
		.io_sources_4_valid(_s_axi__buffered_sourceBuffer_13_io_deq_valid),
		.io_sources_4_bits_addr(_s_axi__buffered_sourceBuffer_13_io_deq_bits_addr),
		.io_sources_4_bits_len(_s_axi__buffered_sourceBuffer_13_io_deq_bits_len),
		.io_sources_4_bits_size(_s_axi__buffered_sourceBuffer_13_io_deq_bits_size),
		.io_sources_4_bits_burst(_s_axi__buffered_sourceBuffer_13_io_deq_bits_burst),
		.io_sources_4_bits_lock(_s_axi__buffered_sourceBuffer_13_io_deq_bits_lock),
		.io_sources_4_bits_cache(_s_axi__buffered_sourceBuffer_13_io_deq_bits_cache),
		.io_sources_4_bits_prot(_s_axi__buffered_sourceBuffer_13_io_deq_bits_prot),
		.io_sources_4_bits_qos(_s_axi__buffered_sourceBuffer_13_io_deq_bits_qos),
		.io_sources_4_bits_region(_s_axi__buffered_sourceBuffer_13_io_deq_bits_region),
		.io_sources_5_ready(_write_arbiter_io_sources_5_ready),
		.io_sources_5_valid(_s_axi__buffered_sourceBuffer_16_io_deq_valid),
		.io_sources_5_bits_addr(_s_axi__buffered_sourceBuffer_16_io_deq_bits_addr),
		.io_sources_5_bits_len(_s_axi__buffered_sourceBuffer_16_io_deq_bits_len),
		.io_sources_5_bits_size(_s_axi__buffered_sourceBuffer_16_io_deq_bits_size),
		.io_sources_5_bits_burst(_s_axi__buffered_sourceBuffer_16_io_deq_bits_burst),
		.io_sources_5_bits_lock(_s_axi__buffered_sourceBuffer_16_io_deq_bits_lock),
		.io_sources_5_bits_cache(_s_axi__buffered_sourceBuffer_16_io_deq_bits_cache),
		.io_sources_5_bits_prot(_s_axi__buffered_sourceBuffer_16_io_deq_bits_prot),
		.io_sources_5_bits_qos(_s_axi__buffered_sourceBuffer_16_io_deq_bits_qos),
		.io_sources_5_bits_region(_s_axi__buffered_sourceBuffer_16_io_deq_bits_region),
		.io_sources_6_ready(_write_arbiter_io_sources_6_ready),
		.io_sources_6_valid(_s_axi__buffered_sourceBuffer_19_io_deq_valid),
		.io_sources_6_bits_addr(_s_axi__buffered_sourceBuffer_19_io_deq_bits_addr),
		.io_sources_6_bits_len(_s_axi__buffered_sourceBuffer_19_io_deq_bits_len),
		.io_sources_6_bits_size(_s_axi__buffered_sourceBuffer_19_io_deq_bits_size),
		.io_sources_6_bits_burst(_s_axi__buffered_sourceBuffer_19_io_deq_bits_burst),
		.io_sources_6_bits_lock(_s_axi__buffered_sourceBuffer_19_io_deq_bits_lock),
		.io_sources_6_bits_cache(_s_axi__buffered_sourceBuffer_19_io_deq_bits_cache),
		.io_sources_6_bits_prot(_s_axi__buffered_sourceBuffer_19_io_deq_bits_prot),
		.io_sources_6_bits_qos(_s_axi__buffered_sourceBuffer_19_io_deq_bits_qos),
		.io_sources_6_bits_region(_s_axi__buffered_sourceBuffer_19_io_deq_bits_region),
		.io_sources_7_ready(_write_arbiter_io_sources_7_ready),
		.io_sources_7_valid(_s_axi__buffered_sourceBuffer_22_io_deq_valid),
		.io_sources_7_bits_addr(_s_axi__buffered_sourceBuffer_22_io_deq_bits_addr),
		.io_sources_7_bits_len(_s_axi__buffered_sourceBuffer_22_io_deq_bits_len),
		.io_sources_7_bits_size(_s_axi__buffered_sourceBuffer_22_io_deq_bits_size),
		.io_sources_7_bits_burst(_s_axi__buffered_sourceBuffer_22_io_deq_bits_burst),
		.io_sources_7_bits_lock(_s_axi__buffered_sourceBuffer_22_io_deq_bits_lock),
		.io_sources_7_bits_cache(_s_axi__buffered_sourceBuffer_22_io_deq_bits_cache),
		.io_sources_7_bits_prot(_s_axi__buffered_sourceBuffer_22_io_deq_bits_prot),
		.io_sources_7_bits_qos(_s_axi__buffered_sourceBuffer_22_io_deq_bits_qos),
		.io_sources_7_bits_region(_s_axi__buffered_sourceBuffer_22_io_deq_bits_region),
		.io_sources_8_ready(_write_arbiter_io_sources_8_ready),
		.io_sources_8_valid(_s_axi__buffered_sourceBuffer_25_io_deq_valid),
		.io_sources_8_bits_addr(_s_axi__buffered_sourceBuffer_25_io_deq_bits_addr),
		.io_sources_8_bits_len(_s_axi__buffered_sourceBuffer_25_io_deq_bits_len),
		.io_sources_8_bits_size(_s_axi__buffered_sourceBuffer_25_io_deq_bits_size),
		.io_sources_8_bits_burst(_s_axi__buffered_sourceBuffer_25_io_deq_bits_burst),
		.io_sources_8_bits_lock(_s_axi__buffered_sourceBuffer_25_io_deq_bits_lock),
		.io_sources_8_bits_cache(_s_axi__buffered_sourceBuffer_25_io_deq_bits_cache),
		.io_sources_8_bits_prot(_s_axi__buffered_sourceBuffer_25_io_deq_bits_prot),
		.io_sources_8_bits_qos(_s_axi__buffered_sourceBuffer_25_io_deq_bits_qos),
		.io_sources_8_bits_region(_s_axi__buffered_sourceBuffer_25_io_deq_bits_region),
		.io_sources_9_ready(_write_arbiter_io_sources_9_ready),
		.io_sources_9_valid(_s_axi__buffered_sourceBuffer_28_io_deq_valid),
		.io_sources_9_bits_addr(_s_axi__buffered_sourceBuffer_28_io_deq_bits_addr),
		.io_sources_9_bits_len(_s_axi__buffered_sourceBuffer_28_io_deq_bits_len),
		.io_sources_9_bits_size(_s_axi__buffered_sourceBuffer_28_io_deq_bits_size),
		.io_sources_9_bits_burst(_s_axi__buffered_sourceBuffer_28_io_deq_bits_burst),
		.io_sources_9_bits_lock(_s_axi__buffered_sourceBuffer_28_io_deq_bits_lock),
		.io_sources_9_bits_cache(_s_axi__buffered_sourceBuffer_28_io_deq_bits_cache),
		.io_sources_9_bits_prot(_s_axi__buffered_sourceBuffer_28_io_deq_bits_prot),
		.io_sources_9_bits_qos(_s_axi__buffered_sourceBuffer_28_io_deq_bits_qos),
		.io_sources_9_bits_region(_s_axi__buffered_sourceBuffer_28_io_deq_bits_region),
		.io_sources_10_ready(_write_arbiter_io_sources_10_ready),
		.io_sources_10_valid(_s_axi__buffered_sourceBuffer_31_io_deq_valid),
		.io_sources_10_bits_addr(_s_axi__buffered_sourceBuffer_31_io_deq_bits_addr),
		.io_sources_10_bits_len(_s_axi__buffered_sourceBuffer_31_io_deq_bits_len),
		.io_sources_10_bits_size(_s_axi__buffered_sourceBuffer_31_io_deq_bits_size),
		.io_sources_10_bits_burst(_s_axi__buffered_sourceBuffer_31_io_deq_bits_burst),
		.io_sources_10_bits_lock(_s_axi__buffered_sourceBuffer_31_io_deq_bits_lock),
		.io_sources_10_bits_cache(_s_axi__buffered_sourceBuffer_31_io_deq_bits_cache),
		.io_sources_10_bits_prot(_s_axi__buffered_sourceBuffer_31_io_deq_bits_prot),
		.io_sources_10_bits_qos(_s_axi__buffered_sourceBuffer_31_io_deq_bits_qos),
		.io_sources_10_bits_region(_s_axi__buffered_sourceBuffer_31_io_deq_bits_region),
		.io_sources_11_ready(_write_arbiter_io_sources_11_ready),
		.io_sources_11_valid(_s_axi__buffered_sourceBuffer_34_io_deq_valid),
		.io_sources_11_bits_addr(_s_axi__buffered_sourceBuffer_34_io_deq_bits_addr),
		.io_sources_11_bits_len(_s_axi__buffered_sourceBuffer_34_io_deq_bits_len),
		.io_sources_11_bits_size(_s_axi__buffered_sourceBuffer_34_io_deq_bits_size),
		.io_sources_11_bits_burst(_s_axi__buffered_sourceBuffer_34_io_deq_bits_burst),
		.io_sources_11_bits_lock(_s_axi__buffered_sourceBuffer_34_io_deq_bits_lock),
		.io_sources_11_bits_cache(_s_axi__buffered_sourceBuffer_34_io_deq_bits_cache),
		.io_sources_11_bits_prot(_s_axi__buffered_sourceBuffer_34_io_deq_bits_prot),
		.io_sources_11_bits_qos(_s_axi__buffered_sourceBuffer_34_io_deq_bits_qos),
		.io_sources_11_bits_region(_s_axi__buffered_sourceBuffer_34_io_deq_bits_region),
		.io_sources_12_ready(_write_arbiter_io_sources_12_ready),
		.io_sources_12_valid(_s_axi__buffered_sourceBuffer_37_io_deq_valid),
		.io_sources_12_bits_addr(_s_axi__buffered_sourceBuffer_37_io_deq_bits_addr),
		.io_sources_12_bits_len(_s_axi__buffered_sourceBuffer_37_io_deq_bits_len),
		.io_sources_12_bits_size(_s_axi__buffered_sourceBuffer_37_io_deq_bits_size),
		.io_sources_12_bits_burst(_s_axi__buffered_sourceBuffer_37_io_deq_bits_burst),
		.io_sources_12_bits_lock(_s_axi__buffered_sourceBuffer_37_io_deq_bits_lock),
		.io_sources_12_bits_cache(_s_axi__buffered_sourceBuffer_37_io_deq_bits_cache),
		.io_sources_12_bits_prot(_s_axi__buffered_sourceBuffer_37_io_deq_bits_prot),
		.io_sources_12_bits_qos(_s_axi__buffered_sourceBuffer_37_io_deq_bits_qos),
		.io_sources_12_bits_region(_s_axi__buffered_sourceBuffer_37_io_deq_bits_region),
		.io_sources_13_ready(_write_arbiter_io_sources_13_ready),
		.io_sources_13_valid(_s_axi__buffered_sourceBuffer_40_io_deq_valid),
		.io_sources_13_bits_addr(_s_axi__buffered_sourceBuffer_40_io_deq_bits_addr),
		.io_sources_13_bits_len(_s_axi__buffered_sourceBuffer_40_io_deq_bits_len),
		.io_sources_13_bits_size(_s_axi__buffered_sourceBuffer_40_io_deq_bits_size),
		.io_sources_13_bits_burst(_s_axi__buffered_sourceBuffer_40_io_deq_bits_burst),
		.io_sources_13_bits_lock(_s_axi__buffered_sourceBuffer_40_io_deq_bits_lock),
		.io_sources_13_bits_cache(_s_axi__buffered_sourceBuffer_40_io_deq_bits_cache),
		.io_sources_13_bits_prot(_s_axi__buffered_sourceBuffer_40_io_deq_bits_prot),
		.io_sources_13_bits_qos(_s_axi__buffered_sourceBuffer_40_io_deq_bits_qos),
		.io_sources_13_bits_region(_s_axi__buffered_sourceBuffer_40_io_deq_bits_region),
		.io_sources_14_ready(_write_arbiter_io_sources_14_ready),
		.io_sources_14_valid(_s_axi__buffered_sourceBuffer_43_io_deq_valid),
		.io_sources_14_bits_addr(_s_axi__buffered_sourceBuffer_43_io_deq_bits_addr),
		.io_sources_14_bits_len(_s_axi__buffered_sourceBuffer_43_io_deq_bits_len),
		.io_sources_14_bits_size(_s_axi__buffered_sourceBuffer_43_io_deq_bits_size),
		.io_sources_14_bits_burst(_s_axi__buffered_sourceBuffer_43_io_deq_bits_burst),
		.io_sources_14_bits_lock(_s_axi__buffered_sourceBuffer_43_io_deq_bits_lock),
		.io_sources_14_bits_cache(_s_axi__buffered_sourceBuffer_43_io_deq_bits_cache),
		.io_sources_14_bits_prot(_s_axi__buffered_sourceBuffer_43_io_deq_bits_prot),
		.io_sources_14_bits_qos(_s_axi__buffered_sourceBuffer_43_io_deq_bits_qos),
		.io_sources_14_bits_region(_s_axi__buffered_sourceBuffer_43_io_deq_bits_region),
		.io_sources_15_ready(_write_arbiter_io_sources_15_ready),
		.io_sources_15_valid(_s_axi__buffered_sourceBuffer_46_io_deq_valid),
		.io_sources_15_bits_addr(_s_axi__buffered_sourceBuffer_46_io_deq_bits_addr),
		.io_sources_15_bits_len(_s_axi__buffered_sourceBuffer_46_io_deq_bits_len),
		.io_sources_15_bits_size(_s_axi__buffered_sourceBuffer_46_io_deq_bits_size),
		.io_sources_15_bits_burst(_s_axi__buffered_sourceBuffer_46_io_deq_bits_burst),
		.io_sources_15_bits_lock(_s_axi__buffered_sourceBuffer_46_io_deq_bits_lock),
		.io_sources_15_bits_cache(_s_axi__buffered_sourceBuffer_46_io_deq_bits_cache),
		.io_sources_15_bits_prot(_s_axi__buffered_sourceBuffer_46_io_deq_bits_prot),
		.io_sources_15_bits_qos(_s_axi__buffered_sourceBuffer_46_io_deq_bits_qos),
		.io_sources_15_bits_region(_s_axi__buffered_sourceBuffer_46_io_deq_bits_region),
		.io_sources_16_ready(_write_arbiter_io_sources_16_ready),
		.io_sources_16_valid(_s_axi__buffered_sourceBuffer_49_io_deq_valid),
		.io_sources_16_bits_addr(_s_axi__buffered_sourceBuffer_49_io_deq_bits_addr),
		.io_sources_16_bits_len(_s_axi__buffered_sourceBuffer_49_io_deq_bits_len),
		.io_sources_16_bits_size(_s_axi__buffered_sourceBuffer_49_io_deq_bits_size),
		.io_sources_16_bits_burst(_s_axi__buffered_sourceBuffer_49_io_deq_bits_burst),
		.io_sources_16_bits_lock(_s_axi__buffered_sourceBuffer_49_io_deq_bits_lock),
		.io_sources_16_bits_cache(_s_axi__buffered_sourceBuffer_49_io_deq_bits_cache),
		.io_sources_16_bits_prot(_s_axi__buffered_sourceBuffer_49_io_deq_bits_prot),
		.io_sources_16_bits_qos(_s_axi__buffered_sourceBuffer_49_io_deq_bits_qos),
		.io_sources_16_bits_region(_s_axi__buffered_sourceBuffer_49_io_deq_bits_region),
		.io_sources_17_ready(_write_arbiter_io_sources_17_ready),
		.io_sources_17_valid(_s_axi__buffered_sourceBuffer_52_io_deq_valid),
		.io_sources_17_bits_addr(_s_axi__buffered_sourceBuffer_52_io_deq_bits_addr),
		.io_sources_17_bits_len(_s_axi__buffered_sourceBuffer_52_io_deq_bits_len),
		.io_sources_17_bits_size(_s_axi__buffered_sourceBuffer_52_io_deq_bits_size),
		.io_sources_17_bits_burst(_s_axi__buffered_sourceBuffer_52_io_deq_bits_burst),
		.io_sources_17_bits_lock(_s_axi__buffered_sourceBuffer_52_io_deq_bits_lock),
		.io_sources_17_bits_cache(_s_axi__buffered_sourceBuffer_52_io_deq_bits_cache),
		.io_sources_17_bits_prot(_s_axi__buffered_sourceBuffer_52_io_deq_bits_prot),
		.io_sources_17_bits_qos(_s_axi__buffered_sourceBuffer_52_io_deq_bits_qos),
		.io_sources_17_bits_region(_s_axi__buffered_sourceBuffer_52_io_deq_bits_region),
		.io_sources_18_ready(_write_arbiter_io_sources_18_ready),
		.io_sources_18_valid(_s_axi__buffered_sourceBuffer_55_io_deq_valid),
		.io_sources_18_bits_addr(_s_axi__buffered_sourceBuffer_55_io_deq_bits_addr),
		.io_sources_18_bits_len(_s_axi__buffered_sourceBuffer_55_io_deq_bits_len),
		.io_sources_18_bits_size(_s_axi__buffered_sourceBuffer_55_io_deq_bits_size),
		.io_sources_18_bits_burst(_s_axi__buffered_sourceBuffer_55_io_deq_bits_burst),
		.io_sources_18_bits_lock(_s_axi__buffered_sourceBuffer_55_io_deq_bits_lock),
		.io_sources_18_bits_cache(_s_axi__buffered_sourceBuffer_55_io_deq_bits_cache),
		.io_sources_18_bits_prot(_s_axi__buffered_sourceBuffer_55_io_deq_bits_prot),
		.io_sources_18_bits_qos(_s_axi__buffered_sourceBuffer_55_io_deq_bits_qos),
		.io_sources_18_bits_region(_s_axi__buffered_sourceBuffer_55_io_deq_bits_region),
		.io_sources_19_ready(_write_arbiter_io_sources_19_ready),
		.io_sources_19_valid(_s_axi__buffered_sourceBuffer_58_io_deq_valid),
		.io_sources_19_bits_addr(_s_axi__buffered_sourceBuffer_58_io_deq_bits_addr),
		.io_sources_19_bits_len(_s_axi__buffered_sourceBuffer_58_io_deq_bits_len),
		.io_sources_19_bits_size(_s_axi__buffered_sourceBuffer_58_io_deq_bits_size),
		.io_sources_19_bits_burst(_s_axi__buffered_sourceBuffer_58_io_deq_bits_burst),
		.io_sources_19_bits_lock(_s_axi__buffered_sourceBuffer_58_io_deq_bits_lock),
		.io_sources_19_bits_cache(_s_axi__buffered_sourceBuffer_58_io_deq_bits_cache),
		.io_sources_19_bits_prot(_s_axi__buffered_sourceBuffer_58_io_deq_bits_prot),
		.io_sources_19_bits_qos(_s_axi__buffered_sourceBuffer_58_io_deq_bits_qos),
		.io_sources_19_bits_region(_s_axi__buffered_sourceBuffer_58_io_deq_bits_region),
		.io_sources_20_ready(_write_arbiter_io_sources_20_ready),
		.io_sources_20_valid(_s_axi__buffered_sourceBuffer_61_io_deq_valid),
		.io_sources_20_bits_addr(_s_axi__buffered_sourceBuffer_61_io_deq_bits_addr),
		.io_sources_20_bits_len(_s_axi__buffered_sourceBuffer_61_io_deq_bits_len),
		.io_sources_20_bits_size(_s_axi__buffered_sourceBuffer_61_io_deq_bits_size),
		.io_sources_20_bits_burst(_s_axi__buffered_sourceBuffer_61_io_deq_bits_burst),
		.io_sources_20_bits_lock(_s_axi__buffered_sourceBuffer_61_io_deq_bits_lock),
		.io_sources_20_bits_cache(_s_axi__buffered_sourceBuffer_61_io_deq_bits_cache),
		.io_sources_20_bits_prot(_s_axi__buffered_sourceBuffer_61_io_deq_bits_prot),
		.io_sources_20_bits_qos(_s_axi__buffered_sourceBuffer_61_io_deq_bits_qos),
		.io_sources_20_bits_region(_s_axi__buffered_sourceBuffer_61_io_deq_bits_region),
		.io_sources_21_ready(_write_arbiter_io_sources_21_ready),
		.io_sources_21_valid(_s_axi__buffered_sourceBuffer_64_io_deq_valid),
		.io_sources_21_bits_addr(_s_axi__buffered_sourceBuffer_64_io_deq_bits_addr),
		.io_sources_21_bits_len(_s_axi__buffered_sourceBuffer_64_io_deq_bits_len),
		.io_sources_21_bits_size(_s_axi__buffered_sourceBuffer_64_io_deq_bits_size),
		.io_sources_21_bits_burst(_s_axi__buffered_sourceBuffer_64_io_deq_bits_burst),
		.io_sources_21_bits_lock(_s_axi__buffered_sourceBuffer_64_io_deq_bits_lock),
		.io_sources_21_bits_cache(_s_axi__buffered_sourceBuffer_64_io_deq_bits_cache),
		.io_sources_21_bits_prot(_s_axi__buffered_sourceBuffer_64_io_deq_bits_prot),
		.io_sources_21_bits_qos(_s_axi__buffered_sourceBuffer_64_io_deq_bits_qos),
		.io_sources_21_bits_region(_s_axi__buffered_sourceBuffer_64_io_deq_bits_region),
		.io_sources_22_ready(_write_arbiter_io_sources_22_ready),
		.io_sources_22_valid(_s_axi__buffered_sourceBuffer_67_io_deq_valid),
		.io_sources_22_bits_addr(_s_axi__buffered_sourceBuffer_67_io_deq_bits_addr),
		.io_sources_22_bits_len(_s_axi__buffered_sourceBuffer_67_io_deq_bits_len),
		.io_sources_22_bits_size(_s_axi__buffered_sourceBuffer_67_io_deq_bits_size),
		.io_sources_22_bits_burst(_s_axi__buffered_sourceBuffer_67_io_deq_bits_burst),
		.io_sources_22_bits_lock(_s_axi__buffered_sourceBuffer_67_io_deq_bits_lock),
		.io_sources_22_bits_cache(_s_axi__buffered_sourceBuffer_67_io_deq_bits_cache),
		.io_sources_22_bits_prot(_s_axi__buffered_sourceBuffer_67_io_deq_bits_prot),
		.io_sources_22_bits_qos(_s_axi__buffered_sourceBuffer_67_io_deq_bits_qos),
		.io_sources_22_bits_region(_s_axi__buffered_sourceBuffer_67_io_deq_bits_region),
		.io_sources_23_ready(_write_arbiter_io_sources_23_ready),
		.io_sources_23_valid(_s_axi__buffered_sourceBuffer_70_io_deq_valid),
		.io_sources_23_bits_addr(_s_axi__buffered_sourceBuffer_70_io_deq_bits_addr),
		.io_sources_23_bits_len(_s_axi__buffered_sourceBuffer_70_io_deq_bits_len),
		.io_sources_23_bits_size(_s_axi__buffered_sourceBuffer_70_io_deq_bits_size),
		.io_sources_23_bits_burst(_s_axi__buffered_sourceBuffer_70_io_deq_bits_burst),
		.io_sources_23_bits_lock(_s_axi__buffered_sourceBuffer_70_io_deq_bits_lock),
		.io_sources_23_bits_cache(_s_axi__buffered_sourceBuffer_70_io_deq_bits_cache),
		.io_sources_23_bits_prot(_s_axi__buffered_sourceBuffer_70_io_deq_bits_prot),
		.io_sources_23_bits_qos(_s_axi__buffered_sourceBuffer_70_io_deq_bits_qos),
		.io_sources_23_bits_region(_s_axi__buffered_sourceBuffer_70_io_deq_bits_region),
		.io_sources_24_ready(_write_arbiter_io_sources_24_ready),
		.io_sources_24_valid(_s_axi__buffered_sourceBuffer_73_io_deq_valid),
		.io_sources_24_bits_addr(_s_axi__buffered_sourceBuffer_73_io_deq_bits_addr),
		.io_sources_24_bits_len(_s_axi__buffered_sourceBuffer_73_io_deq_bits_len),
		.io_sources_24_bits_size(_s_axi__buffered_sourceBuffer_73_io_deq_bits_size),
		.io_sources_24_bits_burst(_s_axi__buffered_sourceBuffer_73_io_deq_bits_burst),
		.io_sources_24_bits_lock(_s_axi__buffered_sourceBuffer_73_io_deq_bits_lock),
		.io_sources_24_bits_cache(_s_axi__buffered_sourceBuffer_73_io_deq_bits_cache),
		.io_sources_24_bits_prot(_s_axi__buffered_sourceBuffer_73_io_deq_bits_prot),
		.io_sources_24_bits_qos(_s_axi__buffered_sourceBuffer_73_io_deq_bits_qos),
		.io_sources_24_bits_region(_s_axi__buffered_sourceBuffer_73_io_deq_bits_region),
		.io_sources_25_ready(_write_arbiter_io_sources_25_ready),
		.io_sources_25_valid(_s_axi__buffered_sourceBuffer_76_io_deq_valid),
		.io_sources_25_bits_addr(_s_axi__buffered_sourceBuffer_76_io_deq_bits_addr),
		.io_sources_25_bits_len(_s_axi__buffered_sourceBuffer_76_io_deq_bits_len),
		.io_sources_25_bits_size(_s_axi__buffered_sourceBuffer_76_io_deq_bits_size),
		.io_sources_25_bits_burst(_s_axi__buffered_sourceBuffer_76_io_deq_bits_burst),
		.io_sources_25_bits_lock(_s_axi__buffered_sourceBuffer_76_io_deq_bits_lock),
		.io_sources_25_bits_cache(_s_axi__buffered_sourceBuffer_76_io_deq_bits_cache),
		.io_sources_25_bits_prot(_s_axi__buffered_sourceBuffer_76_io_deq_bits_prot),
		.io_sources_25_bits_qos(_s_axi__buffered_sourceBuffer_76_io_deq_bits_qos),
		.io_sources_25_bits_region(_s_axi__buffered_sourceBuffer_76_io_deq_bits_region),
		.io_sources_26_ready(_write_arbiter_io_sources_26_ready),
		.io_sources_26_valid(_s_axi__buffered_sourceBuffer_79_io_deq_valid),
		.io_sources_26_bits_addr(_s_axi__buffered_sourceBuffer_79_io_deq_bits_addr),
		.io_sources_26_bits_len(_s_axi__buffered_sourceBuffer_79_io_deq_bits_len),
		.io_sources_26_bits_size(_s_axi__buffered_sourceBuffer_79_io_deq_bits_size),
		.io_sources_26_bits_burst(_s_axi__buffered_sourceBuffer_79_io_deq_bits_burst),
		.io_sources_26_bits_lock(_s_axi__buffered_sourceBuffer_79_io_deq_bits_lock),
		.io_sources_26_bits_cache(_s_axi__buffered_sourceBuffer_79_io_deq_bits_cache),
		.io_sources_26_bits_prot(_s_axi__buffered_sourceBuffer_79_io_deq_bits_prot),
		.io_sources_26_bits_qos(_s_axi__buffered_sourceBuffer_79_io_deq_bits_qos),
		.io_sources_26_bits_region(_s_axi__buffered_sourceBuffer_79_io_deq_bits_region),
		.io_sources_27_ready(_write_arbiter_io_sources_27_ready),
		.io_sources_27_valid(_s_axi__buffered_sourceBuffer_82_io_deq_valid),
		.io_sources_27_bits_addr(_s_axi__buffered_sourceBuffer_82_io_deq_bits_addr),
		.io_sources_27_bits_len(_s_axi__buffered_sourceBuffer_82_io_deq_bits_len),
		.io_sources_27_bits_size(_s_axi__buffered_sourceBuffer_82_io_deq_bits_size),
		.io_sources_27_bits_burst(_s_axi__buffered_sourceBuffer_82_io_deq_bits_burst),
		.io_sources_27_bits_lock(_s_axi__buffered_sourceBuffer_82_io_deq_bits_lock),
		.io_sources_27_bits_cache(_s_axi__buffered_sourceBuffer_82_io_deq_bits_cache),
		.io_sources_27_bits_prot(_s_axi__buffered_sourceBuffer_82_io_deq_bits_prot),
		.io_sources_27_bits_qos(_s_axi__buffered_sourceBuffer_82_io_deq_bits_qos),
		.io_sources_27_bits_region(_s_axi__buffered_sourceBuffer_82_io_deq_bits_region),
		.io_sources_28_ready(_write_arbiter_io_sources_28_ready),
		.io_sources_28_valid(_s_axi__buffered_sourceBuffer_85_io_deq_valid),
		.io_sources_28_bits_addr(_s_axi__buffered_sourceBuffer_85_io_deq_bits_addr),
		.io_sources_28_bits_len(_s_axi__buffered_sourceBuffer_85_io_deq_bits_len),
		.io_sources_28_bits_size(_s_axi__buffered_sourceBuffer_85_io_deq_bits_size),
		.io_sources_28_bits_burst(_s_axi__buffered_sourceBuffer_85_io_deq_bits_burst),
		.io_sources_28_bits_lock(_s_axi__buffered_sourceBuffer_85_io_deq_bits_lock),
		.io_sources_28_bits_cache(_s_axi__buffered_sourceBuffer_85_io_deq_bits_cache),
		.io_sources_28_bits_prot(_s_axi__buffered_sourceBuffer_85_io_deq_bits_prot),
		.io_sources_28_bits_qos(_s_axi__buffered_sourceBuffer_85_io_deq_bits_qos),
		.io_sources_28_bits_region(_s_axi__buffered_sourceBuffer_85_io_deq_bits_region),
		.io_sources_29_ready(_write_arbiter_io_sources_29_ready),
		.io_sources_29_valid(_s_axi__buffered_sourceBuffer_88_io_deq_valid),
		.io_sources_29_bits_addr(_s_axi__buffered_sourceBuffer_88_io_deq_bits_addr),
		.io_sources_29_bits_len(_s_axi__buffered_sourceBuffer_88_io_deq_bits_len),
		.io_sources_29_bits_size(_s_axi__buffered_sourceBuffer_88_io_deq_bits_size),
		.io_sources_29_bits_burst(_s_axi__buffered_sourceBuffer_88_io_deq_bits_burst),
		.io_sources_29_bits_lock(_s_axi__buffered_sourceBuffer_88_io_deq_bits_lock),
		.io_sources_29_bits_cache(_s_axi__buffered_sourceBuffer_88_io_deq_bits_cache),
		.io_sources_29_bits_prot(_s_axi__buffered_sourceBuffer_88_io_deq_bits_prot),
		.io_sources_29_bits_qos(_s_axi__buffered_sourceBuffer_88_io_deq_bits_qos),
		.io_sources_29_bits_region(_s_axi__buffered_sourceBuffer_88_io_deq_bits_region),
		.io_sources_30_ready(_write_arbiter_io_sources_30_ready),
		.io_sources_30_valid(_s_axi__buffered_sourceBuffer_91_io_deq_valid),
		.io_sources_30_bits_addr(_s_axi__buffered_sourceBuffer_91_io_deq_bits_addr),
		.io_sources_30_bits_len(_s_axi__buffered_sourceBuffer_91_io_deq_bits_len),
		.io_sources_30_bits_size(_s_axi__buffered_sourceBuffer_91_io_deq_bits_size),
		.io_sources_30_bits_burst(_s_axi__buffered_sourceBuffer_91_io_deq_bits_burst),
		.io_sources_30_bits_lock(_s_axi__buffered_sourceBuffer_91_io_deq_bits_lock),
		.io_sources_30_bits_cache(_s_axi__buffered_sourceBuffer_91_io_deq_bits_cache),
		.io_sources_30_bits_prot(_s_axi__buffered_sourceBuffer_91_io_deq_bits_prot),
		.io_sources_30_bits_qos(_s_axi__buffered_sourceBuffer_91_io_deq_bits_qos),
		.io_sources_30_bits_region(_s_axi__buffered_sourceBuffer_91_io_deq_bits_region),
		.io_sources_31_ready(_write_arbiter_io_sources_31_ready),
		.io_sources_31_valid(_s_axi__buffered_sourceBuffer_94_io_deq_valid),
		.io_sources_31_bits_addr(_s_axi__buffered_sourceBuffer_94_io_deq_bits_addr),
		.io_sources_31_bits_len(_s_axi__buffered_sourceBuffer_94_io_deq_bits_len),
		.io_sources_31_bits_size(_s_axi__buffered_sourceBuffer_94_io_deq_bits_size),
		.io_sources_31_bits_burst(_s_axi__buffered_sourceBuffer_94_io_deq_bits_burst),
		.io_sources_31_bits_lock(_s_axi__buffered_sourceBuffer_94_io_deq_bits_lock),
		.io_sources_31_bits_cache(_s_axi__buffered_sourceBuffer_94_io_deq_bits_cache),
		.io_sources_31_bits_prot(_s_axi__buffered_sourceBuffer_94_io_deq_bits_prot),
		.io_sources_31_bits_qos(_s_axi__buffered_sourceBuffer_94_io_deq_bits_qos),
		.io_sources_31_bits_region(_s_axi__buffered_sourceBuffer_94_io_deq_bits_region),
		.io_sink_ready(_m_axi__sourceBuffer_1_io_enq_ready),
		.io_sink_valid(_write_arbiter_io_sink_valid),
		.io_sink_bits_id(_write_arbiter_io_sink_bits_id),
		.io_sink_bits_addr(_write_arbiter_io_sink_bits_addr),
		.io_sink_bits_len(_write_arbiter_io_sink_bits_len),
		.io_sink_bits_size(_write_arbiter_io_sink_bits_size),
		.io_sink_bits_burst(_write_arbiter_io_sink_bits_burst),
		.io_sink_bits_lock(_write_arbiter_io_sink_bits_lock),
		.io_sink_bits_cache(_write_arbiter_io_sink_bits_cache),
		.io_sink_bits_prot(_write_arbiter_io_sink_bits_prot),
		.io_sink_bits_qos(_write_arbiter_io_sink_bits_qos),
		.io_sink_bits_region(_write_arbiter_io_sink_bits_region),
		.io_select_ready(_write_portQueue_io_enq_ready),
		.io_select_valid(_write_arbiter_io_select_valid),
		.io_select_bits(_write_arbiter_io_select_bits)
	);
	elasticMux_5 write_mux(
		.io_sources_0_ready(_write_mux_io_sources_0_ready),
		.io_sources_0_valid(_s_axi__buffered_sourceBuffer_2_io_deq_valid),
		.io_sources_0_bits_data(_s_axi__buffered_sourceBuffer_2_io_deq_bits_data),
		.io_sources_0_bits_strb(_s_axi__buffered_sourceBuffer_2_io_deq_bits_strb),
		.io_sources_0_bits_last(_s_axi__buffered_sourceBuffer_2_io_deq_bits_last),
		.io_sources_1_ready(_write_mux_io_sources_1_ready),
		.io_sources_1_valid(_s_axi__buffered_sourceBuffer_5_io_deq_valid),
		.io_sources_1_bits_data(_s_axi__buffered_sourceBuffer_5_io_deq_bits_data),
		.io_sources_1_bits_strb(_s_axi__buffered_sourceBuffer_5_io_deq_bits_strb),
		.io_sources_1_bits_last(_s_axi__buffered_sourceBuffer_5_io_deq_bits_last),
		.io_sources_2_ready(_write_mux_io_sources_2_ready),
		.io_sources_2_valid(_s_axi__buffered_sourceBuffer_8_io_deq_valid),
		.io_sources_2_bits_data(_s_axi__buffered_sourceBuffer_8_io_deq_bits_data),
		.io_sources_2_bits_strb(_s_axi__buffered_sourceBuffer_8_io_deq_bits_strb),
		.io_sources_2_bits_last(_s_axi__buffered_sourceBuffer_8_io_deq_bits_last),
		.io_sources_3_ready(_write_mux_io_sources_3_ready),
		.io_sources_3_valid(_s_axi__buffered_sourceBuffer_11_io_deq_valid),
		.io_sources_3_bits_data(_s_axi__buffered_sourceBuffer_11_io_deq_bits_data),
		.io_sources_3_bits_strb(_s_axi__buffered_sourceBuffer_11_io_deq_bits_strb),
		.io_sources_3_bits_last(_s_axi__buffered_sourceBuffer_11_io_deq_bits_last),
		.io_sources_4_ready(_write_mux_io_sources_4_ready),
		.io_sources_4_valid(_s_axi__buffered_sourceBuffer_14_io_deq_valid),
		.io_sources_4_bits_data(_s_axi__buffered_sourceBuffer_14_io_deq_bits_data),
		.io_sources_4_bits_strb(_s_axi__buffered_sourceBuffer_14_io_deq_bits_strb),
		.io_sources_4_bits_last(_s_axi__buffered_sourceBuffer_14_io_deq_bits_last),
		.io_sources_5_ready(_write_mux_io_sources_5_ready),
		.io_sources_5_valid(_s_axi__buffered_sourceBuffer_17_io_deq_valid),
		.io_sources_5_bits_data(_s_axi__buffered_sourceBuffer_17_io_deq_bits_data),
		.io_sources_5_bits_strb(_s_axi__buffered_sourceBuffer_17_io_deq_bits_strb),
		.io_sources_5_bits_last(_s_axi__buffered_sourceBuffer_17_io_deq_bits_last),
		.io_sources_6_ready(_write_mux_io_sources_6_ready),
		.io_sources_6_valid(_s_axi__buffered_sourceBuffer_20_io_deq_valid),
		.io_sources_6_bits_data(_s_axi__buffered_sourceBuffer_20_io_deq_bits_data),
		.io_sources_6_bits_strb(_s_axi__buffered_sourceBuffer_20_io_deq_bits_strb),
		.io_sources_6_bits_last(_s_axi__buffered_sourceBuffer_20_io_deq_bits_last),
		.io_sources_7_ready(_write_mux_io_sources_7_ready),
		.io_sources_7_valid(_s_axi__buffered_sourceBuffer_23_io_deq_valid),
		.io_sources_7_bits_data(_s_axi__buffered_sourceBuffer_23_io_deq_bits_data),
		.io_sources_7_bits_strb(_s_axi__buffered_sourceBuffer_23_io_deq_bits_strb),
		.io_sources_7_bits_last(_s_axi__buffered_sourceBuffer_23_io_deq_bits_last),
		.io_sources_8_ready(_write_mux_io_sources_8_ready),
		.io_sources_8_valid(_s_axi__buffered_sourceBuffer_26_io_deq_valid),
		.io_sources_8_bits_data(_s_axi__buffered_sourceBuffer_26_io_deq_bits_data),
		.io_sources_8_bits_strb(_s_axi__buffered_sourceBuffer_26_io_deq_bits_strb),
		.io_sources_8_bits_last(_s_axi__buffered_sourceBuffer_26_io_deq_bits_last),
		.io_sources_9_ready(_write_mux_io_sources_9_ready),
		.io_sources_9_valid(_s_axi__buffered_sourceBuffer_29_io_deq_valid),
		.io_sources_9_bits_data(_s_axi__buffered_sourceBuffer_29_io_deq_bits_data),
		.io_sources_9_bits_strb(_s_axi__buffered_sourceBuffer_29_io_deq_bits_strb),
		.io_sources_9_bits_last(_s_axi__buffered_sourceBuffer_29_io_deq_bits_last),
		.io_sources_10_ready(_write_mux_io_sources_10_ready),
		.io_sources_10_valid(_s_axi__buffered_sourceBuffer_32_io_deq_valid),
		.io_sources_10_bits_data(_s_axi__buffered_sourceBuffer_32_io_deq_bits_data),
		.io_sources_10_bits_strb(_s_axi__buffered_sourceBuffer_32_io_deq_bits_strb),
		.io_sources_10_bits_last(_s_axi__buffered_sourceBuffer_32_io_deq_bits_last),
		.io_sources_11_ready(_write_mux_io_sources_11_ready),
		.io_sources_11_valid(_s_axi__buffered_sourceBuffer_35_io_deq_valid),
		.io_sources_11_bits_data(_s_axi__buffered_sourceBuffer_35_io_deq_bits_data),
		.io_sources_11_bits_strb(_s_axi__buffered_sourceBuffer_35_io_deq_bits_strb),
		.io_sources_11_bits_last(_s_axi__buffered_sourceBuffer_35_io_deq_bits_last),
		.io_sources_12_ready(_write_mux_io_sources_12_ready),
		.io_sources_12_valid(_s_axi__buffered_sourceBuffer_38_io_deq_valid),
		.io_sources_12_bits_data(_s_axi__buffered_sourceBuffer_38_io_deq_bits_data),
		.io_sources_12_bits_strb(_s_axi__buffered_sourceBuffer_38_io_deq_bits_strb),
		.io_sources_12_bits_last(_s_axi__buffered_sourceBuffer_38_io_deq_bits_last),
		.io_sources_13_ready(_write_mux_io_sources_13_ready),
		.io_sources_13_valid(_s_axi__buffered_sourceBuffer_41_io_deq_valid),
		.io_sources_13_bits_data(_s_axi__buffered_sourceBuffer_41_io_deq_bits_data),
		.io_sources_13_bits_strb(_s_axi__buffered_sourceBuffer_41_io_deq_bits_strb),
		.io_sources_13_bits_last(_s_axi__buffered_sourceBuffer_41_io_deq_bits_last),
		.io_sources_14_ready(_write_mux_io_sources_14_ready),
		.io_sources_14_valid(_s_axi__buffered_sourceBuffer_44_io_deq_valid),
		.io_sources_14_bits_data(_s_axi__buffered_sourceBuffer_44_io_deq_bits_data),
		.io_sources_14_bits_strb(_s_axi__buffered_sourceBuffer_44_io_deq_bits_strb),
		.io_sources_14_bits_last(_s_axi__buffered_sourceBuffer_44_io_deq_bits_last),
		.io_sources_15_ready(_write_mux_io_sources_15_ready),
		.io_sources_15_valid(_s_axi__buffered_sourceBuffer_47_io_deq_valid),
		.io_sources_15_bits_data(_s_axi__buffered_sourceBuffer_47_io_deq_bits_data),
		.io_sources_15_bits_strb(_s_axi__buffered_sourceBuffer_47_io_deq_bits_strb),
		.io_sources_15_bits_last(_s_axi__buffered_sourceBuffer_47_io_deq_bits_last),
		.io_sources_16_ready(_write_mux_io_sources_16_ready),
		.io_sources_16_valid(_s_axi__buffered_sourceBuffer_50_io_deq_valid),
		.io_sources_16_bits_data(_s_axi__buffered_sourceBuffer_50_io_deq_bits_data),
		.io_sources_16_bits_strb(_s_axi__buffered_sourceBuffer_50_io_deq_bits_strb),
		.io_sources_16_bits_last(_s_axi__buffered_sourceBuffer_50_io_deq_bits_last),
		.io_sources_17_ready(_write_mux_io_sources_17_ready),
		.io_sources_17_valid(_s_axi__buffered_sourceBuffer_53_io_deq_valid),
		.io_sources_17_bits_data(_s_axi__buffered_sourceBuffer_53_io_deq_bits_data),
		.io_sources_17_bits_strb(_s_axi__buffered_sourceBuffer_53_io_deq_bits_strb),
		.io_sources_17_bits_last(_s_axi__buffered_sourceBuffer_53_io_deq_bits_last),
		.io_sources_18_ready(_write_mux_io_sources_18_ready),
		.io_sources_18_valid(_s_axi__buffered_sourceBuffer_56_io_deq_valid),
		.io_sources_18_bits_data(_s_axi__buffered_sourceBuffer_56_io_deq_bits_data),
		.io_sources_18_bits_strb(_s_axi__buffered_sourceBuffer_56_io_deq_bits_strb),
		.io_sources_18_bits_last(_s_axi__buffered_sourceBuffer_56_io_deq_bits_last),
		.io_sources_19_ready(_write_mux_io_sources_19_ready),
		.io_sources_19_valid(_s_axi__buffered_sourceBuffer_59_io_deq_valid),
		.io_sources_19_bits_data(_s_axi__buffered_sourceBuffer_59_io_deq_bits_data),
		.io_sources_19_bits_strb(_s_axi__buffered_sourceBuffer_59_io_deq_bits_strb),
		.io_sources_19_bits_last(_s_axi__buffered_sourceBuffer_59_io_deq_bits_last),
		.io_sources_20_ready(_write_mux_io_sources_20_ready),
		.io_sources_20_valid(_s_axi__buffered_sourceBuffer_62_io_deq_valid),
		.io_sources_20_bits_data(_s_axi__buffered_sourceBuffer_62_io_deq_bits_data),
		.io_sources_20_bits_strb(_s_axi__buffered_sourceBuffer_62_io_deq_bits_strb),
		.io_sources_20_bits_last(_s_axi__buffered_sourceBuffer_62_io_deq_bits_last),
		.io_sources_21_ready(_write_mux_io_sources_21_ready),
		.io_sources_21_valid(_s_axi__buffered_sourceBuffer_65_io_deq_valid),
		.io_sources_21_bits_data(_s_axi__buffered_sourceBuffer_65_io_deq_bits_data),
		.io_sources_21_bits_strb(_s_axi__buffered_sourceBuffer_65_io_deq_bits_strb),
		.io_sources_21_bits_last(_s_axi__buffered_sourceBuffer_65_io_deq_bits_last),
		.io_sources_22_ready(_write_mux_io_sources_22_ready),
		.io_sources_22_valid(_s_axi__buffered_sourceBuffer_68_io_deq_valid),
		.io_sources_22_bits_data(_s_axi__buffered_sourceBuffer_68_io_deq_bits_data),
		.io_sources_22_bits_strb(_s_axi__buffered_sourceBuffer_68_io_deq_bits_strb),
		.io_sources_22_bits_last(_s_axi__buffered_sourceBuffer_68_io_deq_bits_last),
		.io_sources_23_ready(_write_mux_io_sources_23_ready),
		.io_sources_23_valid(_s_axi__buffered_sourceBuffer_71_io_deq_valid),
		.io_sources_23_bits_data(_s_axi__buffered_sourceBuffer_71_io_deq_bits_data),
		.io_sources_23_bits_strb(_s_axi__buffered_sourceBuffer_71_io_deq_bits_strb),
		.io_sources_23_bits_last(_s_axi__buffered_sourceBuffer_71_io_deq_bits_last),
		.io_sources_24_ready(_write_mux_io_sources_24_ready),
		.io_sources_24_valid(_s_axi__buffered_sourceBuffer_74_io_deq_valid),
		.io_sources_24_bits_data(_s_axi__buffered_sourceBuffer_74_io_deq_bits_data),
		.io_sources_24_bits_strb(_s_axi__buffered_sourceBuffer_74_io_deq_bits_strb),
		.io_sources_24_bits_last(_s_axi__buffered_sourceBuffer_74_io_deq_bits_last),
		.io_sources_25_ready(_write_mux_io_sources_25_ready),
		.io_sources_25_valid(_s_axi__buffered_sourceBuffer_77_io_deq_valid),
		.io_sources_25_bits_data(_s_axi__buffered_sourceBuffer_77_io_deq_bits_data),
		.io_sources_25_bits_strb(_s_axi__buffered_sourceBuffer_77_io_deq_bits_strb),
		.io_sources_25_bits_last(_s_axi__buffered_sourceBuffer_77_io_deq_bits_last),
		.io_sources_26_ready(_write_mux_io_sources_26_ready),
		.io_sources_26_valid(_s_axi__buffered_sourceBuffer_80_io_deq_valid),
		.io_sources_26_bits_data(_s_axi__buffered_sourceBuffer_80_io_deq_bits_data),
		.io_sources_26_bits_strb(_s_axi__buffered_sourceBuffer_80_io_deq_bits_strb),
		.io_sources_26_bits_last(_s_axi__buffered_sourceBuffer_80_io_deq_bits_last),
		.io_sources_27_ready(_write_mux_io_sources_27_ready),
		.io_sources_27_valid(_s_axi__buffered_sourceBuffer_83_io_deq_valid),
		.io_sources_27_bits_data(_s_axi__buffered_sourceBuffer_83_io_deq_bits_data),
		.io_sources_27_bits_strb(_s_axi__buffered_sourceBuffer_83_io_deq_bits_strb),
		.io_sources_27_bits_last(_s_axi__buffered_sourceBuffer_83_io_deq_bits_last),
		.io_sources_28_ready(_write_mux_io_sources_28_ready),
		.io_sources_28_valid(_s_axi__buffered_sourceBuffer_86_io_deq_valid),
		.io_sources_28_bits_data(_s_axi__buffered_sourceBuffer_86_io_deq_bits_data),
		.io_sources_28_bits_strb(_s_axi__buffered_sourceBuffer_86_io_deq_bits_strb),
		.io_sources_28_bits_last(_s_axi__buffered_sourceBuffer_86_io_deq_bits_last),
		.io_sources_29_ready(_write_mux_io_sources_29_ready),
		.io_sources_29_valid(_s_axi__buffered_sourceBuffer_89_io_deq_valid),
		.io_sources_29_bits_data(_s_axi__buffered_sourceBuffer_89_io_deq_bits_data),
		.io_sources_29_bits_strb(_s_axi__buffered_sourceBuffer_89_io_deq_bits_strb),
		.io_sources_29_bits_last(_s_axi__buffered_sourceBuffer_89_io_deq_bits_last),
		.io_sources_30_ready(_write_mux_io_sources_30_ready),
		.io_sources_30_valid(_s_axi__buffered_sourceBuffer_92_io_deq_valid),
		.io_sources_30_bits_data(_s_axi__buffered_sourceBuffer_92_io_deq_bits_data),
		.io_sources_30_bits_strb(_s_axi__buffered_sourceBuffer_92_io_deq_bits_strb),
		.io_sources_30_bits_last(_s_axi__buffered_sourceBuffer_92_io_deq_bits_last),
		.io_sources_31_ready(_write_mux_io_sources_31_ready),
		.io_sources_31_valid(_s_axi__buffered_sourceBuffer_95_io_deq_valid),
		.io_sources_31_bits_data(_s_axi__buffered_sourceBuffer_95_io_deq_bits_data),
		.io_sources_31_bits_strb(_s_axi__buffered_sourceBuffer_95_io_deq_bits_strb),
		.io_sources_31_bits_last(_s_axi__buffered_sourceBuffer_95_io_deq_bits_last),
		.io_sink_ready(_m_axi__sourceBuffer_2_io_enq_ready),
		.io_sink_valid(_write_mux_io_sink_valid),
		.io_sink_bits_data(_write_mux_io_sink_bits_data),
		.io_sink_bits_strb(_write_mux_io_sink_bits_strb),
		.io_sink_bits_last(_write_mux_io_sink_bits_last),
		.io_select_ready(_write_mux_io_select_ready),
		.io_select_valid(_write_portQueue_io_deq_valid),
		.io_select_bits(_write_portQueue_io_deq_bits)
	);
	elasticDemux_10 write_demux(
		.io_source_ready(_write_demux_io_source_ready),
		.io_source_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_0),
		.io_sinks_0_ready(_s_axi__buffered_sinkBuffer_1_io_enq_ready),
		.io_sinks_0_valid(_write_demux_io_sinks_0_valid),
		.io_sinks_1_ready(_s_axi__buffered_sinkBuffer_3_io_enq_ready),
		.io_sinks_1_valid(_write_demux_io_sinks_1_valid),
		.io_sinks_2_ready(_s_axi__buffered_sinkBuffer_5_io_enq_ready),
		.io_sinks_2_valid(_write_demux_io_sinks_2_valid),
		.io_sinks_3_ready(_s_axi__buffered_sinkBuffer_7_io_enq_ready),
		.io_sinks_3_valid(_write_demux_io_sinks_3_valid),
		.io_sinks_4_ready(_s_axi__buffered_sinkBuffer_9_io_enq_ready),
		.io_sinks_4_valid(_write_demux_io_sinks_4_valid),
		.io_sinks_5_ready(_s_axi__buffered_sinkBuffer_11_io_enq_ready),
		.io_sinks_5_valid(_write_demux_io_sinks_5_valid),
		.io_sinks_6_ready(_s_axi__buffered_sinkBuffer_13_io_enq_ready),
		.io_sinks_6_valid(_write_demux_io_sinks_6_valid),
		.io_sinks_7_ready(_s_axi__buffered_sinkBuffer_15_io_enq_ready),
		.io_sinks_7_valid(_write_demux_io_sinks_7_valid),
		.io_sinks_8_ready(_s_axi__buffered_sinkBuffer_17_io_enq_ready),
		.io_sinks_8_valid(_write_demux_io_sinks_8_valid),
		.io_sinks_9_ready(_s_axi__buffered_sinkBuffer_19_io_enq_ready),
		.io_sinks_9_valid(_write_demux_io_sinks_9_valid),
		.io_sinks_10_ready(_s_axi__buffered_sinkBuffer_21_io_enq_ready),
		.io_sinks_10_valid(_write_demux_io_sinks_10_valid),
		.io_sinks_11_ready(_s_axi__buffered_sinkBuffer_23_io_enq_ready),
		.io_sinks_11_valid(_write_demux_io_sinks_11_valid),
		.io_sinks_12_ready(_s_axi__buffered_sinkBuffer_25_io_enq_ready),
		.io_sinks_12_valid(_write_demux_io_sinks_12_valid),
		.io_sinks_13_ready(_s_axi__buffered_sinkBuffer_27_io_enq_ready),
		.io_sinks_13_valid(_write_demux_io_sinks_13_valid),
		.io_sinks_14_ready(_s_axi__buffered_sinkBuffer_29_io_enq_ready),
		.io_sinks_14_valid(_write_demux_io_sinks_14_valid),
		.io_sinks_15_ready(_s_axi__buffered_sinkBuffer_31_io_enq_ready),
		.io_sinks_15_valid(_write_demux_io_sinks_15_valid),
		.io_sinks_16_ready(_s_axi__buffered_sinkBuffer_33_io_enq_ready),
		.io_sinks_16_valid(_write_demux_io_sinks_16_valid),
		.io_sinks_17_ready(_s_axi__buffered_sinkBuffer_35_io_enq_ready),
		.io_sinks_17_valid(_write_demux_io_sinks_17_valid),
		.io_sinks_18_ready(_s_axi__buffered_sinkBuffer_37_io_enq_ready),
		.io_sinks_18_valid(_write_demux_io_sinks_18_valid),
		.io_sinks_19_ready(_s_axi__buffered_sinkBuffer_39_io_enq_ready),
		.io_sinks_19_valid(_write_demux_io_sinks_19_valid),
		.io_sinks_20_ready(_s_axi__buffered_sinkBuffer_41_io_enq_ready),
		.io_sinks_20_valid(_write_demux_io_sinks_20_valid),
		.io_sinks_21_ready(_s_axi__buffered_sinkBuffer_43_io_enq_ready),
		.io_sinks_21_valid(_write_demux_io_sinks_21_valid),
		.io_sinks_22_ready(_s_axi__buffered_sinkBuffer_45_io_enq_ready),
		.io_sinks_22_valid(_write_demux_io_sinks_22_valid),
		.io_sinks_23_ready(_s_axi__buffered_sinkBuffer_47_io_enq_ready),
		.io_sinks_23_valid(_write_demux_io_sinks_23_valid),
		.io_sinks_24_ready(_s_axi__buffered_sinkBuffer_49_io_enq_ready),
		.io_sinks_24_valid(_write_demux_io_sinks_24_valid),
		.io_sinks_25_ready(_s_axi__buffered_sinkBuffer_51_io_enq_ready),
		.io_sinks_25_valid(_write_demux_io_sinks_25_valid),
		.io_sinks_26_ready(_s_axi__buffered_sinkBuffer_53_io_enq_ready),
		.io_sinks_26_valid(_write_demux_io_sinks_26_valid),
		.io_sinks_27_ready(_s_axi__buffered_sinkBuffer_55_io_enq_ready),
		.io_sinks_27_valid(_write_demux_io_sinks_27_valid),
		.io_sinks_28_ready(_s_axi__buffered_sinkBuffer_57_io_enq_ready),
		.io_sinks_28_valid(_write_demux_io_sinks_28_valid),
		.io_sinks_29_ready(_s_axi__buffered_sinkBuffer_59_io_enq_ready),
		.io_sinks_29_valid(_write_demux_io_sinks_29_valid),
		.io_sinks_30_ready(_s_axi__buffered_sinkBuffer_61_io_enq_ready),
		.io_sinks_30_valid(_write_demux_io_sinks_30_valid),
		.io_sinks_31_ready(_s_axi__buffered_sinkBuffer_63_io_enq_ready),
		.io_sinks_31_valid(_write_demux_io_sinks_31_valid),
		.io_select_ready(_write_demux_io_select_ready),
		.io_select_valid(_m_axi__sinkBuffer_1_io_deq_valid & ~write_eagerFork_regs_1),
		.io_select_bits(_m_axi__sinkBuffer_1_io_deq_bits_id)
	);
endmodule
module Counter64 (
	clock,
	reset,
	io_signals_0,
	io_signals_1,
	io_signals_2,
	io_signals_3,
	io_signals_4,
	io_signals_5,
	io_signals_6,
	io_signals_7,
	io_signals_8,
	io_signals_9,
	io_signals_10,
	io_signals_11,
	io_signals_12,
	io_signals_13,
	io_signals_14,
	io_signals_15,
	io_signals_16,
	io_signals_17,
	io_signals_18,
	io_signals_19,
	io_signals_20,
	io_signals_21,
	io_signals_22,
	io_signals_23,
	io_signals_24,
	io_signals_25,
	io_signals_26,
	io_signals_27,
	io_signals_28,
	io_signals_29,
	io_signals_30,
	io_signals_31,
	io_signals_32,
	io_signals_33,
	io_signals_34,
	io_signals_35,
	io_signals_36,
	io_signals_37,
	io_signals_38,
	io_signals_39,
	io_signals_40,
	io_signals_41,
	io_signals_42,
	io_signals_43,
	io_signals_44,
	io_signals_45,
	io_signals_46,
	io_signals_47,
	io_signals_48,
	io_signals_49,
	io_signals_50,
	io_signals_51,
	io_signals_52,
	io_signals_53,
	io_signals_54,
	io_signals_55,
	io_signals_56,
	io_signals_57,
	io_signals_58,
	io_signals_59,
	io_signals_60,
	io_signals_61,
	io_signals_62,
	io_signals_63,
	io_signals_64,
	io_signals_65,
	io_signals_66,
	io_signals_67,
	io_signals_68,
	io_signals_69,
	io_signals_70,
	io_signals_71,
	io_signals_72,
	io_signals_73,
	io_signals_74,
	io_signals_75,
	io_signals_76,
	io_signals_77,
	io_signals_78,
	io_signals_79,
	io_signals_80,
	io_signals_81,
	io_signals_82,
	io_signals_83,
	io_signals_84,
	io_signals_85,
	io_signals_86,
	io_signals_87,
	io_signals_88,
	io_signals_89,
	io_signals_90,
	io_signals_91,
	io_signals_92,
	io_signals_93,
	io_signals_94,
	io_signals_95,
	io_signals_96,
	io_signals_97,
	io_signals_98,
	io_signals_99,
	io_signals_100,
	io_signals_101,
	io_signals_102,
	io_signals_103,
	io_signals_104,
	io_signals_105,
	io_signals_106,
	io_signals_107,
	io_signals_108,
	io_signals_109,
	io_signals_110,
	io_signals_111,
	io_signals_112,
	io_signals_113,
	io_signals_114,
	io_signals_115,
	io_signals_116,
	io_signals_117,
	io_signals_118,
	io_signals_119,
	io_signals_120,
	io_signals_121,
	io_signals_122,
	io_signals_123,
	io_signals_124,
	io_signals_125,
	io_signals_126,
	io_signals_127,
	io_counter
);
	input clock;
	input reset;
	input io_signals_0;
	input io_signals_1;
	input io_signals_2;
	input io_signals_3;
	input io_signals_4;
	input io_signals_5;
	input io_signals_6;
	input io_signals_7;
	input io_signals_8;
	input io_signals_9;
	input io_signals_10;
	input io_signals_11;
	input io_signals_12;
	input io_signals_13;
	input io_signals_14;
	input io_signals_15;
	input io_signals_16;
	input io_signals_17;
	input io_signals_18;
	input io_signals_19;
	input io_signals_20;
	input io_signals_21;
	input io_signals_22;
	input io_signals_23;
	input io_signals_24;
	input io_signals_25;
	input io_signals_26;
	input io_signals_27;
	input io_signals_28;
	input io_signals_29;
	input io_signals_30;
	input io_signals_31;
	input io_signals_32;
	input io_signals_33;
	input io_signals_34;
	input io_signals_35;
	input io_signals_36;
	input io_signals_37;
	input io_signals_38;
	input io_signals_39;
	input io_signals_40;
	input io_signals_41;
	input io_signals_42;
	input io_signals_43;
	input io_signals_44;
	input io_signals_45;
	input io_signals_46;
	input io_signals_47;
	input io_signals_48;
	input io_signals_49;
	input io_signals_50;
	input io_signals_51;
	input io_signals_52;
	input io_signals_53;
	input io_signals_54;
	input io_signals_55;
	input io_signals_56;
	input io_signals_57;
	input io_signals_58;
	input io_signals_59;
	input io_signals_60;
	input io_signals_61;
	input io_signals_62;
	input io_signals_63;
	input io_signals_64;
	input io_signals_65;
	input io_signals_66;
	input io_signals_67;
	input io_signals_68;
	input io_signals_69;
	input io_signals_70;
	input io_signals_71;
	input io_signals_72;
	input io_signals_73;
	input io_signals_74;
	input io_signals_75;
	input io_signals_76;
	input io_signals_77;
	input io_signals_78;
	input io_signals_79;
	input io_signals_80;
	input io_signals_81;
	input io_signals_82;
	input io_signals_83;
	input io_signals_84;
	input io_signals_85;
	input io_signals_86;
	input io_signals_87;
	input io_signals_88;
	input io_signals_89;
	input io_signals_90;
	input io_signals_91;
	input io_signals_92;
	input io_signals_93;
	input io_signals_94;
	input io_signals_95;
	input io_signals_96;
	input io_signals_97;
	input io_signals_98;
	input io_signals_99;
	input io_signals_100;
	input io_signals_101;
	input io_signals_102;
	input io_signals_103;
	input io_signals_104;
	input io_signals_105;
	input io_signals_106;
	input io_signals_107;
	input io_signals_108;
	input io_signals_109;
	input io_signals_110;
	input io_signals_111;
	input io_signals_112;
	input io_signals_113;
	input io_signals_114;
	input io_signals_115;
	input io_signals_116;
	input io_signals_117;
	input io_signals_118;
	input io_signals_119;
	input io_signals_120;
	input io_signals_121;
	input io_signals_122;
	input io_signals_123;
	input io_signals_124;
	input io_signals_125;
	input io_signals_126;
	input io_signals_127;
	output wire [63:0] io_counter;
	reg [63:0] counter;
	always @(posedge clock)
		if (reset)
			counter <= 64'h0000000000000000;
		else
			counter <= counter + {56'h00000000000000, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_0} + {1'h0, io_signals_1}} + {1'h0, {1'h0, io_signals_2} + {1'h0, io_signals_3}}} + {1'h0, {1'h0, {1'h0, io_signals_4} + {1'h0, io_signals_5}} + {1'h0, {1'h0, io_signals_6} + {1'h0, io_signals_7}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_8} + {1'h0, io_signals_9}} + {1'h0, {1'h0, io_signals_10} + {1'h0, io_signals_11}}} + {1'h0, {1'h0, {1'h0, io_signals_12} + {1'h0, io_signals_13}} + {1'h0, {1'h0, io_signals_14} + {1'h0, io_signals_15}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_16} + {1'h0, io_signals_17}} + {1'h0, {1'h0, io_signals_18} + {1'h0, io_signals_19}}} + {1'h0, {1'h0, {1'h0, io_signals_20} + {1'h0, io_signals_21}} + {1'h0, {1'h0, io_signals_22} + {1'h0, io_signals_23}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_24} + {1'h0, io_signals_25}} + {1'h0, {1'h0, io_signals_26} + {1'h0, io_signals_27}}} + {1'h0, {1'h0, {1'h0, io_signals_28} + {1'h0, io_signals_29}} + {1'h0, {1'h0, io_signals_30} + {1'h0, io_signals_31}}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_32} + {1'h0, io_signals_33}} + {1'h0, {1'h0, io_signals_34} + {1'h0, io_signals_35}}} + {1'h0, {1'h0, {1'h0, io_signals_36} + {1'h0, io_signals_37}} + {1'h0, {1'h0, io_signals_38} + {1'h0, io_signals_39}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_40} + {1'h0, io_signals_41}} + {1'h0, {1'h0, io_signals_42} + {1'h0, io_signals_43}}} + {1'h0, {1'h0, {1'h0, io_signals_44} + {1'h0, io_signals_45}} + {1'h0, {1'h0, io_signals_46} + {1'h0, io_signals_47}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_48} + {1'h0, io_signals_49}} + {1'h0, {1'h0, io_signals_50} + {1'h0, io_signals_51}}} + {1'h0, {1'h0, {1'h0, io_signals_52} + {1'h0, io_signals_53}} + {1'h0, {1'h0, io_signals_54} + {1'h0, io_signals_55}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_56} + {1'h0, io_signals_57}} + {1'h0, {1'h0, io_signals_58} + {1'h0, io_signals_59}}} + {1'h0, {1'h0, {1'h0, io_signals_60} + {1'h0, io_signals_61}} + {1'h0, {1'h0, io_signals_62} + {1'h0, io_signals_63}}}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_64} + {1'h0, io_signals_65}} + {1'h0, {1'h0, io_signals_66} + {1'h0, io_signals_67}}} + {1'h0, {1'h0, {1'h0, io_signals_68} + {1'h0, io_signals_69}} + {1'h0, {1'h0, io_signals_70} + {1'h0, io_signals_71}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_72} + {1'h0, io_signals_73}} + {1'h0, {1'h0, io_signals_74} + {1'h0, io_signals_75}}} + {1'h0, {1'h0, {1'h0, io_signals_76} + {1'h0, io_signals_77}} + {1'h0, {1'h0, io_signals_78} + {1'h0, io_signals_79}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_80} + {1'h0, io_signals_81}} + {1'h0, {1'h0, io_signals_82} + {1'h0, io_signals_83}}} + {1'h0, {1'h0, {1'h0, io_signals_84} + {1'h0, io_signals_85}} + {1'h0, {1'h0, io_signals_86} + {1'h0, io_signals_87}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_88} + {1'h0, io_signals_89}} + {1'h0, {1'h0, io_signals_90} + {1'h0, io_signals_91}}} + {1'h0, {1'h0, {1'h0, io_signals_92} + {1'h0, io_signals_93}} + {1'h0, {1'h0, io_signals_94} + {1'h0, io_signals_95}}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_96} + {1'h0, io_signals_97}} + {1'h0, {1'h0, io_signals_98} + {1'h0, io_signals_99}}} + {1'h0, {1'h0, {1'h0, io_signals_100} + {1'h0, io_signals_101}} + {1'h0, {1'h0, io_signals_102} + {1'h0, io_signals_103}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_104} + {1'h0, io_signals_105}} + {1'h0, {1'h0, io_signals_106} + {1'h0, io_signals_107}}} + {1'h0, {1'h0, {1'h0, io_signals_108} + {1'h0, io_signals_109}} + {1'h0, {1'h0, io_signals_110} + {1'h0, io_signals_111}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_112} + {1'h0, io_signals_113}} + {1'h0, {1'h0, io_signals_114} + {1'h0, io_signals_115}}} + {1'h0, {1'h0, {1'h0, io_signals_116} + {1'h0, io_signals_117}} + {1'h0, {1'h0, io_signals_118} + {1'h0, io_signals_119}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_120} + {1'h0, io_signals_121}} + {1'h0, {1'h0, io_signals_122} + {1'h0, io_signals_123}}} + {1'h0, {1'h0, {1'h0, io_signals_124} + {1'h0, io_signals_125}} + {1'h0, {1'h0, io_signals_126} + {1'h0, io_signals_127}}}}}}}};
	assign io_counter = counter;
endmodule
module ArgumentNotifier (
	clock,
	reset,
	io_export_argIn_0_TREADY,
	io_export_argIn_0_TVALID,
	io_export_argIn_0_TDATA,
	io_export_argIn_1_TREADY,
	io_export_argIn_1_TVALID,
	io_export_argIn_1_TDATA,
	io_export_argIn_2_TREADY,
	io_export_argIn_2_TVALID,
	io_export_argIn_2_TDATA,
	io_export_argIn_3_TREADY,
	io_export_argIn_3_TVALID,
	io_export_argIn_3_TDATA,
	io_export_argIn_4_TREADY,
	io_export_argIn_4_TVALID,
	io_export_argIn_4_TDATA,
	io_export_argIn_5_TREADY,
	io_export_argIn_5_TVALID,
	io_export_argIn_5_TDATA,
	io_export_argIn_6_TREADY,
	io_export_argIn_6_TVALID,
	io_export_argIn_6_TDATA,
	io_export_argIn_7_TREADY,
	io_export_argIn_7_TVALID,
	io_export_argIn_7_TDATA,
	io_export_argIn_8_TREADY,
	io_export_argIn_8_TVALID,
	io_export_argIn_8_TDATA,
	io_export_argIn_9_TREADY,
	io_export_argIn_9_TVALID,
	io_export_argIn_9_TDATA,
	io_export_argIn_10_TREADY,
	io_export_argIn_10_TVALID,
	io_export_argIn_10_TDATA,
	io_export_argIn_11_TREADY,
	io_export_argIn_11_TVALID,
	io_export_argIn_11_TDATA,
	io_export_argIn_12_TREADY,
	io_export_argIn_12_TVALID,
	io_export_argIn_12_TDATA,
	io_export_argIn_13_TREADY,
	io_export_argIn_13_TVALID,
	io_export_argIn_13_TDATA,
	io_export_argIn_14_TREADY,
	io_export_argIn_14_TVALID,
	io_export_argIn_14_TDATA,
	io_export_argIn_15_TREADY,
	io_export_argIn_15_TVALID,
	io_export_argIn_15_TDATA,
	io_export_argIn_16_TREADY,
	io_export_argIn_16_TVALID,
	io_export_argIn_16_TDATA,
	io_export_argIn_17_TREADY,
	io_export_argIn_17_TVALID,
	io_export_argIn_17_TDATA,
	io_export_argIn_18_TREADY,
	io_export_argIn_18_TVALID,
	io_export_argIn_18_TDATA,
	io_export_argIn_19_TREADY,
	io_export_argIn_19_TVALID,
	io_export_argIn_19_TDATA,
	io_export_argIn_20_TREADY,
	io_export_argIn_20_TVALID,
	io_export_argIn_20_TDATA,
	io_export_argIn_21_TREADY,
	io_export_argIn_21_TVALID,
	io_export_argIn_21_TDATA,
	io_export_argIn_22_TREADY,
	io_export_argIn_22_TVALID,
	io_export_argIn_22_TDATA,
	io_export_argIn_23_TREADY,
	io_export_argIn_23_TVALID,
	io_export_argIn_23_TDATA,
	io_export_argIn_24_TREADY,
	io_export_argIn_24_TVALID,
	io_export_argIn_24_TDATA,
	io_export_argIn_25_TREADY,
	io_export_argIn_25_TVALID,
	io_export_argIn_25_TDATA,
	io_export_argIn_26_TREADY,
	io_export_argIn_26_TVALID,
	io_export_argIn_26_TDATA,
	io_export_argIn_27_TREADY,
	io_export_argIn_27_TVALID,
	io_export_argIn_27_TDATA,
	io_export_argIn_28_TREADY,
	io_export_argIn_28_TVALID,
	io_export_argIn_28_TDATA,
	io_export_argIn_29_TREADY,
	io_export_argIn_29_TVALID,
	io_export_argIn_29_TDATA,
	io_export_argIn_30_TREADY,
	io_export_argIn_30_TVALID,
	io_export_argIn_30_TDATA,
	io_export_argIn_31_TREADY,
	io_export_argIn_31_TVALID,
	io_export_argIn_31_TDATA,
	io_export_argIn_32_TREADY,
	io_export_argIn_32_TVALID,
	io_export_argIn_32_TDATA,
	io_export_argIn_33_TREADY,
	io_export_argIn_33_TVALID,
	io_export_argIn_33_TDATA,
	io_export_argIn_34_TREADY,
	io_export_argIn_34_TVALID,
	io_export_argIn_34_TDATA,
	io_export_argIn_35_TREADY,
	io_export_argIn_35_TVALID,
	io_export_argIn_35_TDATA,
	io_export_argIn_36_TREADY,
	io_export_argIn_36_TVALID,
	io_export_argIn_36_TDATA,
	io_export_argIn_37_TREADY,
	io_export_argIn_37_TVALID,
	io_export_argIn_37_TDATA,
	io_export_argIn_38_TREADY,
	io_export_argIn_38_TVALID,
	io_export_argIn_38_TDATA,
	io_export_argIn_39_TREADY,
	io_export_argIn_39_TVALID,
	io_export_argIn_39_TDATA,
	io_export_argIn_40_TREADY,
	io_export_argIn_40_TVALID,
	io_export_argIn_40_TDATA,
	io_export_argIn_41_TREADY,
	io_export_argIn_41_TVALID,
	io_export_argIn_41_TDATA,
	io_export_argIn_42_TREADY,
	io_export_argIn_42_TVALID,
	io_export_argIn_42_TDATA,
	io_export_argIn_43_TREADY,
	io_export_argIn_43_TVALID,
	io_export_argIn_43_TDATA,
	io_export_argIn_44_TREADY,
	io_export_argIn_44_TVALID,
	io_export_argIn_44_TDATA,
	io_export_argIn_45_TREADY,
	io_export_argIn_45_TVALID,
	io_export_argIn_45_TDATA,
	io_export_argIn_46_TREADY,
	io_export_argIn_46_TVALID,
	io_export_argIn_46_TDATA,
	io_export_argIn_47_TREADY,
	io_export_argIn_47_TVALID,
	io_export_argIn_47_TDATA,
	io_export_argIn_48_TREADY,
	io_export_argIn_48_TVALID,
	io_export_argIn_48_TDATA,
	io_export_argIn_49_TREADY,
	io_export_argIn_49_TVALID,
	io_export_argIn_49_TDATA,
	io_export_argIn_50_TREADY,
	io_export_argIn_50_TVALID,
	io_export_argIn_50_TDATA,
	io_export_argIn_51_TREADY,
	io_export_argIn_51_TVALID,
	io_export_argIn_51_TDATA,
	io_export_argIn_52_TREADY,
	io_export_argIn_52_TVALID,
	io_export_argIn_52_TDATA,
	io_export_argIn_53_TREADY,
	io_export_argIn_53_TVALID,
	io_export_argIn_53_TDATA,
	io_export_argIn_54_TREADY,
	io_export_argIn_54_TVALID,
	io_export_argIn_54_TDATA,
	io_export_argIn_55_TREADY,
	io_export_argIn_55_TVALID,
	io_export_argIn_55_TDATA,
	io_export_argIn_56_TREADY,
	io_export_argIn_56_TVALID,
	io_export_argIn_56_TDATA,
	io_export_argIn_57_TREADY,
	io_export_argIn_57_TVALID,
	io_export_argIn_57_TDATA,
	io_export_argIn_58_TREADY,
	io_export_argIn_58_TVALID,
	io_export_argIn_58_TDATA,
	io_export_argIn_59_TREADY,
	io_export_argIn_59_TVALID,
	io_export_argIn_59_TDATA,
	io_export_argIn_60_TREADY,
	io_export_argIn_60_TVALID,
	io_export_argIn_60_TDATA,
	io_export_argIn_61_TREADY,
	io_export_argIn_61_TVALID,
	io_export_argIn_61_TDATA,
	io_export_argIn_62_TREADY,
	io_export_argIn_62_TVALID,
	io_export_argIn_62_TDATA,
	io_export_argIn_63_TREADY,
	io_export_argIn_63_TVALID,
	io_export_argIn_63_TDATA,
	io_export_argIn_64_TREADY,
	io_export_argIn_64_TVALID,
	io_export_argIn_64_TDATA,
	io_export_argIn_65_TREADY,
	io_export_argIn_65_TVALID,
	io_export_argIn_65_TDATA,
	io_export_argIn_66_TREADY,
	io_export_argIn_66_TVALID,
	io_export_argIn_66_TDATA,
	io_export_argIn_67_TREADY,
	io_export_argIn_67_TVALID,
	io_export_argIn_67_TDATA,
	io_export_argIn_68_TREADY,
	io_export_argIn_68_TVALID,
	io_export_argIn_68_TDATA,
	io_export_argIn_69_TREADY,
	io_export_argIn_69_TVALID,
	io_export_argIn_69_TDATA,
	io_export_argIn_70_TREADY,
	io_export_argIn_70_TVALID,
	io_export_argIn_70_TDATA,
	io_export_argIn_71_TREADY,
	io_export_argIn_71_TVALID,
	io_export_argIn_71_TDATA,
	io_export_argIn_72_TREADY,
	io_export_argIn_72_TVALID,
	io_export_argIn_72_TDATA,
	io_export_argIn_73_TREADY,
	io_export_argIn_73_TVALID,
	io_export_argIn_73_TDATA,
	io_export_argIn_74_TREADY,
	io_export_argIn_74_TVALID,
	io_export_argIn_74_TDATA,
	io_export_argIn_75_TREADY,
	io_export_argIn_75_TVALID,
	io_export_argIn_75_TDATA,
	io_export_argIn_76_TREADY,
	io_export_argIn_76_TVALID,
	io_export_argIn_76_TDATA,
	io_export_argIn_77_TREADY,
	io_export_argIn_77_TVALID,
	io_export_argIn_77_TDATA,
	io_export_argIn_78_TREADY,
	io_export_argIn_78_TVALID,
	io_export_argIn_78_TDATA,
	io_export_argIn_79_TREADY,
	io_export_argIn_79_TVALID,
	io_export_argIn_79_TDATA,
	io_export_argIn_80_TREADY,
	io_export_argIn_80_TVALID,
	io_export_argIn_80_TDATA,
	io_export_argIn_81_TREADY,
	io_export_argIn_81_TVALID,
	io_export_argIn_81_TDATA,
	io_export_argIn_82_TREADY,
	io_export_argIn_82_TVALID,
	io_export_argIn_82_TDATA,
	io_export_argIn_83_TREADY,
	io_export_argIn_83_TVALID,
	io_export_argIn_83_TDATA,
	io_export_argIn_84_TREADY,
	io_export_argIn_84_TVALID,
	io_export_argIn_84_TDATA,
	io_export_argIn_85_TREADY,
	io_export_argIn_85_TVALID,
	io_export_argIn_85_TDATA,
	io_export_argIn_86_TREADY,
	io_export_argIn_86_TVALID,
	io_export_argIn_86_TDATA,
	io_export_argIn_87_TREADY,
	io_export_argIn_87_TVALID,
	io_export_argIn_87_TDATA,
	io_export_argIn_88_TREADY,
	io_export_argIn_88_TVALID,
	io_export_argIn_88_TDATA,
	io_export_argIn_89_TREADY,
	io_export_argIn_89_TVALID,
	io_export_argIn_89_TDATA,
	io_export_argIn_90_TREADY,
	io_export_argIn_90_TVALID,
	io_export_argIn_90_TDATA,
	io_export_argIn_91_TREADY,
	io_export_argIn_91_TVALID,
	io_export_argIn_91_TDATA,
	io_export_argIn_92_TREADY,
	io_export_argIn_92_TVALID,
	io_export_argIn_92_TDATA,
	io_export_argIn_93_TREADY,
	io_export_argIn_93_TVALID,
	io_export_argIn_93_TDATA,
	io_export_argIn_94_TREADY,
	io_export_argIn_94_TVALID,
	io_export_argIn_94_TDATA,
	io_export_argIn_95_TREADY,
	io_export_argIn_95_TVALID,
	io_export_argIn_95_TDATA,
	io_export_argIn_96_TREADY,
	io_export_argIn_96_TVALID,
	io_export_argIn_96_TDATA,
	io_export_argIn_97_TREADY,
	io_export_argIn_97_TVALID,
	io_export_argIn_97_TDATA,
	io_export_argIn_98_TREADY,
	io_export_argIn_98_TVALID,
	io_export_argIn_98_TDATA,
	io_export_argIn_99_TREADY,
	io_export_argIn_99_TVALID,
	io_export_argIn_99_TDATA,
	io_export_argIn_100_TREADY,
	io_export_argIn_100_TVALID,
	io_export_argIn_100_TDATA,
	io_export_argIn_101_TREADY,
	io_export_argIn_101_TVALID,
	io_export_argIn_101_TDATA,
	io_export_argIn_102_TREADY,
	io_export_argIn_102_TVALID,
	io_export_argIn_102_TDATA,
	io_export_argIn_103_TREADY,
	io_export_argIn_103_TVALID,
	io_export_argIn_103_TDATA,
	io_export_argIn_104_TREADY,
	io_export_argIn_104_TVALID,
	io_export_argIn_104_TDATA,
	io_export_argIn_105_TREADY,
	io_export_argIn_105_TVALID,
	io_export_argIn_105_TDATA,
	io_export_argIn_106_TREADY,
	io_export_argIn_106_TVALID,
	io_export_argIn_106_TDATA,
	io_export_argIn_107_TREADY,
	io_export_argIn_107_TVALID,
	io_export_argIn_107_TDATA,
	io_export_argIn_108_TREADY,
	io_export_argIn_108_TVALID,
	io_export_argIn_108_TDATA,
	io_export_argIn_109_TREADY,
	io_export_argIn_109_TVALID,
	io_export_argIn_109_TDATA,
	io_export_argIn_110_TREADY,
	io_export_argIn_110_TVALID,
	io_export_argIn_110_TDATA,
	io_export_argIn_111_TREADY,
	io_export_argIn_111_TVALID,
	io_export_argIn_111_TDATA,
	io_export_argIn_112_TREADY,
	io_export_argIn_112_TVALID,
	io_export_argIn_112_TDATA,
	io_export_argIn_113_TREADY,
	io_export_argIn_113_TVALID,
	io_export_argIn_113_TDATA,
	io_export_argIn_114_TREADY,
	io_export_argIn_114_TVALID,
	io_export_argIn_114_TDATA,
	io_export_argIn_115_TREADY,
	io_export_argIn_115_TVALID,
	io_export_argIn_115_TDATA,
	io_export_argIn_116_TREADY,
	io_export_argIn_116_TVALID,
	io_export_argIn_116_TDATA,
	io_export_argIn_117_TREADY,
	io_export_argIn_117_TVALID,
	io_export_argIn_117_TDATA,
	io_export_argIn_118_TREADY,
	io_export_argIn_118_TVALID,
	io_export_argIn_118_TDATA,
	io_export_argIn_119_TREADY,
	io_export_argIn_119_TVALID,
	io_export_argIn_119_TDATA,
	io_export_argIn_120_TREADY,
	io_export_argIn_120_TVALID,
	io_export_argIn_120_TDATA,
	io_export_argIn_121_TREADY,
	io_export_argIn_121_TVALID,
	io_export_argIn_121_TDATA,
	io_export_argIn_122_TREADY,
	io_export_argIn_122_TVALID,
	io_export_argIn_122_TDATA,
	io_export_argIn_123_TREADY,
	io_export_argIn_123_TVALID,
	io_export_argIn_123_TDATA,
	io_export_argIn_124_TREADY,
	io_export_argIn_124_TVALID,
	io_export_argIn_124_TDATA,
	io_export_argIn_125_TREADY,
	io_export_argIn_125_TVALID,
	io_export_argIn_125_TDATA,
	io_export_argIn_126_TREADY,
	io_export_argIn_126_TVALID,
	io_export_argIn_126_TDATA,
	io_export_argIn_127_TREADY,
	io_export_argIn_127_TVALID,
	io_export_argIn_127_TDATA,
	connStealNtw_0_ctrl_serveStealReq_valid,
	connStealNtw_0_ctrl_serveStealReq_ready,
	connStealNtw_0_data_qOutTask_ready,
	connStealNtw_0_data_qOutTask_valid,
	connStealNtw_0_data_qOutTask_bits,
	connStealNtw_1_ctrl_serveStealReq_valid,
	connStealNtw_1_ctrl_serveStealReq_ready,
	connStealNtw_1_data_qOutTask_ready,
	connStealNtw_1_data_qOutTask_valid,
	connStealNtw_1_data_qOutTask_bits,
	connStealNtw_2_ctrl_serveStealReq_valid,
	connStealNtw_2_ctrl_serveStealReq_ready,
	connStealNtw_2_data_qOutTask_ready,
	connStealNtw_2_data_qOutTask_valid,
	connStealNtw_2_data_qOutTask_bits,
	connStealNtw_3_ctrl_serveStealReq_valid,
	connStealNtw_3_ctrl_serveStealReq_ready,
	connStealNtw_3_data_qOutTask_ready,
	connStealNtw_3_data_qOutTask_valid,
	connStealNtw_3_data_qOutTask_bits,
	connStealNtw_4_ctrl_serveStealReq_valid,
	connStealNtw_4_ctrl_serveStealReq_ready,
	connStealNtw_4_data_qOutTask_ready,
	connStealNtw_4_data_qOutTask_valid,
	connStealNtw_4_data_qOutTask_bits,
	connStealNtw_5_ctrl_serveStealReq_valid,
	connStealNtw_5_ctrl_serveStealReq_ready,
	connStealNtw_5_data_qOutTask_ready,
	connStealNtw_5_data_qOutTask_valid,
	connStealNtw_5_data_qOutTask_bits,
	connStealNtw_6_ctrl_serveStealReq_valid,
	connStealNtw_6_ctrl_serveStealReq_ready,
	connStealNtw_6_data_qOutTask_ready,
	connStealNtw_6_data_qOutTask_valid,
	connStealNtw_6_data_qOutTask_bits,
	connStealNtw_7_ctrl_serveStealReq_valid,
	connStealNtw_7_ctrl_serveStealReq_ready,
	connStealNtw_7_data_qOutTask_ready,
	connStealNtw_7_data_qOutTask_valid,
	connStealNtw_7_data_qOutTask_bits,
	connStealNtw_8_ctrl_serveStealReq_valid,
	connStealNtw_8_ctrl_serveStealReq_ready,
	connStealNtw_8_data_qOutTask_ready,
	connStealNtw_8_data_qOutTask_valid,
	connStealNtw_8_data_qOutTask_bits,
	connStealNtw_9_ctrl_serveStealReq_valid,
	connStealNtw_9_ctrl_serveStealReq_ready,
	connStealNtw_9_data_qOutTask_ready,
	connStealNtw_9_data_qOutTask_valid,
	connStealNtw_9_data_qOutTask_bits,
	connStealNtw_10_ctrl_serveStealReq_valid,
	connStealNtw_10_ctrl_serveStealReq_ready,
	connStealNtw_10_data_qOutTask_ready,
	connStealNtw_10_data_qOutTask_valid,
	connStealNtw_10_data_qOutTask_bits,
	connStealNtw_11_ctrl_serveStealReq_valid,
	connStealNtw_11_ctrl_serveStealReq_ready,
	connStealNtw_11_data_qOutTask_ready,
	connStealNtw_11_data_qOutTask_valid,
	connStealNtw_11_data_qOutTask_bits,
	connStealNtw_12_ctrl_serveStealReq_valid,
	connStealNtw_12_ctrl_serveStealReq_ready,
	connStealNtw_12_data_qOutTask_ready,
	connStealNtw_12_data_qOutTask_valid,
	connStealNtw_12_data_qOutTask_bits,
	connStealNtw_13_ctrl_serveStealReq_valid,
	connStealNtw_13_ctrl_serveStealReq_ready,
	connStealNtw_13_data_qOutTask_ready,
	connStealNtw_13_data_qOutTask_valid,
	connStealNtw_13_data_qOutTask_bits,
	connStealNtw_14_ctrl_serveStealReq_valid,
	connStealNtw_14_ctrl_serveStealReq_ready,
	connStealNtw_14_data_qOutTask_ready,
	connStealNtw_14_data_qOutTask_valid,
	connStealNtw_14_data_qOutTask_bits,
	connStealNtw_15_ctrl_serveStealReq_valid,
	connStealNtw_15_ctrl_serveStealReq_ready,
	connStealNtw_15_data_qOutTask_ready,
	connStealNtw_15_data_qOutTask_valid,
	connStealNtw_15_data_qOutTask_bits,
	axi_full_argRoute_0_ar_ready,
	axi_full_argRoute_0_ar_valid,
	axi_full_argRoute_0_ar_bits_id,
	axi_full_argRoute_0_ar_bits_addr,
	axi_full_argRoute_0_ar_bits_len,
	axi_full_argRoute_0_ar_bits_size,
	axi_full_argRoute_0_ar_bits_burst,
	axi_full_argRoute_0_ar_bits_lock,
	axi_full_argRoute_0_ar_bits_cache,
	axi_full_argRoute_0_ar_bits_prot,
	axi_full_argRoute_0_ar_bits_qos,
	axi_full_argRoute_0_ar_bits_region,
	axi_full_argRoute_0_r_ready,
	axi_full_argRoute_0_r_valid,
	axi_full_argRoute_0_r_bits_id,
	axi_full_argRoute_0_r_bits_data,
	axi_full_argRoute_0_r_bits_resp,
	axi_full_argRoute_0_r_bits_last,
	axi_full_argRoute_0_aw_ready,
	axi_full_argRoute_0_aw_valid,
	axi_full_argRoute_0_aw_bits_id,
	axi_full_argRoute_0_aw_bits_addr,
	axi_full_argRoute_0_aw_bits_len,
	axi_full_argRoute_0_aw_bits_size,
	axi_full_argRoute_0_aw_bits_burst,
	axi_full_argRoute_0_aw_bits_lock,
	axi_full_argRoute_0_aw_bits_cache,
	axi_full_argRoute_0_aw_bits_prot,
	axi_full_argRoute_0_aw_bits_qos,
	axi_full_argRoute_0_aw_bits_region,
	axi_full_argRoute_0_w_ready,
	axi_full_argRoute_0_w_valid,
	axi_full_argRoute_0_w_bits_data,
	axi_full_argRoute_0_w_bits_strb,
	axi_full_argRoute_0_w_bits_last,
	axi_full_argRoute_0_b_ready,
	axi_full_argRoute_0_b_valid,
	axi_full_argRoute_0_b_bits_id,
	axi_full_argRoute_0_b_bits_resp
);
	input clock;
	input reset;
	output wire io_export_argIn_0_TREADY;
	input io_export_argIn_0_TVALID;
	input [63:0] io_export_argIn_0_TDATA;
	output wire io_export_argIn_1_TREADY;
	input io_export_argIn_1_TVALID;
	input [63:0] io_export_argIn_1_TDATA;
	output wire io_export_argIn_2_TREADY;
	input io_export_argIn_2_TVALID;
	input [63:0] io_export_argIn_2_TDATA;
	output wire io_export_argIn_3_TREADY;
	input io_export_argIn_3_TVALID;
	input [63:0] io_export_argIn_3_TDATA;
	output wire io_export_argIn_4_TREADY;
	input io_export_argIn_4_TVALID;
	input [63:0] io_export_argIn_4_TDATA;
	output wire io_export_argIn_5_TREADY;
	input io_export_argIn_5_TVALID;
	input [63:0] io_export_argIn_5_TDATA;
	output wire io_export_argIn_6_TREADY;
	input io_export_argIn_6_TVALID;
	input [63:0] io_export_argIn_6_TDATA;
	output wire io_export_argIn_7_TREADY;
	input io_export_argIn_7_TVALID;
	input [63:0] io_export_argIn_7_TDATA;
	output wire io_export_argIn_8_TREADY;
	input io_export_argIn_8_TVALID;
	input [63:0] io_export_argIn_8_TDATA;
	output wire io_export_argIn_9_TREADY;
	input io_export_argIn_9_TVALID;
	input [63:0] io_export_argIn_9_TDATA;
	output wire io_export_argIn_10_TREADY;
	input io_export_argIn_10_TVALID;
	input [63:0] io_export_argIn_10_TDATA;
	output wire io_export_argIn_11_TREADY;
	input io_export_argIn_11_TVALID;
	input [63:0] io_export_argIn_11_TDATA;
	output wire io_export_argIn_12_TREADY;
	input io_export_argIn_12_TVALID;
	input [63:0] io_export_argIn_12_TDATA;
	output wire io_export_argIn_13_TREADY;
	input io_export_argIn_13_TVALID;
	input [63:0] io_export_argIn_13_TDATA;
	output wire io_export_argIn_14_TREADY;
	input io_export_argIn_14_TVALID;
	input [63:0] io_export_argIn_14_TDATA;
	output wire io_export_argIn_15_TREADY;
	input io_export_argIn_15_TVALID;
	input [63:0] io_export_argIn_15_TDATA;
	output wire io_export_argIn_16_TREADY;
	input io_export_argIn_16_TVALID;
	input [63:0] io_export_argIn_16_TDATA;
	output wire io_export_argIn_17_TREADY;
	input io_export_argIn_17_TVALID;
	input [63:0] io_export_argIn_17_TDATA;
	output wire io_export_argIn_18_TREADY;
	input io_export_argIn_18_TVALID;
	input [63:0] io_export_argIn_18_TDATA;
	output wire io_export_argIn_19_TREADY;
	input io_export_argIn_19_TVALID;
	input [63:0] io_export_argIn_19_TDATA;
	output wire io_export_argIn_20_TREADY;
	input io_export_argIn_20_TVALID;
	input [63:0] io_export_argIn_20_TDATA;
	output wire io_export_argIn_21_TREADY;
	input io_export_argIn_21_TVALID;
	input [63:0] io_export_argIn_21_TDATA;
	output wire io_export_argIn_22_TREADY;
	input io_export_argIn_22_TVALID;
	input [63:0] io_export_argIn_22_TDATA;
	output wire io_export_argIn_23_TREADY;
	input io_export_argIn_23_TVALID;
	input [63:0] io_export_argIn_23_TDATA;
	output wire io_export_argIn_24_TREADY;
	input io_export_argIn_24_TVALID;
	input [63:0] io_export_argIn_24_TDATA;
	output wire io_export_argIn_25_TREADY;
	input io_export_argIn_25_TVALID;
	input [63:0] io_export_argIn_25_TDATA;
	output wire io_export_argIn_26_TREADY;
	input io_export_argIn_26_TVALID;
	input [63:0] io_export_argIn_26_TDATA;
	output wire io_export_argIn_27_TREADY;
	input io_export_argIn_27_TVALID;
	input [63:0] io_export_argIn_27_TDATA;
	output wire io_export_argIn_28_TREADY;
	input io_export_argIn_28_TVALID;
	input [63:0] io_export_argIn_28_TDATA;
	output wire io_export_argIn_29_TREADY;
	input io_export_argIn_29_TVALID;
	input [63:0] io_export_argIn_29_TDATA;
	output wire io_export_argIn_30_TREADY;
	input io_export_argIn_30_TVALID;
	input [63:0] io_export_argIn_30_TDATA;
	output wire io_export_argIn_31_TREADY;
	input io_export_argIn_31_TVALID;
	input [63:0] io_export_argIn_31_TDATA;
	output wire io_export_argIn_32_TREADY;
	input io_export_argIn_32_TVALID;
	input [63:0] io_export_argIn_32_TDATA;
	output wire io_export_argIn_33_TREADY;
	input io_export_argIn_33_TVALID;
	input [63:0] io_export_argIn_33_TDATA;
	output wire io_export_argIn_34_TREADY;
	input io_export_argIn_34_TVALID;
	input [63:0] io_export_argIn_34_TDATA;
	output wire io_export_argIn_35_TREADY;
	input io_export_argIn_35_TVALID;
	input [63:0] io_export_argIn_35_TDATA;
	output wire io_export_argIn_36_TREADY;
	input io_export_argIn_36_TVALID;
	input [63:0] io_export_argIn_36_TDATA;
	output wire io_export_argIn_37_TREADY;
	input io_export_argIn_37_TVALID;
	input [63:0] io_export_argIn_37_TDATA;
	output wire io_export_argIn_38_TREADY;
	input io_export_argIn_38_TVALID;
	input [63:0] io_export_argIn_38_TDATA;
	output wire io_export_argIn_39_TREADY;
	input io_export_argIn_39_TVALID;
	input [63:0] io_export_argIn_39_TDATA;
	output wire io_export_argIn_40_TREADY;
	input io_export_argIn_40_TVALID;
	input [63:0] io_export_argIn_40_TDATA;
	output wire io_export_argIn_41_TREADY;
	input io_export_argIn_41_TVALID;
	input [63:0] io_export_argIn_41_TDATA;
	output wire io_export_argIn_42_TREADY;
	input io_export_argIn_42_TVALID;
	input [63:0] io_export_argIn_42_TDATA;
	output wire io_export_argIn_43_TREADY;
	input io_export_argIn_43_TVALID;
	input [63:0] io_export_argIn_43_TDATA;
	output wire io_export_argIn_44_TREADY;
	input io_export_argIn_44_TVALID;
	input [63:0] io_export_argIn_44_TDATA;
	output wire io_export_argIn_45_TREADY;
	input io_export_argIn_45_TVALID;
	input [63:0] io_export_argIn_45_TDATA;
	output wire io_export_argIn_46_TREADY;
	input io_export_argIn_46_TVALID;
	input [63:0] io_export_argIn_46_TDATA;
	output wire io_export_argIn_47_TREADY;
	input io_export_argIn_47_TVALID;
	input [63:0] io_export_argIn_47_TDATA;
	output wire io_export_argIn_48_TREADY;
	input io_export_argIn_48_TVALID;
	input [63:0] io_export_argIn_48_TDATA;
	output wire io_export_argIn_49_TREADY;
	input io_export_argIn_49_TVALID;
	input [63:0] io_export_argIn_49_TDATA;
	output wire io_export_argIn_50_TREADY;
	input io_export_argIn_50_TVALID;
	input [63:0] io_export_argIn_50_TDATA;
	output wire io_export_argIn_51_TREADY;
	input io_export_argIn_51_TVALID;
	input [63:0] io_export_argIn_51_TDATA;
	output wire io_export_argIn_52_TREADY;
	input io_export_argIn_52_TVALID;
	input [63:0] io_export_argIn_52_TDATA;
	output wire io_export_argIn_53_TREADY;
	input io_export_argIn_53_TVALID;
	input [63:0] io_export_argIn_53_TDATA;
	output wire io_export_argIn_54_TREADY;
	input io_export_argIn_54_TVALID;
	input [63:0] io_export_argIn_54_TDATA;
	output wire io_export_argIn_55_TREADY;
	input io_export_argIn_55_TVALID;
	input [63:0] io_export_argIn_55_TDATA;
	output wire io_export_argIn_56_TREADY;
	input io_export_argIn_56_TVALID;
	input [63:0] io_export_argIn_56_TDATA;
	output wire io_export_argIn_57_TREADY;
	input io_export_argIn_57_TVALID;
	input [63:0] io_export_argIn_57_TDATA;
	output wire io_export_argIn_58_TREADY;
	input io_export_argIn_58_TVALID;
	input [63:0] io_export_argIn_58_TDATA;
	output wire io_export_argIn_59_TREADY;
	input io_export_argIn_59_TVALID;
	input [63:0] io_export_argIn_59_TDATA;
	output wire io_export_argIn_60_TREADY;
	input io_export_argIn_60_TVALID;
	input [63:0] io_export_argIn_60_TDATA;
	output wire io_export_argIn_61_TREADY;
	input io_export_argIn_61_TVALID;
	input [63:0] io_export_argIn_61_TDATA;
	output wire io_export_argIn_62_TREADY;
	input io_export_argIn_62_TVALID;
	input [63:0] io_export_argIn_62_TDATA;
	output wire io_export_argIn_63_TREADY;
	input io_export_argIn_63_TVALID;
	input [63:0] io_export_argIn_63_TDATA;
	output wire io_export_argIn_64_TREADY;
	input io_export_argIn_64_TVALID;
	input [63:0] io_export_argIn_64_TDATA;
	output wire io_export_argIn_65_TREADY;
	input io_export_argIn_65_TVALID;
	input [63:0] io_export_argIn_65_TDATA;
	output wire io_export_argIn_66_TREADY;
	input io_export_argIn_66_TVALID;
	input [63:0] io_export_argIn_66_TDATA;
	output wire io_export_argIn_67_TREADY;
	input io_export_argIn_67_TVALID;
	input [63:0] io_export_argIn_67_TDATA;
	output wire io_export_argIn_68_TREADY;
	input io_export_argIn_68_TVALID;
	input [63:0] io_export_argIn_68_TDATA;
	output wire io_export_argIn_69_TREADY;
	input io_export_argIn_69_TVALID;
	input [63:0] io_export_argIn_69_TDATA;
	output wire io_export_argIn_70_TREADY;
	input io_export_argIn_70_TVALID;
	input [63:0] io_export_argIn_70_TDATA;
	output wire io_export_argIn_71_TREADY;
	input io_export_argIn_71_TVALID;
	input [63:0] io_export_argIn_71_TDATA;
	output wire io_export_argIn_72_TREADY;
	input io_export_argIn_72_TVALID;
	input [63:0] io_export_argIn_72_TDATA;
	output wire io_export_argIn_73_TREADY;
	input io_export_argIn_73_TVALID;
	input [63:0] io_export_argIn_73_TDATA;
	output wire io_export_argIn_74_TREADY;
	input io_export_argIn_74_TVALID;
	input [63:0] io_export_argIn_74_TDATA;
	output wire io_export_argIn_75_TREADY;
	input io_export_argIn_75_TVALID;
	input [63:0] io_export_argIn_75_TDATA;
	output wire io_export_argIn_76_TREADY;
	input io_export_argIn_76_TVALID;
	input [63:0] io_export_argIn_76_TDATA;
	output wire io_export_argIn_77_TREADY;
	input io_export_argIn_77_TVALID;
	input [63:0] io_export_argIn_77_TDATA;
	output wire io_export_argIn_78_TREADY;
	input io_export_argIn_78_TVALID;
	input [63:0] io_export_argIn_78_TDATA;
	output wire io_export_argIn_79_TREADY;
	input io_export_argIn_79_TVALID;
	input [63:0] io_export_argIn_79_TDATA;
	output wire io_export_argIn_80_TREADY;
	input io_export_argIn_80_TVALID;
	input [63:0] io_export_argIn_80_TDATA;
	output wire io_export_argIn_81_TREADY;
	input io_export_argIn_81_TVALID;
	input [63:0] io_export_argIn_81_TDATA;
	output wire io_export_argIn_82_TREADY;
	input io_export_argIn_82_TVALID;
	input [63:0] io_export_argIn_82_TDATA;
	output wire io_export_argIn_83_TREADY;
	input io_export_argIn_83_TVALID;
	input [63:0] io_export_argIn_83_TDATA;
	output wire io_export_argIn_84_TREADY;
	input io_export_argIn_84_TVALID;
	input [63:0] io_export_argIn_84_TDATA;
	output wire io_export_argIn_85_TREADY;
	input io_export_argIn_85_TVALID;
	input [63:0] io_export_argIn_85_TDATA;
	output wire io_export_argIn_86_TREADY;
	input io_export_argIn_86_TVALID;
	input [63:0] io_export_argIn_86_TDATA;
	output wire io_export_argIn_87_TREADY;
	input io_export_argIn_87_TVALID;
	input [63:0] io_export_argIn_87_TDATA;
	output wire io_export_argIn_88_TREADY;
	input io_export_argIn_88_TVALID;
	input [63:0] io_export_argIn_88_TDATA;
	output wire io_export_argIn_89_TREADY;
	input io_export_argIn_89_TVALID;
	input [63:0] io_export_argIn_89_TDATA;
	output wire io_export_argIn_90_TREADY;
	input io_export_argIn_90_TVALID;
	input [63:0] io_export_argIn_90_TDATA;
	output wire io_export_argIn_91_TREADY;
	input io_export_argIn_91_TVALID;
	input [63:0] io_export_argIn_91_TDATA;
	output wire io_export_argIn_92_TREADY;
	input io_export_argIn_92_TVALID;
	input [63:0] io_export_argIn_92_TDATA;
	output wire io_export_argIn_93_TREADY;
	input io_export_argIn_93_TVALID;
	input [63:0] io_export_argIn_93_TDATA;
	output wire io_export_argIn_94_TREADY;
	input io_export_argIn_94_TVALID;
	input [63:0] io_export_argIn_94_TDATA;
	output wire io_export_argIn_95_TREADY;
	input io_export_argIn_95_TVALID;
	input [63:0] io_export_argIn_95_TDATA;
	output wire io_export_argIn_96_TREADY;
	input io_export_argIn_96_TVALID;
	input [63:0] io_export_argIn_96_TDATA;
	output wire io_export_argIn_97_TREADY;
	input io_export_argIn_97_TVALID;
	input [63:0] io_export_argIn_97_TDATA;
	output wire io_export_argIn_98_TREADY;
	input io_export_argIn_98_TVALID;
	input [63:0] io_export_argIn_98_TDATA;
	output wire io_export_argIn_99_TREADY;
	input io_export_argIn_99_TVALID;
	input [63:0] io_export_argIn_99_TDATA;
	output wire io_export_argIn_100_TREADY;
	input io_export_argIn_100_TVALID;
	input [63:0] io_export_argIn_100_TDATA;
	output wire io_export_argIn_101_TREADY;
	input io_export_argIn_101_TVALID;
	input [63:0] io_export_argIn_101_TDATA;
	output wire io_export_argIn_102_TREADY;
	input io_export_argIn_102_TVALID;
	input [63:0] io_export_argIn_102_TDATA;
	output wire io_export_argIn_103_TREADY;
	input io_export_argIn_103_TVALID;
	input [63:0] io_export_argIn_103_TDATA;
	output wire io_export_argIn_104_TREADY;
	input io_export_argIn_104_TVALID;
	input [63:0] io_export_argIn_104_TDATA;
	output wire io_export_argIn_105_TREADY;
	input io_export_argIn_105_TVALID;
	input [63:0] io_export_argIn_105_TDATA;
	output wire io_export_argIn_106_TREADY;
	input io_export_argIn_106_TVALID;
	input [63:0] io_export_argIn_106_TDATA;
	output wire io_export_argIn_107_TREADY;
	input io_export_argIn_107_TVALID;
	input [63:0] io_export_argIn_107_TDATA;
	output wire io_export_argIn_108_TREADY;
	input io_export_argIn_108_TVALID;
	input [63:0] io_export_argIn_108_TDATA;
	output wire io_export_argIn_109_TREADY;
	input io_export_argIn_109_TVALID;
	input [63:0] io_export_argIn_109_TDATA;
	output wire io_export_argIn_110_TREADY;
	input io_export_argIn_110_TVALID;
	input [63:0] io_export_argIn_110_TDATA;
	output wire io_export_argIn_111_TREADY;
	input io_export_argIn_111_TVALID;
	input [63:0] io_export_argIn_111_TDATA;
	output wire io_export_argIn_112_TREADY;
	input io_export_argIn_112_TVALID;
	input [63:0] io_export_argIn_112_TDATA;
	output wire io_export_argIn_113_TREADY;
	input io_export_argIn_113_TVALID;
	input [63:0] io_export_argIn_113_TDATA;
	output wire io_export_argIn_114_TREADY;
	input io_export_argIn_114_TVALID;
	input [63:0] io_export_argIn_114_TDATA;
	output wire io_export_argIn_115_TREADY;
	input io_export_argIn_115_TVALID;
	input [63:0] io_export_argIn_115_TDATA;
	output wire io_export_argIn_116_TREADY;
	input io_export_argIn_116_TVALID;
	input [63:0] io_export_argIn_116_TDATA;
	output wire io_export_argIn_117_TREADY;
	input io_export_argIn_117_TVALID;
	input [63:0] io_export_argIn_117_TDATA;
	output wire io_export_argIn_118_TREADY;
	input io_export_argIn_118_TVALID;
	input [63:0] io_export_argIn_118_TDATA;
	output wire io_export_argIn_119_TREADY;
	input io_export_argIn_119_TVALID;
	input [63:0] io_export_argIn_119_TDATA;
	output wire io_export_argIn_120_TREADY;
	input io_export_argIn_120_TVALID;
	input [63:0] io_export_argIn_120_TDATA;
	output wire io_export_argIn_121_TREADY;
	input io_export_argIn_121_TVALID;
	input [63:0] io_export_argIn_121_TDATA;
	output wire io_export_argIn_122_TREADY;
	input io_export_argIn_122_TVALID;
	input [63:0] io_export_argIn_122_TDATA;
	output wire io_export_argIn_123_TREADY;
	input io_export_argIn_123_TVALID;
	input [63:0] io_export_argIn_123_TDATA;
	output wire io_export_argIn_124_TREADY;
	input io_export_argIn_124_TVALID;
	input [63:0] io_export_argIn_124_TDATA;
	output wire io_export_argIn_125_TREADY;
	input io_export_argIn_125_TVALID;
	input [63:0] io_export_argIn_125_TDATA;
	output wire io_export_argIn_126_TREADY;
	input io_export_argIn_126_TVALID;
	input [63:0] io_export_argIn_126_TDATA;
	output wire io_export_argIn_127_TREADY;
	input io_export_argIn_127_TVALID;
	input [63:0] io_export_argIn_127_TDATA;
	output wire connStealNtw_0_ctrl_serveStealReq_valid;
	input connStealNtw_0_ctrl_serveStealReq_ready;
	input connStealNtw_0_data_qOutTask_ready;
	output wire connStealNtw_0_data_qOutTask_valid;
	output wire [255:0] connStealNtw_0_data_qOutTask_bits;
	output wire connStealNtw_1_ctrl_serveStealReq_valid;
	input connStealNtw_1_ctrl_serveStealReq_ready;
	input connStealNtw_1_data_qOutTask_ready;
	output wire connStealNtw_1_data_qOutTask_valid;
	output wire [255:0] connStealNtw_1_data_qOutTask_bits;
	output wire connStealNtw_2_ctrl_serveStealReq_valid;
	input connStealNtw_2_ctrl_serveStealReq_ready;
	input connStealNtw_2_data_qOutTask_ready;
	output wire connStealNtw_2_data_qOutTask_valid;
	output wire [255:0] connStealNtw_2_data_qOutTask_bits;
	output wire connStealNtw_3_ctrl_serveStealReq_valid;
	input connStealNtw_3_ctrl_serveStealReq_ready;
	input connStealNtw_3_data_qOutTask_ready;
	output wire connStealNtw_3_data_qOutTask_valid;
	output wire [255:0] connStealNtw_3_data_qOutTask_bits;
	output wire connStealNtw_4_ctrl_serveStealReq_valid;
	input connStealNtw_4_ctrl_serveStealReq_ready;
	input connStealNtw_4_data_qOutTask_ready;
	output wire connStealNtw_4_data_qOutTask_valid;
	output wire [255:0] connStealNtw_4_data_qOutTask_bits;
	output wire connStealNtw_5_ctrl_serveStealReq_valid;
	input connStealNtw_5_ctrl_serveStealReq_ready;
	input connStealNtw_5_data_qOutTask_ready;
	output wire connStealNtw_5_data_qOutTask_valid;
	output wire [255:0] connStealNtw_5_data_qOutTask_bits;
	output wire connStealNtw_6_ctrl_serveStealReq_valid;
	input connStealNtw_6_ctrl_serveStealReq_ready;
	input connStealNtw_6_data_qOutTask_ready;
	output wire connStealNtw_6_data_qOutTask_valid;
	output wire [255:0] connStealNtw_6_data_qOutTask_bits;
	output wire connStealNtw_7_ctrl_serveStealReq_valid;
	input connStealNtw_7_ctrl_serveStealReq_ready;
	input connStealNtw_7_data_qOutTask_ready;
	output wire connStealNtw_7_data_qOutTask_valid;
	output wire [255:0] connStealNtw_7_data_qOutTask_bits;
	output wire connStealNtw_8_ctrl_serveStealReq_valid;
	input connStealNtw_8_ctrl_serveStealReq_ready;
	input connStealNtw_8_data_qOutTask_ready;
	output wire connStealNtw_8_data_qOutTask_valid;
	output wire [255:0] connStealNtw_8_data_qOutTask_bits;
	output wire connStealNtw_9_ctrl_serveStealReq_valid;
	input connStealNtw_9_ctrl_serveStealReq_ready;
	input connStealNtw_9_data_qOutTask_ready;
	output wire connStealNtw_9_data_qOutTask_valid;
	output wire [255:0] connStealNtw_9_data_qOutTask_bits;
	output wire connStealNtw_10_ctrl_serveStealReq_valid;
	input connStealNtw_10_ctrl_serveStealReq_ready;
	input connStealNtw_10_data_qOutTask_ready;
	output wire connStealNtw_10_data_qOutTask_valid;
	output wire [255:0] connStealNtw_10_data_qOutTask_bits;
	output wire connStealNtw_11_ctrl_serveStealReq_valid;
	input connStealNtw_11_ctrl_serveStealReq_ready;
	input connStealNtw_11_data_qOutTask_ready;
	output wire connStealNtw_11_data_qOutTask_valid;
	output wire [255:0] connStealNtw_11_data_qOutTask_bits;
	output wire connStealNtw_12_ctrl_serveStealReq_valid;
	input connStealNtw_12_ctrl_serveStealReq_ready;
	input connStealNtw_12_data_qOutTask_ready;
	output wire connStealNtw_12_data_qOutTask_valid;
	output wire [255:0] connStealNtw_12_data_qOutTask_bits;
	output wire connStealNtw_13_ctrl_serveStealReq_valid;
	input connStealNtw_13_ctrl_serveStealReq_ready;
	input connStealNtw_13_data_qOutTask_ready;
	output wire connStealNtw_13_data_qOutTask_valid;
	output wire [255:0] connStealNtw_13_data_qOutTask_bits;
	output wire connStealNtw_14_ctrl_serveStealReq_valid;
	input connStealNtw_14_ctrl_serveStealReq_ready;
	input connStealNtw_14_data_qOutTask_ready;
	output wire connStealNtw_14_data_qOutTask_valid;
	output wire [255:0] connStealNtw_14_data_qOutTask_bits;
	output wire connStealNtw_15_ctrl_serveStealReq_valid;
	input connStealNtw_15_ctrl_serveStealReq_ready;
	input connStealNtw_15_data_qOutTask_ready;
	output wire connStealNtw_15_data_qOutTask_valid;
	output wire [255:0] connStealNtw_15_data_qOutTask_bits;
	input axi_full_argRoute_0_ar_ready;
	output wire axi_full_argRoute_0_ar_valid;
	output wire [4:0] axi_full_argRoute_0_ar_bits_id;
	output wire [63:0] axi_full_argRoute_0_ar_bits_addr;
	output wire [7:0] axi_full_argRoute_0_ar_bits_len;
	output wire [2:0] axi_full_argRoute_0_ar_bits_size;
	output wire [1:0] axi_full_argRoute_0_ar_bits_burst;
	output wire axi_full_argRoute_0_ar_bits_lock;
	output wire [3:0] axi_full_argRoute_0_ar_bits_cache;
	output wire [2:0] axi_full_argRoute_0_ar_bits_prot;
	output wire [3:0] axi_full_argRoute_0_ar_bits_qos;
	output wire [3:0] axi_full_argRoute_0_ar_bits_region;
	output wire axi_full_argRoute_0_r_ready;
	input axi_full_argRoute_0_r_valid;
	input [4:0] axi_full_argRoute_0_r_bits_id;
	input [31:0] axi_full_argRoute_0_r_bits_data;
	input [1:0] axi_full_argRoute_0_r_bits_resp;
	input axi_full_argRoute_0_r_bits_last;
	input axi_full_argRoute_0_aw_ready;
	output wire axi_full_argRoute_0_aw_valid;
	output wire [4:0] axi_full_argRoute_0_aw_bits_id;
	output wire [63:0] axi_full_argRoute_0_aw_bits_addr;
	output wire [7:0] axi_full_argRoute_0_aw_bits_len;
	output wire [2:0] axi_full_argRoute_0_aw_bits_size;
	output wire [1:0] axi_full_argRoute_0_aw_bits_burst;
	output wire axi_full_argRoute_0_aw_bits_lock;
	output wire [3:0] axi_full_argRoute_0_aw_bits_cache;
	output wire [2:0] axi_full_argRoute_0_aw_bits_prot;
	output wire [3:0] axi_full_argRoute_0_aw_bits_qos;
	output wire [3:0] axi_full_argRoute_0_aw_bits_region;
	input axi_full_argRoute_0_w_ready;
	output wire axi_full_argRoute_0_w_valid;
	output wire [31:0] axi_full_argRoute_0_w_bits_data;
	output wire [3:0] axi_full_argRoute_0_w_bits_strb;
	output wire axi_full_argRoute_0_w_bits_last;
	output wire axi_full_argRoute_0_b_ready;
	input axi_full_argRoute_0_b_valid;
	input [4:0] axi_full_argRoute_0_b_bits_id;
	input [1:0] axi_full_argRoute_0_b_bits_resp;
	wire _axis_stream_converters_in_127_io_dataIn_TREADY;
	wire _axis_stream_converters_in_127_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_127_io_dataOut_TDATA;
	wire _axis_stream_converters_in_126_io_dataIn_TREADY;
	wire _axis_stream_converters_in_126_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_126_io_dataOut_TDATA;
	wire _axis_stream_converters_in_125_io_dataIn_TREADY;
	wire _axis_stream_converters_in_125_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_125_io_dataOut_TDATA;
	wire _axis_stream_converters_in_124_io_dataIn_TREADY;
	wire _axis_stream_converters_in_124_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_124_io_dataOut_TDATA;
	wire _axis_stream_converters_in_123_io_dataIn_TREADY;
	wire _axis_stream_converters_in_123_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_123_io_dataOut_TDATA;
	wire _axis_stream_converters_in_122_io_dataIn_TREADY;
	wire _axis_stream_converters_in_122_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_122_io_dataOut_TDATA;
	wire _axis_stream_converters_in_121_io_dataIn_TREADY;
	wire _axis_stream_converters_in_121_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_121_io_dataOut_TDATA;
	wire _axis_stream_converters_in_120_io_dataIn_TREADY;
	wire _axis_stream_converters_in_120_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_120_io_dataOut_TDATA;
	wire _axis_stream_converters_in_119_io_dataIn_TREADY;
	wire _axis_stream_converters_in_119_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_119_io_dataOut_TDATA;
	wire _axis_stream_converters_in_118_io_dataIn_TREADY;
	wire _axis_stream_converters_in_118_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_118_io_dataOut_TDATA;
	wire _axis_stream_converters_in_117_io_dataIn_TREADY;
	wire _axis_stream_converters_in_117_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_117_io_dataOut_TDATA;
	wire _axis_stream_converters_in_116_io_dataIn_TREADY;
	wire _axis_stream_converters_in_116_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_116_io_dataOut_TDATA;
	wire _axis_stream_converters_in_115_io_dataIn_TREADY;
	wire _axis_stream_converters_in_115_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_115_io_dataOut_TDATA;
	wire _axis_stream_converters_in_114_io_dataIn_TREADY;
	wire _axis_stream_converters_in_114_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_114_io_dataOut_TDATA;
	wire _axis_stream_converters_in_113_io_dataIn_TREADY;
	wire _axis_stream_converters_in_113_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_113_io_dataOut_TDATA;
	wire _axis_stream_converters_in_112_io_dataIn_TREADY;
	wire _axis_stream_converters_in_112_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_112_io_dataOut_TDATA;
	wire _axis_stream_converters_in_111_io_dataIn_TREADY;
	wire _axis_stream_converters_in_111_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_111_io_dataOut_TDATA;
	wire _axis_stream_converters_in_110_io_dataIn_TREADY;
	wire _axis_stream_converters_in_110_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_110_io_dataOut_TDATA;
	wire _axis_stream_converters_in_109_io_dataIn_TREADY;
	wire _axis_stream_converters_in_109_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_109_io_dataOut_TDATA;
	wire _axis_stream_converters_in_108_io_dataIn_TREADY;
	wire _axis_stream_converters_in_108_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_108_io_dataOut_TDATA;
	wire _axis_stream_converters_in_107_io_dataIn_TREADY;
	wire _axis_stream_converters_in_107_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_107_io_dataOut_TDATA;
	wire _axis_stream_converters_in_106_io_dataIn_TREADY;
	wire _axis_stream_converters_in_106_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_106_io_dataOut_TDATA;
	wire _axis_stream_converters_in_105_io_dataIn_TREADY;
	wire _axis_stream_converters_in_105_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_105_io_dataOut_TDATA;
	wire _axis_stream_converters_in_104_io_dataIn_TREADY;
	wire _axis_stream_converters_in_104_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_104_io_dataOut_TDATA;
	wire _axis_stream_converters_in_103_io_dataIn_TREADY;
	wire _axis_stream_converters_in_103_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_103_io_dataOut_TDATA;
	wire _axis_stream_converters_in_102_io_dataIn_TREADY;
	wire _axis_stream_converters_in_102_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_102_io_dataOut_TDATA;
	wire _axis_stream_converters_in_101_io_dataIn_TREADY;
	wire _axis_stream_converters_in_101_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_101_io_dataOut_TDATA;
	wire _axis_stream_converters_in_100_io_dataIn_TREADY;
	wire _axis_stream_converters_in_100_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_100_io_dataOut_TDATA;
	wire _axis_stream_converters_in_99_io_dataIn_TREADY;
	wire _axis_stream_converters_in_99_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_99_io_dataOut_TDATA;
	wire _axis_stream_converters_in_98_io_dataIn_TREADY;
	wire _axis_stream_converters_in_98_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_98_io_dataOut_TDATA;
	wire _axis_stream_converters_in_97_io_dataIn_TREADY;
	wire _axis_stream_converters_in_97_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_97_io_dataOut_TDATA;
	wire _axis_stream_converters_in_96_io_dataIn_TREADY;
	wire _axis_stream_converters_in_96_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_96_io_dataOut_TDATA;
	wire _axis_stream_converters_in_95_io_dataIn_TREADY;
	wire _axis_stream_converters_in_95_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_95_io_dataOut_TDATA;
	wire _axis_stream_converters_in_94_io_dataIn_TREADY;
	wire _axis_stream_converters_in_94_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_94_io_dataOut_TDATA;
	wire _axis_stream_converters_in_93_io_dataIn_TREADY;
	wire _axis_stream_converters_in_93_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_93_io_dataOut_TDATA;
	wire _axis_stream_converters_in_92_io_dataIn_TREADY;
	wire _axis_stream_converters_in_92_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_92_io_dataOut_TDATA;
	wire _axis_stream_converters_in_91_io_dataIn_TREADY;
	wire _axis_stream_converters_in_91_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_91_io_dataOut_TDATA;
	wire _axis_stream_converters_in_90_io_dataIn_TREADY;
	wire _axis_stream_converters_in_90_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_90_io_dataOut_TDATA;
	wire _axis_stream_converters_in_89_io_dataIn_TREADY;
	wire _axis_stream_converters_in_89_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_89_io_dataOut_TDATA;
	wire _axis_stream_converters_in_88_io_dataIn_TREADY;
	wire _axis_stream_converters_in_88_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_88_io_dataOut_TDATA;
	wire _axis_stream_converters_in_87_io_dataIn_TREADY;
	wire _axis_stream_converters_in_87_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_87_io_dataOut_TDATA;
	wire _axis_stream_converters_in_86_io_dataIn_TREADY;
	wire _axis_stream_converters_in_86_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_86_io_dataOut_TDATA;
	wire _axis_stream_converters_in_85_io_dataIn_TREADY;
	wire _axis_stream_converters_in_85_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_85_io_dataOut_TDATA;
	wire _axis_stream_converters_in_84_io_dataIn_TREADY;
	wire _axis_stream_converters_in_84_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_84_io_dataOut_TDATA;
	wire _axis_stream_converters_in_83_io_dataIn_TREADY;
	wire _axis_stream_converters_in_83_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_83_io_dataOut_TDATA;
	wire _axis_stream_converters_in_82_io_dataIn_TREADY;
	wire _axis_stream_converters_in_82_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_82_io_dataOut_TDATA;
	wire _axis_stream_converters_in_81_io_dataIn_TREADY;
	wire _axis_stream_converters_in_81_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_81_io_dataOut_TDATA;
	wire _axis_stream_converters_in_80_io_dataIn_TREADY;
	wire _axis_stream_converters_in_80_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_80_io_dataOut_TDATA;
	wire _axis_stream_converters_in_79_io_dataIn_TREADY;
	wire _axis_stream_converters_in_79_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_79_io_dataOut_TDATA;
	wire _axis_stream_converters_in_78_io_dataIn_TREADY;
	wire _axis_stream_converters_in_78_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_78_io_dataOut_TDATA;
	wire _axis_stream_converters_in_77_io_dataIn_TREADY;
	wire _axis_stream_converters_in_77_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_77_io_dataOut_TDATA;
	wire _axis_stream_converters_in_76_io_dataIn_TREADY;
	wire _axis_stream_converters_in_76_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_76_io_dataOut_TDATA;
	wire _axis_stream_converters_in_75_io_dataIn_TREADY;
	wire _axis_stream_converters_in_75_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_75_io_dataOut_TDATA;
	wire _axis_stream_converters_in_74_io_dataIn_TREADY;
	wire _axis_stream_converters_in_74_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_74_io_dataOut_TDATA;
	wire _axis_stream_converters_in_73_io_dataIn_TREADY;
	wire _axis_stream_converters_in_73_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_73_io_dataOut_TDATA;
	wire _axis_stream_converters_in_72_io_dataIn_TREADY;
	wire _axis_stream_converters_in_72_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_72_io_dataOut_TDATA;
	wire _axis_stream_converters_in_71_io_dataIn_TREADY;
	wire _axis_stream_converters_in_71_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_71_io_dataOut_TDATA;
	wire _axis_stream_converters_in_70_io_dataIn_TREADY;
	wire _axis_stream_converters_in_70_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_70_io_dataOut_TDATA;
	wire _axis_stream_converters_in_69_io_dataIn_TREADY;
	wire _axis_stream_converters_in_69_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_69_io_dataOut_TDATA;
	wire _axis_stream_converters_in_68_io_dataIn_TREADY;
	wire _axis_stream_converters_in_68_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_68_io_dataOut_TDATA;
	wire _axis_stream_converters_in_67_io_dataIn_TREADY;
	wire _axis_stream_converters_in_67_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_67_io_dataOut_TDATA;
	wire _axis_stream_converters_in_66_io_dataIn_TREADY;
	wire _axis_stream_converters_in_66_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_66_io_dataOut_TDATA;
	wire _axis_stream_converters_in_65_io_dataIn_TREADY;
	wire _axis_stream_converters_in_65_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_65_io_dataOut_TDATA;
	wire _axis_stream_converters_in_64_io_dataIn_TREADY;
	wire _axis_stream_converters_in_64_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_64_io_dataOut_TDATA;
	wire _axis_stream_converters_in_63_io_dataIn_TREADY;
	wire _axis_stream_converters_in_63_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_63_io_dataOut_TDATA;
	wire _axis_stream_converters_in_62_io_dataIn_TREADY;
	wire _axis_stream_converters_in_62_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_62_io_dataOut_TDATA;
	wire _axis_stream_converters_in_61_io_dataIn_TREADY;
	wire _axis_stream_converters_in_61_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_61_io_dataOut_TDATA;
	wire _axis_stream_converters_in_60_io_dataIn_TREADY;
	wire _axis_stream_converters_in_60_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_60_io_dataOut_TDATA;
	wire _axis_stream_converters_in_59_io_dataIn_TREADY;
	wire _axis_stream_converters_in_59_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_59_io_dataOut_TDATA;
	wire _axis_stream_converters_in_58_io_dataIn_TREADY;
	wire _axis_stream_converters_in_58_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_58_io_dataOut_TDATA;
	wire _axis_stream_converters_in_57_io_dataIn_TREADY;
	wire _axis_stream_converters_in_57_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_57_io_dataOut_TDATA;
	wire _axis_stream_converters_in_56_io_dataIn_TREADY;
	wire _axis_stream_converters_in_56_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_56_io_dataOut_TDATA;
	wire _axis_stream_converters_in_55_io_dataIn_TREADY;
	wire _axis_stream_converters_in_55_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_55_io_dataOut_TDATA;
	wire _axis_stream_converters_in_54_io_dataIn_TREADY;
	wire _axis_stream_converters_in_54_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_54_io_dataOut_TDATA;
	wire _axis_stream_converters_in_53_io_dataIn_TREADY;
	wire _axis_stream_converters_in_53_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_53_io_dataOut_TDATA;
	wire _axis_stream_converters_in_52_io_dataIn_TREADY;
	wire _axis_stream_converters_in_52_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_52_io_dataOut_TDATA;
	wire _axis_stream_converters_in_51_io_dataIn_TREADY;
	wire _axis_stream_converters_in_51_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_51_io_dataOut_TDATA;
	wire _axis_stream_converters_in_50_io_dataIn_TREADY;
	wire _axis_stream_converters_in_50_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_50_io_dataOut_TDATA;
	wire _axis_stream_converters_in_49_io_dataIn_TREADY;
	wire _axis_stream_converters_in_49_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_49_io_dataOut_TDATA;
	wire _axis_stream_converters_in_48_io_dataIn_TREADY;
	wire _axis_stream_converters_in_48_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_48_io_dataOut_TDATA;
	wire _axis_stream_converters_in_47_io_dataIn_TREADY;
	wire _axis_stream_converters_in_47_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_47_io_dataOut_TDATA;
	wire _axis_stream_converters_in_46_io_dataIn_TREADY;
	wire _axis_stream_converters_in_46_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_46_io_dataOut_TDATA;
	wire _axis_stream_converters_in_45_io_dataIn_TREADY;
	wire _axis_stream_converters_in_45_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_45_io_dataOut_TDATA;
	wire _axis_stream_converters_in_44_io_dataIn_TREADY;
	wire _axis_stream_converters_in_44_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_44_io_dataOut_TDATA;
	wire _axis_stream_converters_in_43_io_dataIn_TREADY;
	wire _axis_stream_converters_in_43_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_43_io_dataOut_TDATA;
	wire _axis_stream_converters_in_42_io_dataIn_TREADY;
	wire _axis_stream_converters_in_42_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_42_io_dataOut_TDATA;
	wire _axis_stream_converters_in_41_io_dataIn_TREADY;
	wire _axis_stream_converters_in_41_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_41_io_dataOut_TDATA;
	wire _axis_stream_converters_in_40_io_dataIn_TREADY;
	wire _axis_stream_converters_in_40_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_40_io_dataOut_TDATA;
	wire _axis_stream_converters_in_39_io_dataIn_TREADY;
	wire _axis_stream_converters_in_39_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_39_io_dataOut_TDATA;
	wire _axis_stream_converters_in_38_io_dataIn_TREADY;
	wire _axis_stream_converters_in_38_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_38_io_dataOut_TDATA;
	wire _axis_stream_converters_in_37_io_dataIn_TREADY;
	wire _axis_stream_converters_in_37_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_37_io_dataOut_TDATA;
	wire _axis_stream_converters_in_36_io_dataIn_TREADY;
	wire _axis_stream_converters_in_36_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_36_io_dataOut_TDATA;
	wire _axis_stream_converters_in_35_io_dataIn_TREADY;
	wire _axis_stream_converters_in_35_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_35_io_dataOut_TDATA;
	wire _axis_stream_converters_in_34_io_dataIn_TREADY;
	wire _axis_stream_converters_in_34_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_34_io_dataOut_TDATA;
	wire _axis_stream_converters_in_33_io_dataIn_TREADY;
	wire _axis_stream_converters_in_33_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_33_io_dataOut_TDATA;
	wire _axis_stream_converters_in_32_io_dataIn_TREADY;
	wire _axis_stream_converters_in_32_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_32_io_dataOut_TDATA;
	wire _axis_stream_converters_in_31_io_dataIn_TREADY;
	wire _axis_stream_converters_in_31_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_31_io_dataOut_TDATA;
	wire _axis_stream_converters_in_30_io_dataIn_TREADY;
	wire _axis_stream_converters_in_30_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_30_io_dataOut_TDATA;
	wire _axis_stream_converters_in_29_io_dataIn_TREADY;
	wire _axis_stream_converters_in_29_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_29_io_dataOut_TDATA;
	wire _axis_stream_converters_in_28_io_dataIn_TREADY;
	wire _axis_stream_converters_in_28_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_28_io_dataOut_TDATA;
	wire _axis_stream_converters_in_27_io_dataIn_TREADY;
	wire _axis_stream_converters_in_27_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_27_io_dataOut_TDATA;
	wire _axis_stream_converters_in_26_io_dataIn_TREADY;
	wire _axis_stream_converters_in_26_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_26_io_dataOut_TDATA;
	wire _axis_stream_converters_in_25_io_dataIn_TREADY;
	wire _axis_stream_converters_in_25_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_25_io_dataOut_TDATA;
	wire _axis_stream_converters_in_24_io_dataIn_TREADY;
	wire _axis_stream_converters_in_24_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_24_io_dataOut_TDATA;
	wire _axis_stream_converters_in_23_io_dataIn_TREADY;
	wire _axis_stream_converters_in_23_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_23_io_dataOut_TDATA;
	wire _axis_stream_converters_in_22_io_dataIn_TREADY;
	wire _axis_stream_converters_in_22_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_22_io_dataOut_TDATA;
	wire _axis_stream_converters_in_21_io_dataIn_TREADY;
	wire _axis_stream_converters_in_21_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_21_io_dataOut_TDATA;
	wire _axis_stream_converters_in_20_io_dataIn_TREADY;
	wire _axis_stream_converters_in_20_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_20_io_dataOut_TDATA;
	wire _axis_stream_converters_in_19_io_dataIn_TREADY;
	wire _axis_stream_converters_in_19_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_19_io_dataOut_TDATA;
	wire _axis_stream_converters_in_18_io_dataIn_TREADY;
	wire _axis_stream_converters_in_18_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_18_io_dataOut_TDATA;
	wire _axis_stream_converters_in_17_io_dataIn_TREADY;
	wire _axis_stream_converters_in_17_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_17_io_dataOut_TDATA;
	wire _axis_stream_converters_in_16_io_dataIn_TREADY;
	wire _axis_stream_converters_in_16_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_16_io_dataOut_TDATA;
	wire _axis_stream_converters_in_15_io_dataIn_TREADY;
	wire _axis_stream_converters_in_15_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_15_io_dataOut_TDATA;
	wire _axis_stream_converters_in_14_io_dataIn_TREADY;
	wire _axis_stream_converters_in_14_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_14_io_dataOut_TDATA;
	wire _axis_stream_converters_in_13_io_dataIn_TREADY;
	wire _axis_stream_converters_in_13_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_13_io_dataOut_TDATA;
	wire _axis_stream_converters_in_12_io_dataIn_TREADY;
	wire _axis_stream_converters_in_12_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_12_io_dataOut_TDATA;
	wire _axis_stream_converters_in_11_io_dataIn_TREADY;
	wire _axis_stream_converters_in_11_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_11_io_dataOut_TDATA;
	wire _axis_stream_converters_in_10_io_dataIn_TREADY;
	wire _axis_stream_converters_in_10_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_10_io_dataOut_TDATA;
	wire _axis_stream_converters_in_9_io_dataIn_TREADY;
	wire _axis_stream_converters_in_9_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_9_io_dataOut_TDATA;
	wire _axis_stream_converters_in_8_io_dataIn_TREADY;
	wire _axis_stream_converters_in_8_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_8_io_dataOut_TDATA;
	wire _axis_stream_converters_in_7_io_dataIn_TREADY;
	wire _axis_stream_converters_in_7_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_7_io_dataOut_TDATA;
	wire _axis_stream_converters_in_6_io_dataIn_TREADY;
	wire _axis_stream_converters_in_6_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_6_io_dataOut_TDATA;
	wire _axis_stream_converters_in_5_io_dataIn_TREADY;
	wire _axis_stream_converters_in_5_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_5_io_dataOut_TDATA;
	wire _axis_stream_converters_in_4_io_dataIn_TREADY;
	wire _axis_stream_converters_in_4_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_4_io_dataOut_TDATA;
	wire _axis_stream_converters_in_3_io_dataIn_TREADY;
	wire _axis_stream_converters_in_3_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_3_io_dataOut_TDATA;
	wire _axis_stream_converters_in_2_io_dataIn_TREADY;
	wire _axis_stream_converters_in_2_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_2_io_dataOut_TDATA;
	wire _axis_stream_converters_in_1_io_dataIn_TREADY;
	wire _axis_stream_converters_in_1_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_1_io_dataOut_TDATA;
	wire _axis_stream_converters_in_0_io_dataIn_TREADY;
	wire _axis_stream_converters_in_0_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_0_io_dataOut_TDATA;
	wire _mux_s_axi_0_ar_ready;
	wire _mux_s_axi_0_r_valid;
	wire [31:0] _mux_s_axi_0_r_bits_data;
	wire _mux_s_axi_0_aw_ready;
	wire _mux_s_axi_0_w_ready;
	wire _mux_s_axi_0_b_valid;
	wire _mux_s_axi_1_ar_ready;
	wire _mux_s_axi_1_r_valid;
	wire [31:0] _mux_s_axi_1_r_bits_data;
	wire _mux_s_axi_1_aw_ready;
	wire _mux_s_axi_1_w_ready;
	wire _mux_s_axi_1_b_valid;
	wire _mux_s_axi_2_ar_ready;
	wire _mux_s_axi_2_r_valid;
	wire [31:0] _mux_s_axi_2_r_bits_data;
	wire _mux_s_axi_2_aw_ready;
	wire _mux_s_axi_2_w_ready;
	wire _mux_s_axi_2_b_valid;
	wire _mux_s_axi_3_ar_ready;
	wire _mux_s_axi_3_r_valid;
	wire [31:0] _mux_s_axi_3_r_bits_data;
	wire _mux_s_axi_3_aw_ready;
	wire _mux_s_axi_3_w_ready;
	wire _mux_s_axi_3_b_valid;
	wire _mux_s_axi_4_ar_ready;
	wire _mux_s_axi_4_r_valid;
	wire [31:0] _mux_s_axi_4_r_bits_data;
	wire _mux_s_axi_4_aw_ready;
	wire _mux_s_axi_4_w_ready;
	wire _mux_s_axi_4_b_valid;
	wire _mux_s_axi_5_ar_ready;
	wire _mux_s_axi_5_r_valid;
	wire [31:0] _mux_s_axi_5_r_bits_data;
	wire _mux_s_axi_5_aw_ready;
	wire _mux_s_axi_5_w_ready;
	wire _mux_s_axi_5_b_valid;
	wire _mux_s_axi_6_ar_ready;
	wire _mux_s_axi_6_r_valid;
	wire [31:0] _mux_s_axi_6_r_bits_data;
	wire _mux_s_axi_6_aw_ready;
	wire _mux_s_axi_6_w_ready;
	wire _mux_s_axi_6_b_valid;
	wire _mux_s_axi_7_ar_ready;
	wire _mux_s_axi_7_r_valid;
	wire [31:0] _mux_s_axi_7_r_bits_data;
	wire _mux_s_axi_7_aw_ready;
	wire _mux_s_axi_7_w_ready;
	wire _mux_s_axi_7_b_valid;
	wire _mux_s_axi_8_ar_ready;
	wire _mux_s_axi_8_r_valid;
	wire [31:0] _mux_s_axi_8_r_bits_data;
	wire _mux_s_axi_8_aw_ready;
	wire _mux_s_axi_8_w_ready;
	wire _mux_s_axi_8_b_valid;
	wire _mux_s_axi_9_ar_ready;
	wire _mux_s_axi_9_r_valid;
	wire [31:0] _mux_s_axi_9_r_bits_data;
	wire _mux_s_axi_9_aw_ready;
	wire _mux_s_axi_9_w_ready;
	wire _mux_s_axi_9_b_valid;
	wire _mux_s_axi_10_ar_ready;
	wire _mux_s_axi_10_r_valid;
	wire [31:0] _mux_s_axi_10_r_bits_data;
	wire _mux_s_axi_10_aw_ready;
	wire _mux_s_axi_10_w_ready;
	wire _mux_s_axi_10_b_valid;
	wire _mux_s_axi_11_ar_ready;
	wire _mux_s_axi_11_r_valid;
	wire [31:0] _mux_s_axi_11_r_bits_data;
	wire _mux_s_axi_11_aw_ready;
	wire _mux_s_axi_11_w_ready;
	wire _mux_s_axi_11_b_valid;
	wire _mux_s_axi_12_ar_ready;
	wire _mux_s_axi_12_r_valid;
	wire [31:0] _mux_s_axi_12_r_bits_data;
	wire _mux_s_axi_12_aw_ready;
	wire _mux_s_axi_12_w_ready;
	wire _mux_s_axi_12_b_valid;
	wire _mux_s_axi_13_ar_ready;
	wire _mux_s_axi_13_r_valid;
	wire [31:0] _mux_s_axi_13_r_bits_data;
	wire _mux_s_axi_13_aw_ready;
	wire _mux_s_axi_13_w_ready;
	wire _mux_s_axi_13_b_valid;
	wire _mux_s_axi_14_ar_ready;
	wire _mux_s_axi_14_r_valid;
	wire [31:0] _mux_s_axi_14_r_bits_data;
	wire _mux_s_axi_14_aw_ready;
	wire _mux_s_axi_14_w_ready;
	wire _mux_s_axi_14_b_valid;
	wire _mux_s_axi_15_ar_ready;
	wire _mux_s_axi_15_r_valid;
	wire [31:0] _mux_s_axi_15_r_bits_data;
	wire _mux_s_axi_15_aw_ready;
	wire _mux_s_axi_15_w_ready;
	wire _mux_s_axi_15_b_valid;
	wire _mux_s_axi_16_ar_ready;
	wire _mux_s_axi_16_r_valid;
	wire [31:0] _mux_s_axi_16_r_bits_data;
	wire _mux_s_axi_17_ar_ready;
	wire _mux_s_axi_17_r_valid;
	wire [31:0] _mux_s_axi_17_r_bits_data;
	wire _mux_s_axi_18_ar_ready;
	wire _mux_s_axi_18_r_valid;
	wire [31:0] _mux_s_axi_18_r_bits_data;
	wire _mux_s_axi_19_ar_ready;
	wire _mux_s_axi_19_r_valid;
	wire [31:0] _mux_s_axi_19_r_bits_data;
	wire _mux_s_axi_20_ar_ready;
	wire _mux_s_axi_20_r_valid;
	wire [31:0] _mux_s_axi_20_r_bits_data;
	wire _mux_s_axi_21_ar_ready;
	wire _mux_s_axi_21_r_valid;
	wire [31:0] _mux_s_axi_21_r_bits_data;
	wire _mux_s_axi_22_ar_ready;
	wire _mux_s_axi_22_r_valid;
	wire [31:0] _mux_s_axi_22_r_bits_data;
	wire _mux_s_axi_23_ar_ready;
	wire _mux_s_axi_23_r_valid;
	wire [31:0] _mux_s_axi_23_r_bits_data;
	wire _mux_s_axi_24_ar_ready;
	wire _mux_s_axi_24_r_valid;
	wire [31:0] _mux_s_axi_24_r_bits_data;
	wire _mux_s_axi_25_ar_ready;
	wire _mux_s_axi_25_r_valid;
	wire [31:0] _mux_s_axi_25_r_bits_data;
	wire _mux_s_axi_26_ar_ready;
	wire _mux_s_axi_26_r_valid;
	wire [31:0] _mux_s_axi_26_r_bits_data;
	wire _mux_s_axi_27_ar_ready;
	wire _mux_s_axi_27_r_valid;
	wire [31:0] _mux_s_axi_27_r_bits_data;
	wire _mux_s_axi_28_ar_ready;
	wire _mux_s_axi_28_r_valid;
	wire [31:0] _mux_s_axi_28_r_bits_data;
	wire _mux_s_axi_29_ar_ready;
	wire _mux_s_axi_29_r_valid;
	wire [31:0] _mux_s_axi_29_r_bits_data;
	wire _mux_s_axi_30_ar_ready;
	wire _mux_s_axi_30_r_valid;
	wire [31:0] _mux_s_axi_30_r_bits_data;
	wire _mux_s_axi_31_ar_ready;
	wire _mux_s_axi_31_r_valid;
	wire [31:0] _mux_s_axi_31_r_bits_data;
	wire _argRouteRvmReadOnly_15_io_read_address_ready;
	wire _argRouteRvmReadOnly_15_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_15_io_read_data_bits;
	wire _argRouteRvmReadOnly_15_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_15_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_15_axi_r_ready;
	wire _argRouteRvmReadOnly_14_io_read_address_ready;
	wire _argRouteRvmReadOnly_14_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_14_io_read_data_bits;
	wire _argRouteRvmReadOnly_14_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_14_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_14_axi_r_ready;
	wire _argRouteRvmReadOnly_13_io_read_address_ready;
	wire _argRouteRvmReadOnly_13_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_13_io_read_data_bits;
	wire _argRouteRvmReadOnly_13_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_13_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_13_axi_r_ready;
	wire _argRouteRvmReadOnly_12_io_read_address_ready;
	wire _argRouteRvmReadOnly_12_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_12_io_read_data_bits;
	wire _argRouteRvmReadOnly_12_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_12_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_12_axi_r_ready;
	wire _argRouteRvmReadOnly_11_io_read_address_ready;
	wire _argRouteRvmReadOnly_11_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_11_io_read_data_bits;
	wire _argRouteRvmReadOnly_11_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_11_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_11_axi_r_ready;
	wire _argRouteRvmReadOnly_10_io_read_address_ready;
	wire _argRouteRvmReadOnly_10_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_10_io_read_data_bits;
	wire _argRouteRvmReadOnly_10_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_10_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_10_axi_r_ready;
	wire _argRouteRvmReadOnly_9_io_read_address_ready;
	wire _argRouteRvmReadOnly_9_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_9_io_read_data_bits;
	wire _argRouteRvmReadOnly_9_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_9_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_9_axi_r_ready;
	wire _argRouteRvmReadOnly_8_io_read_address_ready;
	wire _argRouteRvmReadOnly_8_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_8_io_read_data_bits;
	wire _argRouteRvmReadOnly_8_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_8_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_8_axi_r_ready;
	wire _argRouteRvmReadOnly_7_io_read_address_ready;
	wire _argRouteRvmReadOnly_7_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_7_io_read_data_bits;
	wire _argRouteRvmReadOnly_7_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_7_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_7_axi_r_ready;
	wire _argRouteRvmReadOnly_6_io_read_address_ready;
	wire _argRouteRvmReadOnly_6_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_6_io_read_data_bits;
	wire _argRouteRvmReadOnly_6_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_6_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_6_axi_r_ready;
	wire _argRouteRvmReadOnly_5_io_read_address_ready;
	wire _argRouteRvmReadOnly_5_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_5_io_read_data_bits;
	wire _argRouteRvmReadOnly_5_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_5_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_5_axi_r_ready;
	wire _argRouteRvmReadOnly_4_io_read_address_ready;
	wire _argRouteRvmReadOnly_4_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_4_io_read_data_bits;
	wire _argRouteRvmReadOnly_4_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_4_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_4_axi_r_ready;
	wire _argRouteRvmReadOnly_3_io_read_address_ready;
	wire _argRouteRvmReadOnly_3_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_3_io_read_data_bits;
	wire _argRouteRvmReadOnly_3_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_3_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_3_axi_r_ready;
	wire _argRouteRvmReadOnly_2_io_read_address_ready;
	wire _argRouteRvmReadOnly_2_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_2_io_read_data_bits;
	wire _argRouteRvmReadOnly_2_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_2_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_2_axi_r_ready;
	wire _argRouteRvmReadOnly_1_io_read_address_ready;
	wire _argRouteRvmReadOnly_1_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_1_io_read_data_bits;
	wire _argRouteRvmReadOnly_1_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_1_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_1_axi_r_ready;
	wire _argRouteRvmReadOnly_0_io_read_address_ready;
	wire _argRouteRvmReadOnly_0_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_0_io_read_data_bits;
	wire _argRouteRvmReadOnly_0_axi_ar_valid;
	wire [63:0] _argRouteRvmReadOnly_0_axi_ar_bits_addr;
	wire _argRouteRvmReadOnly_0_axi_r_ready;
	wire _argRouteRvm_15_io_read_address_ready;
	wire _argRouteRvm_15_io_read_data_valid;
	wire [31:0] _argRouteRvm_15_io_read_data_bits;
	wire _argRouteRvm_15_io_write_address_ready;
	wire _argRouteRvm_15_io_write_data_ready;
	wire _argRouteRvm_15_axi_ar_valid;
	wire [63:0] _argRouteRvm_15_axi_ar_bits_addr;
	wire _argRouteRvm_15_axi_r_ready;
	wire _argRouteRvm_15_axi_aw_valid;
	wire [63:0] _argRouteRvm_15_axi_aw_bits_addr;
	wire _argRouteRvm_15_axi_w_valid;
	wire [31:0] _argRouteRvm_15_axi_w_bits_data;
	wire _argRouteRvm_14_io_read_address_ready;
	wire _argRouteRvm_14_io_read_data_valid;
	wire [31:0] _argRouteRvm_14_io_read_data_bits;
	wire _argRouteRvm_14_io_write_address_ready;
	wire _argRouteRvm_14_io_write_data_ready;
	wire _argRouteRvm_14_axi_ar_valid;
	wire [63:0] _argRouteRvm_14_axi_ar_bits_addr;
	wire _argRouteRvm_14_axi_r_ready;
	wire _argRouteRvm_14_axi_aw_valid;
	wire [63:0] _argRouteRvm_14_axi_aw_bits_addr;
	wire _argRouteRvm_14_axi_w_valid;
	wire [31:0] _argRouteRvm_14_axi_w_bits_data;
	wire _argRouteRvm_13_io_read_address_ready;
	wire _argRouteRvm_13_io_read_data_valid;
	wire [31:0] _argRouteRvm_13_io_read_data_bits;
	wire _argRouteRvm_13_io_write_address_ready;
	wire _argRouteRvm_13_io_write_data_ready;
	wire _argRouteRvm_13_axi_ar_valid;
	wire [63:0] _argRouteRvm_13_axi_ar_bits_addr;
	wire _argRouteRvm_13_axi_r_ready;
	wire _argRouteRvm_13_axi_aw_valid;
	wire [63:0] _argRouteRvm_13_axi_aw_bits_addr;
	wire _argRouteRvm_13_axi_w_valid;
	wire [31:0] _argRouteRvm_13_axi_w_bits_data;
	wire _argRouteRvm_12_io_read_address_ready;
	wire _argRouteRvm_12_io_read_data_valid;
	wire [31:0] _argRouteRvm_12_io_read_data_bits;
	wire _argRouteRvm_12_io_write_address_ready;
	wire _argRouteRvm_12_io_write_data_ready;
	wire _argRouteRvm_12_axi_ar_valid;
	wire [63:0] _argRouteRvm_12_axi_ar_bits_addr;
	wire _argRouteRvm_12_axi_r_ready;
	wire _argRouteRvm_12_axi_aw_valid;
	wire [63:0] _argRouteRvm_12_axi_aw_bits_addr;
	wire _argRouteRvm_12_axi_w_valid;
	wire [31:0] _argRouteRvm_12_axi_w_bits_data;
	wire _argRouteRvm_11_io_read_address_ready;
	wire _argRouteRvm_11_io_read_data_valid;
	wire [31:0] _argRouteRvm_11_io_read_data_bits;
	wire _argRouteRvm_11_io_write_address_ready;
	wire _argRouteRvm_11_io_write_data_ready;
	wire _argRouteRvm_11_axi_ar_valid;
	wire [63:0] _argRouteRvm_11_axi_ar_bits_addr;
	wire _argRouteRvm_11_axi_r_ready;
	wire _argRouteRvm_11_axi_aw_valid;
	wire [63:0] _argRouteRvm_11_axi_aw_bits_addr;
	wire _argRouteRvm_11_axi_w_valid;
	wire [31:0] _argRouteRvm_11_axi_w_bits_data;
	wire _argRouteRvm_10_io_read_address_ready;
	wire _argRouteRvm_10_io_read_data_valid;
	wire [31:0] _argRouteRvm_10_io_read_data_bits;
	wire _argRouteRvm_10_io_write_address_ready;
	wire _argRouteRvm_10_io_write_data_ready;
	wire _argRouteRvm_10_axi_ar_valid;
	wire [63:0] _argRouteRvm_10_axi_ar_bits_addr;
	wire _argRouteRvm_10_axi_r_ready;
	wire _argRouteRvm_10_axi_aw_valid;
	wire [63:0] _argRouteRvm_10_axi_aw_bits_addr;
	wire _argRouteRvm_10_axi_w_valid;
	wire [31:0] _argRouteRvm_10_axi_w_bits_data;
	wire _argRouteRvm_9_io_read_address_ready;
	wire _argRouteRvm_9_io_read_data_valid;
	wire [31:0] _argRouteRvm_9_io_read_data_bits;
	wire _argRouteRvm_9_io_write_address_ready;
	wire _argRouteRvm_9_io_write_data_ready;
	wire _argRouteRvm_9_axi_ar_valid;
	wire [63:0] _argRouteRvm_9_axi_ar_bits_addr;
	wire _argRouteRvm_9_axi_r_ready;
	wire _argRouteRvm_9_axi_aw_valid;
	wire [63:0] _argRouteRvm_9_axi_aw_bits_addr;
	wire _argRouteRvm_9_axi_w_valid;
	wire [31:0] _argRouteRvm_9_axi_w_bits_data;
	wire _argRouteRvm_8_io_read_address_ready;
	wire _argRouteRvm_8_io_read_data_valid;
	wire [31:0] _argRouteRvm_8_io_read_data_bits;
	wire _argRouteRvm_8_io_write_address_ready;
	wire _argRouteRvm_8_io_write_data_ready;
	wire _argRouteRvm_8_axi_ar_valid;
	wire [63:0] _argRouteRvm_8_axi_ar_bits_addr;
	wire _argRouteRvm_8_axi_r_ready;
	wire _argRouteRvm_8_axi_aw_valid;
	wire [63:0] _argRouteRvm_8_axi_aw_bits_addr;
	wire _argRouteRvm_8_axi_w_valid;
	wire [31:0] _argRouteRvm_8_axi_w_bits_data;
	wire _argRouteRvm_7_io_read_address_ready;
	wire _argRouteRvm_7_io_read_data_valid;
	wire [31:0] _argRouteRvm_7_io_read_data_bits;
	wire _argRouteRvm_7_io_write_address_ready;
	wire _argRouteRvm_7_io_write_data_ready;
	wire _argRouteRvm_7_axi_ar_valid;
	wire [63:0] _argRouteRvm_7_axi_ar_bits_addr;
	wire _argRouteRvm_7_axi_r_ready;
	wire _argRouteRvm_7_axi_aw_valid;
	wire [63:0] _argRouteRvm_7_axi_aw_bits_addr;
	wire _argRouteRvm_7_axi_w_valid;
	wire [31:0] _argRouteRvm_7_axi_w_bits_data;
	wire _argRouteRvm_6_io_read_address_ready;
	wire _argRouteRvm_6_io_read_data_valid;
	wire [31:0] _argRouteRvm_6_io_read_data_bits;
	wire _argRouteRvm_6_io_write_address_ready;
	wire _argRouteRvm_6_io_write_data_ready;
	wire _argRouteRvm_6_axi_ar_valid;
	wire [63:0] _argRouteRvm_6_axi_ar_bits_addr;
	wire _argRouteRvm_6_axi_r_ready;
	wire _argRouteRvm_6_axi_aw_valid;
	wire [63:0] _argRouteRvm_6_axi_aw_bits_addr;
	wire _argRouteRvm_6_axi_w_valid;
	wire [31:0] _argRouteRvm_6_axi_w_bits_data;
	wire _argRouteRvm_5_io_read_address_ready;
	wire _argRouteRvm_5_io_read_data_valid;
	wire [31:0] _argRouteRvm_5_io_read_data_bits;
	wire _argRouteRvm_5_io_write_address_ready;
	wire _argRouteRvm_5_io_write_data_ready;
	wire _argRouteRvm_5_axi_ar_valid;
	wire [63:0] _argRouteRvm_5_axi_ar_bits_addr;
	wire _argRouteRvm_5_axi_r_ready;
	wire _argRouteRvm_5_axi_aw_valid;
	wire [63:0] _argRouteRvm_5_axi_aw_bits_addr;
	wire _argRouteRvm_5_axi_w_valid;
	wire [31:0] _argRouteRvm_5_axi_w_bits_data;
	wire _argRouteRvm_4_io_read_address_ready;
	wire _argRouteRvm_4_io_read_data_valid;
	wire [31:0] _argRouteRvm_4_io_read_data_bits;
	wire _argRouteRvm_4_io_write_address_ready;
	wire _argRouteRvm_4_io_write_data_ready;
	wire _argRouteRvm_4_axi_ar_valid;
	wire [63:0] _argRouteRvm_4_axi_ar_bits_addr;
	wire _argRouteRvm_4_axi_r_ready;
	wire _argRouteRvm_4_axi_aw_valid;
	wire [63:0] _argRouteRvm_4_axi_aw_bits_addr;
	wire _argRouteRvm_4_axi_w_valid;
	wire [31:0] _argRouteRvm_4_axi_w_bits_data;
	wire _argRouteRvm_3_io_read_address_ready;
	wire _argRouteRvm_3_io_read_data_valid;
	wire [31:0] _argRouteRvm_3_io_read_data_bits;
	wire _argRouteRvm_3_io_write_address_ready;
	wire _argRouteRvm_3_io_write_data_ready;
	wire _argRouteRvm_3_axi_ar_valid;
	wire [63:0] _argRouteRvm_3_axi_ar_bits_addr;
	wire _argRouteRvm_3_axi_r_ready;
	wire _argRouteRvm_3_axi_aw_valid;
	wire [63:0] _argRouteRvm_3_axi_aw_bits_addr;
	wire _argRouteRvm_3_axi_w_valid;
	wire [31:0] _argRouteRvm_3_axi_w_bits_data;
	wire _argRouteRvm_2_io_read_address_ready;
	wire _argRouteRvm_2_io_read_data_valid;
	wire [31:0] _argRouteRvm_2_io_read_data_bits;
	wire _argRouteRvm_2_io_write_address_ready;
	wire _argRouteRvm_2_io_write_data_ready;
	wire _argRouteRvm_2_axi_ar_valid;
	wire [63:0] _argRouteRvm_2_axi_ar_bits_addr;
	wire _argRouteRvm_2_axi_r_ready;
	wire _argRouteRvm_2_axi_aw_valid;
	wire [63:0] _argRouteRvm_2_axi_aw_bits_addr;
	wire _argRouteRvm_2_axi_w_valid;
	wire [31:0] _argRouteRvm_2_axi_w_bits_data;
	wire _argRouteRvm_1_io_read_address_ready;
	wire _argRouteRvm_1_io_read_data_valid;
	wire [31:0] _argRouteRvm_1_io_read_data_bits;
	wire _argRouteRvm_1_io_write_address_ready;
	wire _argRouteRvm_1_io_write_data_ready;
	wire _argRouteRvm_1_axi_ar_valid;
	wire [63:0] _argRouteRvm_1_axi_ar_bits_addr;
	wire _argRouteRvm_1_axi_r_ready;
	wire _argRouteRvm_1_axi_aw_valid;
	wire [63:0] _argRouteRvm_1_axi_aw_bits_addr;
	wire _argRouteRvm_1_axi_w_valid;
	wire [31:0] _argRouteRvm_1_axi_w_bits_data;
	wire _argRouteRvm_0_io_read_address_ready;
	wire _argRouteRvm_0_io_read_data_valid;
	wire [31:0] _argRouteRvm_0_io_read_data_bits;
	wire _argRouteRvm_0_io_write_address_ready;
	wire _argRouteRvm_0_io_write_data_ready;
	wire _argRouteRvm_0_axi_ar_valid;
	wire [63:0] _argRouteRvm_0_axi_ar_bits_addr;
	wire _argRouteRvm_0_axi_r_ready;
	wire _argRouteRvm_0_axi_aw_valid;
	wire [63:0] _argRouteRvm_0_axi_aw_bits_addr;
	wire _argRouteRvm_0_axi_w_valid;
	wire [31:0] _argRouteRvm_0_axi_w_bits_data;
	wire _argRouteServers_15_io_connNetwork_ready;
	wire _argRouteServers_15_io_read_address_valid;
	wire [63:0] _argRouteServers_15_io_read_address_bits;
	wire _argRouteServers_15_io_read_data_ready;
	wire _argRouteServers_15_io_write_address_valid;
	wire [63:0] _argRouteServers_15_io_write_address_bits;
	wire _argRouteServers_15_io_write_data_valid;
	wire [31:0] _argRouteServers_15_io_write_data_bits;
	wire _argRouteServers_15_io_read_address_task_valid;
	wire [63:0] _argRouteServers_15_io_read_address_task_bits;
	wire _argRouteServers_15_io_read_data_task_ready;
	wire _argRouteServers_14_io_connNetwork_ready;
	wire _argRouteServers_14_io_read_address_valid;
	wire [63:0] _argRouteServers_14_io_read_address_bits;
	wire _argRouteServers_14_io_read_data_ready;
	wire _argRouteServers_14_io_write_address_valid;
	wire [63:0] _argRouteServers_14_io_write_address_bits;
	wire _argRouteServers_14_io_write_data_valid;
	wire [31:0] _argRouteServers_14_io_write_data_bits;
	wire _argRouteServers_14_io_read_address_task_valid;
	wire [63:0] _argRouteServers_14_io_read_address_task_bits;
	wire _argRouteServers_14_io_read_data_task_ready;
	wire _argRouteServers_13_io_connNetwork_ready;
	wire _argRouteServers_13_io_read_address_valid;
	wire [63:0] _argRouteServers_13_io_read_address_bits;
	wire _argRouteServers_13_io_read_data_ready;
	wire _argRouteServers_13_io_write_address_valid;
	wire [63:0] _argRouteServers_13_io_write_address_bits;
	wire _argRouteServers_13_io_write_data_valid;
	wire [31:0] _argRouteServers_13_io_write_data_bits;
	wire _argRouteServers_13_io_read_address_task_valid;
	wire [63:0] _argRouteServers_13_io_read_address_task_bits;
	wire _argRouteServers_13_io_read_data_task_ready;
	wire _argRouteServers_12_io_connNetwork_ready;
	wire _argRouteServers_12_io_read_address_valid;
	wire [63:0] _argRouteServers_12_io_read_address_bits;
	wire _argRouteServers_12_io_read_data_ready;
	wire _argRouteServers_12_io_write_address_valid;
	wire [63:0] _argRouteServers_12_io_write_address_bits;
	wire _argRouteServers_12_io_write_data_valid;
	wire [31:0] _argRouteServers_12_io_write_data_bits;
	wire _argRouteServers_12_io_read_address_task_valid;
	wire [63:0] _argRouteServers_12_io_read_address_task_bits;
	wire _argRouteServers_12_io_read_data_task_ready;
	wire _argRouteServers_11_io_connNetwork_ready;
	wire _argRouteServers_11_io_read_address_valid;
	wire [63:0] _argRouteServers_11_io_read_address_bits;
	wire _argRouteServers_11_io_read_data_ready;
	wire _argRouteServers_11_io_write_address_valid;
	wire [63:0] _argRouteServers_11_io_write_address_bits;
	wire _argRouteServers_11_io_write_data_valid;
	wire [31:0] _argRouteServers_11_io_write_data_bits;
	wire _argRouteServers_11_io_read_address_task_valid;
	wire [63:0] _argRouteServers_11_io_read_address_task_bits;
	wire _argRouteServers_11_io_read_data_task_ready;
	wire _argRouteServers_10_io_connNetwork_ready;
	wire _argRouteServers_10_io_read_address_valid;
	wire [63:0] _argRouteServers_10_io_read_address_bits;
	wire _argRouteServers_10_io_read_data_ready;
	wire _argRouteServers_10_io_write_address_valid;
	wire [63:0] _argRouteServers_10_io_write_address_bits;
	wire _argRouteServers_10_io_write_data_valid;
	wire [31:0] _argRouteServers_10_io_write_data_bits;
	wire _argRouteServers_10_io_read_address_task_valid;
	wire [63:0] _argRouteServers_10_io_read_address_task_bits;
	wire _argRouteServers_10_io_read_data_task_ready;
	wire _argRouteServers_9_io_connNetwork_ready;
	wire _argRouteServers_9_io_read_address_valid;
	wire [63:0] _argRouteServers_9_io_read_address_bits;
	wire _argRouteServers_9_io_read_data_ready;
	wire _argRouteServers_9_io_write_address_valid;
	wire [63:0] _argRouteServers_9_io_write_address_bits;
	wire _argRouteServers_9_io_write_data_valid;
	wire [31:0] _argRouteServers_9_io_write_data_bits;
	wire _argRouteServers_9_io_read_address_task_valid;
	wire [63:0] _argRouteServers_9_io_read_address_task_bits;
	wire _argRouteServers_9_io_read_data_task_ready;
	wire _argRouteServers_8_io_connNetwork_ready;
	wire _argRouteServers_8_io_read_address_valid;
	wire [63:0] _argRouteServers_8_io_read_address_bits;
	wire _argRouteServers_8_io_read_data_ready;
	wire _argRouteServers_8_io_write_address_valid;
	wire [63:0] _argRouteServers_8_io_write_address_bits;
	wire _argRouteServers_8_io_write_data_valid;
	wire [31:0] _argRouteServers_8_io_write_data_bits;
	wire _argRouteServers_8_io_read_address_task_valid;
	wire [63:0] _argRouteServers_8_io_read_address_task_bits;
	wire _argRouteServers_8_io_read_data_task_ready;
	wire _argRouteServers_7_io_connNetwork_ready;
	wire _argRouteServers_7_io_read_address_valid;
	wire [63:0] _argRouteServers_7_io_read_address_bits;
	wire _argRouteServers_7_io_read_data_ready;
	wire _argRouteServers_7_io_write_address_valid;
	wire [63:0] _argRouteServers_7_io_write_address_bits;
	wire _argRouteServers_7_io_write_data_valid;
	wire [31:0] _argRouteServers_7_io_write_data_bits;
	wire _argRouteServers_7_io_read_address_task_valid;
	wire [63:0] _argRouteServers_7_io_read_address_task_bits;
	wire _argRouteServers_7_io_read_data_task_ready;
	wire _argRouteServers_6_io_connNetwork_ready;
	wire _argRouteServers_6_io_read_address_valid;
	wire [63:0] _argRouteServers_6_io_read_address_bits;
	wire _argRouteServers_6_io_read_data_ready;
	wire _argRouteServers_6_io_write_address_valid;
	wire [63:0] _argRouteServers_6_io_write_address_bits;
	wire _argRouteServers_6_io_write_data_valid;
	wire [31:0] _argRouteServers_6_io_write_data_bits;
	wire _argRouteServers_6_io_read_address_task_valid;
	wire [63:0] _argRouteServers_6_io_read_address_task_bits;
	wire _argRouteServers_6_io_read_data_task_ready;
	wire _argRouteServers_5_io_connNetwork_ready;
	wire _argRouteServers_5_io_read_address_valid;
	wire [63:0] _argRouteServers_5_io_read_address_bits;
	wire _argRouteServers_5_io_read_data_ready;
	wire _argRouteServers_5_io_write_address_valid;
	wire [63:0] _argRouteServers_5_io_write_address_bits;
	wire _argRouteServers_5_io_write_data_valid;
	wire [31:0] _argRouteServers_5_io_write_data_bits;
	wire _argRouteServers_5_io_read_address_task_valid;
	wire [63:0] _argRouteServers_5_io_read_address_task_bits;
	wire _argRouteServers_5_io_read_data_task_ready;
	wire _argRouteServers_4_io_connNetwork_ready;
	wire _argRouteServers_4_io_read_address_valid;
	wire [63:0] _argRouteServers_4_io_read_address_bits;
	wire _argRouteServers_4_io_read_data_ready;
	wire _argRouteServers_4_io_write_address_valid;
	wire [63:0] _argRouteServers_4_io_write_address_bits;
	wire _argRouteServers_4_io_write_data_valid;
	wire [31:0] _argRouteServers_4_io_write_data_bits;
	wire _argRouteServers_4_io_read_address_task_valid;
	wire [63:0] _argRouteServers_4_io_read_address_task_bits;
	wire _argRouteServers_4_io_read_data_task_ready;
	wire _argRouteServers_3_io_connNetwork_ready;
	wire _argRouteServers_3_io_read_address_valid;
	wire [63:0] _argRouteServers_3_io_read_address_bits;
	wire _argRouteServers_3_io_read_data_ready;
	wire _argRouteServers_3_io_write_address_valid;
	wire [63:0] _argRouteServers_3_io_write_address_bits;
	wire _argRouteServers_3_io_write_data_valid;
	wire [31:0] _argRouteServers_3_io_write_data_bits;
	wire _argRouteServers_3_io_read_address_task_valid;
	wire [63:0] _argRouteServers_3_io_read_address_task_bits;
	wire _argRouteServers_3_io_read_data_task_ready;
	wire _argRouteServers_2_io_connNetwork_ready;
	wire _argRouteServers_2_io_read_address_valid;
	wire [63:0] _argRouteServers_2_io_read_address_bits;
	wire _argRouteServers_2_io_read_data_ready;
	wire _argRouteServers_2_io_write_address_valid;
	wire [63:0] _argRouteServers_2_io_write_address_bits;
	wire _argRouteServers_2_io_write_data_valid;
	wire [31:0] _argRouteServers_2_io_write_data_bits;
	wire _argRouteServers_2_io_read_address_task_valid;
	wire [63:0] _argRouteServers_2_io_read_address_task_bits;
	wire _argRouteServers_2_io_read_data_task_ready;
	wire _argRouteServers_1_io_connNetwork_ready;
	wire _argRouteServers_1_io_read_address_valid;
	wire [63:0] _argRouteServers_1_io_read_address_bits;
	wire _argRouteServers_1_io_read_data_ready;
	wire _argRouteServers_1_io_write_address_valid;
	wire [63:0] _argRouteServers_1_io_write_address_bits;
	wire _argRouteServers_1_io_write_data_valid;
	wire [31:0] _argRouteServers_1_io_write_data_bits;
	wire _argRouteServers_1_io_read_address_task_valid;
	wire [63:0] _argRouteServers_1_io_read_address_task_bits;
	wire _argRouteServers_1_io_read_data_task_ready;
	wire _argRouteServers_0_io_connNetwork_ready;
	wire _argRouteServers_0_io_read_address_valid;
	wire [63:0] _argRouteServers_0_io_read_address_bits;
	wire _argRouteServers_0_io_read_data_ready;
	wire _argRouteServers_0_io_write_address_valid;
	wire [63:0] _argRouteServers_0_io_write_address_bits;
	wire _argRouteServers_0_io_write_data_valid;
	wire [31:0] _argRouteServers_0_io_write_data_bits;
	wire _argRouteServers_0_io_read_address_task_valid;
	wire [63:0] _argRouteServers_0_io_read_address_task_bits;
	wire _argRouteServers_0_io_read_data_task_ready;
	wire _argSide_io_connVAS_0_valid;
	wire [63:0] _argSide_io_connVAS_0_bits;
	wire _argSide_io_connVAS_1_valid;
	wire [63:0] _argSide_io_connVAS_1_bits;
	wire _argSide_io_connVAS_2_valid;
	wire [63:0] _argSide_io_connVAS_2_bits;
	wire _argSide_io_connVAS_3_valid;
	wire [63:0] _argSide_io_connVAS_3_bits;
	wire _argSide_io_connVAS_4_valid;
	wire [63:0] _argSide_io_connVAS_4_bits;
	wire _argSide_io_connVAS_5_valid;
	wire [63:0] _argSide_io_connVAS_5_bits;
	wire _argSide_io_connVAS_6_valid;
	wire [63:0] _argSide_io_connVAS_6_bits;
	wire _argSide_io_connVAS_7_valid;
	wire [63:0] _argSide_io_connVAS_7_bits;
	wire _argSide_io_connVAS_8_valid;
	wire [63:0] _argSide_io_connVAS_8_bits;
	wire _argSide_io_connVAS_9_valid;
	wire [63:0] _argSide_io_connVAS_9_bits;
	wire _argSide_io_connVAS_10_valid;
	wire [63:0] _argSide_io_connVAS_10_bits;
	wire _argSide_io_connVAS_11_valid;
	wire [63:0] _argSide_io_connVAS_11_bits;
	wire _argSide_io_connVAS_12_valid;
	wire [63:0] _argSide_io_connVAS_12_bits;
	wire _argSide_io_connVAS_13_valid;
	wire [63:0] _argSide_io_connVAS_13_bits;
	wire _argSide_io_connVAS_14_valid;
	wire [63:0] _argSide_io_connVAS_14_bits;
	wire _argSide_io_connVAS_15_valid;
	wire [63:0] _argSide_io_connVAS_15_bits;
	wire _argSide_io_connPE_0_ready;
	wire _argSide_io_connPE_1_ready;
	wire _argSide_io_connPE_2_ready;
	wire _argSide_io_connPE_3_ready;
	wire _argSide_io_connPE_4_ready;
	wire _argSide_io_connPE_5_ready;
	wire _argSide_io_connPE_6_ready;
	wire _argSide_io_connPE_7_ready;
	wire _argSide_io_connPE_8_ready;
	wire _argSide_io_connPE_9_ready;
	wire _argSide_io_connPE_10_ready;
	wire _argSide_io_connPE_11_ready;
	wire _argSide_io_connPE_12_ready;
	wire _argSide_io_connPE_13_ready;
	wire _argSide_io_connPE_14_ready;
	wire _argSide_io_connPE_15_ready;
	wire _argSide_io_connPE_16_ready;
	wire _argSide_io_connPE_17_ready;
	wire _argSide_io_connPE_18_ready;
	wire _argSide_io_connPE_19_ready;
	wire _argSide_io_connPE_20_ready;
	wire _argSide_io_connPE_21_ready;
	wire _argSide_io_connPE_22_ready;
	wire _argSide_io_connPE_23_ready;
	wire _argSide_io_connPE_24_ready;
	wire _argSide_io_connPE_25_ready;
	wire _argSide_io_connPE_26_ready;
	wire _argSide_io_connPE_27_ready;
	wire _argSide_io_connPE_28_ready;
	wire _argSide_io_connPE_29_ready;
	wire _argSide_io_connPE_30_ready;
	wire _argSide_io_connPE_31_ready;
	wire _argSide_io_connPE_32_ready;
	wire _argSide_io_connPE_33_ready;
	wire _argSide_io_connPE_34_ready;
	wire _argSide_io_connPE_35_ready;
	wire _argSide_io_connPE_36_ready;
	wire _argSide_io_connPE_37_ready;
	wire _argSide_io_connPE_38_ready;
	wire _argSide_io_connPE_39_ready;
	wire _argSide_io_connPE_40_ready;
	wire _argSide_io_connPE_41_ready;
	wire _argSide_io_connPE_42_ready;
	wire _argSide_io_connPE_43_ready;
	wire _argSide_io_connPE_44_ready;
	wire _argSide_io_connPE_45_ready;
	wire _argSide_io_connPE_46_ready;
	wire _argSide_io_connPE_47_ready;
	wire _argSide_io_connPE_48_ready;
	wire _argSide_io_connPE_49_ready;
	wire _argSide_io_connPE_50_ready;
	wire _argSide_io_connPE_51_ready;
	wire _argSide_io_connPE_52_ready;
	wire _argSide_io_connPE_53_ready;
	wire _argSide_io_connPE_54_ready;
	wire _argSide_io_connPE_55_ready;
	wire _argSide_io_connPE_56_ready;
	wire _argSide_io_connPE_57_ready;
	wire _argSide_io_connPE_58_ready;
	wire _argSide_io_connPE_59_ready;
	wire _argSide_io_connPE_60_ready;
	wire _argSide_io_connPE_61_ready;
	wire _argSide_io_connPE_62_ready;
	wire _argSide_io_connPE_63_ready;
	wire _argSide_io_connPE_64_ready;
	wire _argSide_io_connPE_65_ready;
	wire _argSide_io_connPE_66_ready;
	wire _argSide_io_connPE_67_ready;
	wire _argSide_io_connPE_68_ready;
	wire _argSide_io_connPE_69_ready;
	wire _argSide_io_connPE_70_ready;
	wire _argSide_io_connPE_71_ready;
	wire _argSide_io_connPE_72_ready;
	wire _argSide_io_connPE_73_ready;
	wire _argSide_io_connPE_74_ready;
	wire _argSide_io_connPE_75_ready;
	wire _argSide_io_connPE_76_ready;
	wire _argSide_io_connPE_77_ready;
	wire _argSide_io_connPE_78_ready;
	wire _argSide_io_connPE_79_ready;
	wire _argSide_io_connPE_80_ready;
	wire _argSide_io_connPE_81_ready;
	wire _argSide_io_connPE_82_ready;
	wire _argSide_io_connPE_83_ready;
	wire _argSide_io_connPE_84_ready;
	wire _argSide_io_connPE_85_ready;
	wire _argSide_io_connPE_86_ready;
	wire _argSide_io_connPE_87_ready;
	wire _argSide_io_connPE_88_ready;
	wire _argSide_io_connPE_89_ready;
	wire _argSide_io_connPE_90_ready;
	wire _argSide_io_connPE_91_ready;
	wire _argSide_io_connPE_92_ready;
	wire _argSide_io_connPE_93_ready;
	wire _argSide_io_connPE_94_ready;
	wire _argSide_io_connPE_95_ready;
	wire _argSide_io_connPE_96_ready;
	wire _argSide_io_connPE_97_ready;
	wire _argSide_io_connPE_98_ready;
	wire _argSide_io_connPE_99_ready;
	wire _argSide_io_connPE_100_ready;
	wire _argSide_io_connPE_101_ready;
	wire _argSide_io_connPE_102_ready;
	wire _argSide_io_connPE_103_ready;
	wire _argSide_io_connPE_104_ready;
	wire _argSide_io_connPE_105_ready;
	wire _argSide_io_connPE_106_ready;
	wire _argSide_io_connPE_107_ready;
	wire _argSide_io_connPE_108_ready;
	wire _argSide_io_connPE_109_ready;
	wire _argSide_io_connPE_110_ready;
	wire _argSide_io_connPE_111_ready;
	wire _argSide_io_connPE_112_ready;
	wire _argSide_io_connPE_113_ready;
	wire _argSide_io_connPE_114_ready;
	wire _argSide_io_connPE_115_ready;
	wire _argSide_io_connPE_116_ready;
	wire _argSide_io_connPE_117_ready;
	wire _argSide_io_connPE_118_ready;
	wire _argSide_io_connPE_119_ready;
	wire _argSide_io_connPE_120_ready;
	wire _argSide_io_connPE_121_ready;
	wire _argSide_io_connPE_122_ready;
	wire _argSide_io_connPE_123_ready;
	wire _argSide_io_connPE_124_ready;
	wire _argSide_io_connPE_125_ready;
	wire _argSide_io_connPE_126_ready;
	wire _argSide_io_connPE_127_ready;
	ArgumentNotifierNetwork argSide(
		.clock(clock),
		.reset(reset),
		.io_connVAS_0_ready(_argRouteServers_0_io_connNetwork_ready),
		.io_connVAS_0_valid(_argSide_io_connVAS_0_valid),
		.io_connVAS_0_bits(_argSide_io_connVAS_0_bits),
		.io_connVAS_1_ready(_argRouteServers_1_io_connNetwork_ready),
		.io_connVAS_1_valid(_argSide_io_connVAS_1_valid),
		.io_connVAS_1_bits(_argSide_io_connVAS_1_bits),
		.io_connVAS_2_ready(_argRouteServers_2_io_connNetwork_ready),
		.io_connVAS_2_valid(_argSide_io_connVAS_2_valid),
		.io_connVAS_2_bits(_argSide_io_connVAS_2_bits),
		.io_connVAS_3_ready(_argRouteServers_3_io_connNetwork_ready),
		.io_connVAS_3_valid(_argSide_io_connVAS_3_valid),
		.io_connVAS_3_bits(_argSide_io_connVAS_3_bits),
		.io_connVAS_4_ready(_argRouteServers_4_io_connNetwork_ready),
		.io_connVAS_4_valid(_argSide_io_connVAS_4_valid),
		.io_connVAS_4_bits(_argSide_io_connVAS_4_bits),
		.io_connVAS_5_ready(_argRouteServers_5_io_connNetwork_ready),
		.io_connVAS_5_valid(_argSide_io_connVAS_5_valid),
		.io_connVAS_5_bits(_argSide_io_connVAS_5_bits),
		.io_connVAS_6_ready(_argRouteServers_6_io_connNetwork_ready),
		.io_connVAS_6_valid(_argSide_io_connVAS_6_valid),
		.io_connVAS_6_bits(_argSide_io_connVAS_6_bits),
		.io_connVAS_7_ready(_argRouteServers_7_io_connNetwork_ready),
		.io_connVAS_7_valid(_argSide_io_connVAS_7_valid),
		.io_connVAS_7_bits(_argSide_io_connVAS_7_bits),
		.io_connVAS_8_ready(_argRouteServers_8_io_connNetwork_ready),
		.io_connVAS_8_valid(_argSide_io_connVAS_8_valid),
		.io_connVAS_8_bits(_argSide_io_connVAS_8_bits),
		.io_connVAS_9_ready(_argRouteServers_9_io_connNetwork_ready),
		.io_connVAS_9_valid(_argSide_io_connVAS_9_valid),
		.io_connVAS_9_bits(_argSide_io_connVAS_9_bits),
		.io_connVAS_10_ready(_argRouteServers_10_io_connNetwork_ready),
		.io_connVAS_10_valid(_argSide_io_connVAS_10_valid),
		.io_connVAS_10_bits(_argSide_io_connVAS_10_bits),
		.io_connVAS_11_ready(_argRouteServers_11_io_connNetwork_ready),
		.io_connVAS_11_valid(_argSide_io_connVAS_11_valid),
		.io_connVAS_11_bits(_argSide_io_connVAS_11_bits),
		.io_connVAS_12_ready(_argRouteServers_12_io_connNetwork_ready),
		.io_connVAS_12_valid(_argSide_io_connVAS_12_valid),
		.io_connVAS_12_bits(_argSide_io_connVAS_12_bits),
		.io_connVAS_13_ready(_argRouteServers_13_io_connNetwork_ready),
		.io_connVAS_13_valid(_argSide_io_connVAS_13_valid),
		.io_connVAS_13_bits(_argSide_io_connVAS_13_bits),
		.io_connVAS_14_ready(_argRouteServers_14_io_connNetwork_ready),
		.io_connVAS_14_valid(_argSide_io_connVAS_14_valid),
		.io_connVAS_14_bits(_argSide_io_connVAS_14_bits),
		.io_connVAS_15_ready(_argRouteServers_15_io_connNetwork_ready),
		.io_connVAS_15_valid(_argSide_io_connVAS_15_valid),
		.io_connVAS_15_bits(_argSide_io_connVAS_15_bits),
		.io_connPE_0_ready(_argSide_io_connPE_0_ready),
		.io_connPE_0_valid(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_connPE_0_bits(_axis_stream_converters_in_0_io_dataOut_TDATA),
		.io_connPE_1_ready(_argSide_io_connPE_1_ready),
		.io_connPE_1_valid(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_connPE_1_bits(_axis_stream_converters_in_1_io_dataOut_TDATA),
		.io_connPE_2_ready(_argSide_io_connPE_2_ready),
		.io_connPE_2_valid(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_connPE_2_bits(_axis_stream_converters_in_2_io_dataOut_TDATA),
		.io_connPE_3_ready(_argSide_io_connPE_3_ready),
		.io_connPE_3_valid(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_connPE_3_bits(_axis_stream_converters_in_3_io_dataOut_TDATA),
		.io_connPE_4_ready(_argSide_io_connPE_4_ready),
		.io_connPE_4_valid(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_connPE_4_bits(_axis_stream_converters_in_4_io_dataOut_TDATA),
		.io_connPE_5_ready(_argSide_io_connPE_5_ready),
		.io_connPE_5_valid(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_connPE_5_bits(_axis_stream_converters_in_5_io_dataOut_TDATA),
		.io_connPE_6_ready(_argSide_io_connPE_6_ready),
		.io_connPE_6_valid(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_connPE_6_bits(_axis_stream_converters_in_6_io_dataOut_TDATA),
		.io_connPE_7_ready(_argSide_io_connPE_7_ready),
		.io_connPE_7_valid(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_connPE_7_bits(_axis_stream_converters_in_7_io_dataOut_TDATA),
		.io_connPE_8_ready(_argSide_io_connPE_8_ready),
		.io_connPE_8_valid(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_connPE_8_bits(_axis_stream_converters_in_8_io_dataOut_TDATA),
		.io_connPE_9_ready(_argSide_io_connPE_9_ready),
		.io_connPE_9_valid(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_connPE_9_bits(_axis_stream_converters_in_9_io_dataOut_TDATA),
		.io_connPE_10_ready(_argSide_io_connPE_10_ready),
		.io_connPE_10_valid(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_connPE_10_bits(_axis_stream_converters_in_10_io_dataOut_TDATA),
		.io_connPE_11_ready(_argSide_io_connPE_11_ready),
		.io_connPE_11_valid(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_connPE_11_bits(_axis_stream_converters_in_11_io_dataOut_TDATA),
		.io_connPE_12_ready(_argSide_io_connPE_12_ready),
		.io_connPE_12_valid(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_connPE_12_bits(_axis_stream_converters_in_12_io_dataOut_TDATA),
		.io_connPE_13_ready(_argSide_io_connPE_13_ready),
		.io_connPE_13_valid(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_connPE_13_bits(_axis_stream_converters_in_13_io_dataOut_TDATA),
		.io_connPE_14_ready(_argSide_io_connPE_14_ready),
		.io_connPE_14_valid(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_connPE_14_bits(_axis_stream_converters_in_14_io_dataOut_TDATA),
		.io_connPE_15_ready(_argSide_io_connPE_15_ready),
		.io_connPE_15_valid(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_connPE_15_bits(_axis_stream_converters_in_15_io_dataOut_TDATA),
		.io_connPE_16_ready(_argSide_io_connPE_16_ready),
		.io_connPE_16_valid(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_connPE_16_bits(_axis_stream_converters_in_16_io_dataOut_TDATA),
		.io_connPE_17_ready(_argSide_io_connPE_17_ready),
		.io_connPE_17_valid(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_connPE_17_bits(_axis_stream_converters_in_17_io_dataOut_TDATA),
		.io_connPE_18_ready(_argSide_io_connPE_18_ready),
		.io_connPE_18_valid(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_connPE_18_bits(_axis_stream_converters_in_18_io_dataOut_TDATA),
		.io_connPE_19_ready(_argSide_io_connPE_19_ready),
		.io_connPE_19_valid(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_connPE_19_bits(_axis_stream_converters_in_19_io_dataOut_TDATA),
		.io_connPE_20_ready(_argSide_io_connPE_20_ready),
		.io_connPE_20_valid(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_connPE_20_bits(_axis_stream_converters_in_20_io_dataOut_TDATA),
		.io_connPE_21_ready(_argSide_io_connPE_21_ready),
		.io_connPE_21_valid(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_connPE_21_bits(_axis_stream_converters_in_21_io_dataOut_TDATA),
		.io_connPE_22_ready(_argSide_io_connPE_22_ready),
		.io_connPE_22_valid(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_connPE_22_bits(_axis_stream_converters_in_22_io_dataOut_TDATA),
		.io_connPE_23_ready(_argSide_io_connPE_23_ready),
		.io_connPE_23_valid(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_connPE_23_bits(_axis_stream_converters_in_23_io_dataOut_TDATA),
		.io_connPE_24_ready(_argSide_io_connPE_24_ready),
		.io_connPE_24_valid(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_connPE_24_bits(_axis_stream_converters_in_24_io_dataOut_TDATA),
		.io_connPE_25_ready(_argSide_io_connPE_25_ready),
		.io_connPE_25_valid(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_connPE_25_bits(_axis_stream_converters_in_25_io_dataOut_TDATA),
		.io_connPE_26_ready(_argSide_io_connPE_26_ready),
		.io_connPE_26_valid(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_connPE_26_bits(_axis_stream_converters_in_26_io_dataOut_TDATA),
		.io_connPE_27_ready(_argSide_io_connPE_27_ready),
		.io_connPE_27_valid(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_connPE_27_bits(_axis_stream_converters_in_27_io_dataOut_TDATA),
		.io_connPE_28_ready(_argSide_io_connPE_28_ready),
		.io_connPE_28_valid(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_connPE_28_bits(_axis_stream_converters_in_28_io_dataOut_TDATA),
		.io_connPE_29_ready(_argSide_io_connPE_29_ready),
		.io_connPE_29_valid(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_connPE_29_bits(_axis_stream_converters_in_29_io_dataOut_TDATA),
		.io_connPE_30_ready(_argSide_io_connPE_30_ready),
		.io_connPE_30_valid(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_connPE_30_bits(_axis_stream_converters_in_30_io_dataOut_TDATA),
		.io_connPE_31_ready(_argSide_io_connPE_31_ready),
		.io_connPE_31_valid(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_connPE_31_bits(_axis_stream_converters_in_31_io_dataOut_TDATA),
		.io_connPE_32_ready(_argSide_io_connPE_32_ready),
		.io_connPE_32_valid(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_connPE_32_bits(_axis_stream_converters_in_32_io_dataOut_TDATA),
		.io_connPE_33_ready(_argSide_io_connPE_33_ready),
		.io_connPE_33_valid(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_connPE_33_bits(_axis_stream_converters_in_33_io_dataOut_TDATA),
		.io_connPE_34_ready(_argSide_io_connPE_34_ready),
		.io_connPE_34_valid(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_connPE_34_bits(_axis_stream_converters_in_34_io_dataOut_TDATA),
		.io_connPE_35_ready(_argSide_io_connPE_35_ready),
		.io_connPE_35_valid(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_connPE_35_bits(_axis_stream_converters_in_35_io_dataOut_TDATA),
		.io_connPE_36_ready(_argSide_io_connPE_36_ready),
		.io_connPE_36_valid(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_connPE_36_bits(_axis_stream_converters_in_36_io_dataOut_TDATA),
		.io_connPE_37_ready(_argSide_io_connPE_37_ready),
		.io_connPE_37_valid(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_connPE_37_bits(_axis_stream_converters_in_37_io_dataOut_TDATA),
		.io_connPE_38_ready(_argSide_io_connPE_38_ready),
		.io_connPE_38_valid(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_connPE_38_bits(_axis_stream_converters_in_38_io_dataOut_TDATA),
		.io_connPE_39_ready(_argSide_io_connPE_39_ready),
		.io_connPE_39_valid(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_connPE_39_bits(_axis_stream_converters_in_39_io_dataOut_TDATA),
		.io_connPE_40_ready(_argSide_io_connPE_40_ready),
		.io_connPE_40_valid(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_connPE_40_bits(_axis_stream_converters_in_40_io_dataOut_TDATA),
		.io_connPE_41_ready(_argSide_io_connPE_41_ready),
		.io_connPE_41_valid(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_connPE_41_bits(_axis_stream_converters_in_41_io_dataOut_TDATA),
		.io_connPE_42_ready(_argSide_io_connPE_42_ready),
		.io_connPE_42_valid(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_connPE_42_bits(_axis_stream_converters_in_42_io_dataOut_TDATA),
		.io_connPE_43_ready(_argSide_io_connPE_43_ready),
		.io_connPE_43_valid(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_connPE_43_bits(_axis_stream_converters_in_43_io_dataOut_TDATA),
		.io_connPE_44_ready(_argSide_io_connPE_44_ready),
		.io_connPE_44_valid(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_connPE_44_bits(_axis_stream_converters_in_44_io_dataOut_TDATA),
		.io_connPE_45_ready(_argSide_io_connPE_45_ready),
		.io_connPE_45_valid(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_connPE_45_bits(_axis_stream_converters_in_45_io_dataOut_TDATA),
		.io_connPE_46_ready(_argSide_io_connPE_46_ready),
		.io_connPE_46_valid(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_connPE_46_bits(_axis_stream_converters_in_46_io_dataOut_TDATA),
		.io_connPE_47_ready(_argSide_io_connPE_47_ready),
		.io_connPE_47_valid(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_connPE_47_bits(_axis_stream_converters_in_47_io_dataOut_TDATA),
		.io_connPE_48_ready(_argSide_io_connPE_48_ready),
		.io_connPE_48_valid(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_connPE_48_bits(_axis_stream_converters_in_48_io_dataOut_TDATA),
		.io_connPE_49_ready(_argSide_io_connPE_49_ready),
		.io_connPE_49_valid(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_connPE_49_bits(_axis_stream_converters_in_49_io_dataOut_TDATA),
		.io_connPE_50_ready(_argSide_io_connPE_50_ready),
		.io_connPE_50_valid(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_connPE_50_bits(_axis_stream_converters_in_50_io_dataOut_TDATA),
		.io_connPE_51_ready(_argSide_io_connPE_51_ready),
		.io_connPE_51_valid(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_connPE_51_bits(_axis_stream_converters_in_51_io_dataOut_TDATA),
		.io_connPE_52_ready(_argSide_io_connPE_52_ready),
		.io_connPE_52_valid(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_connPE_52_bits(_axis_stream_converters_in_52_io_dataOut_TDATA),
		.io_connPE_53_ready(_argSide_io_connPE_53_ready),
		.io_connPE_53_valid(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_connPE_53_bits(_axis_stream_converters_in_53_io_dataOut_TDATA),
		.io_connPE_54_ready(_argSide_io_connPE_54_ready),
		.io_connPE_54_valid(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_connPE_54_bits(_axis_stream_converters_in_54_io_dataOut_TDATA),
		.io_connPE_55_ready(_argSide_io_connPE_55_ready),
		.io_connPE_55_valid(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_connPE_55_bits(_axis_stream_converters_in_55_io_dataOut_TDATA),
		.io_connPE_56_ready(_argSide_io_connPE_56_ready),
		.io_connPE_56_valid(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_connPE_56_bits(_axis_stream_converters_in_56_io_dataOut_TDATA),
		.io_connPE_57_ready(_argSide_io_connPE_57_ready),
		.io_connPE_57_valid(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_connPE_57_bits(_axis_stream_converters_in_57_io_dataOut_TDATA),
		.io_connPE_58_ready(_argSide_io_connPE_58_ready),
		.io_connPE_58_valid(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_connPE_58_bits(_axis_stream_converters_in_58_io_dataOut_TDATA),
		.io_connPE_59_ready(_argSide_io_connPE_59_ready),
		.io_connPE_59_valid(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_connPE_59_bits(_axis_stream_converters_in_59_io_dataOut_TDATA),
		.io_connPE_60_ready(_argSide_io_connPE_60_ready),
		.io_connPE_60_valid(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_connPE_60_bits(_axis_stream_converters_in_60_io_dataOut_TDATA),
		.io_connPE_61_ready(_argSide_io_connPE_61_ready),
		.io_connPE_61_valid(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_connPE_61_bits(_axis_stream_converters_in_61_io_dataOut_TDATA),
		.io_connPE_62_ready(_argSide_io_connPE_62_ready),
		.io_connPE_62_valid(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_connPE_62_bits(_axis_stream_converters_in_62_io_dataOut_TDATA),
		.io_connPE_63_ready(_argSide_io_connPE_63_ready),
		.io_connPE_63_valid(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_connPE_63_bits(_axis_stream_converters_in_63_io_dataOut_TDATA),
		.io_connPE_64_ready(_argSide_io_connPE_64_ready),
		.io_connPE_64_valid(_axis_stream_converters_in_64_io_dataOut_TVALID),
		.io_connPE_64_bits(_axis_stream_converters_in_64_io_dataOut_TDATA),
		.io_connPE_65_ready(_argSide_io_connPE_65_ready),
		.io_connPE_65_valid(_axis_stream_converters_in_65_io_dataOut_TVALID),
		.io_connPE_65_bits(_axis_stream_converters_in_65_io_dataOut_TDATA),
		.io_connPE_66_ready(_argSide_io_connPE_66_ready),
		.io_connPE_66_valid(_axis_stream_converters_in_66_io_dataOut_TVALID),
		.io_connPE_66_bits(_axis_stream_converters_in_66_io_dataOut_TDATA),
		.io_connPE_67_ready(_argSide_io_connPE_67_ready),
		.io_connPE_67_valid(_axis_stream_converters_in_67_io_dataOut_TVALID),
		.io_connPE_67_bits(_axis_stream_converters_in_67_io_dataOut_TDATA),
		.io_connPE_68_ready(_argSide_io_connPE_68_ready),
		.io_connPE_68_valid(_axis_stream_converters_in_68_io_dataOut_TVALID),
		.io_connPE_68_bits(_axis_stream_converters_in_68_io_dataOut_TDATA),
		.io_connPE_69_ready(_argSide_io_connPE_69_ready),
		.io_connPE_69_valid(_axis_stream_converters_in_69_io_dataOut_TVALID),
		.io_connPE_69_bits(_axis_stream_converters_in_69_io_dataOut_TDATA),
		.io_connPE_70_ready(_argSide_io_connPE_70_ready),
		.io_connPE_70_valid(_axis_stream_converters_in_70_io_dataOut_TVALID),
		.io_connPE_70_bits(_axis_stream_converters_in_70_io_dataOut_TDATA),
		.io_connPE_71_ready(_argSide_io_connPE_71_ready),
		.io_connPE_71_valid(_axis_stream_converters_in_71_io_dataOut_TVALID),
		.io_connPE_71_bits(_axis_stream_converters_in_71_io_dataOut_TDATA),
		.io_connPE_72_ready(_argSide_io_connPE_72_ready),
		.io_connPE_72_valid(_axis_stream_converters_in_72_io_dataOut_TVALID),
		.io_connPE_72_bits(_axis_stream_converters_in_72_io_dataOut_TDATA),
		.io_connPE_73_ready(_argSide_io_connPE_73_ready),
		.io_connPE_73_valid(_axis_stream_converters_in_73_io_dataOut_TVALID),
		.io_connPE_73_bits(_axis_stream_converters_in_73_io_dataOut_TDATA),
		.io_connPE_74_ready(_argSide_io_connPE_74_ready),
		.io_connPE_74_valid(_axis_stream_converters_in_74_io_dataOut_TVALID),
		.io_connPE_74_bits(_axis_stream_converters_in_74_io_dataOut_TDATA),
		.io_connPE_75_ready(_argSide_io_connPE_75_ready),
		.io_connPE_75_valid(_axis_stream_converters_in_75_io_dataOut_TVALID),
		.io_connPE_75_bits(_axis_stream_converters_in_75_io_dataOut_TDATA),
		.io_connPE_76_ready(_argSide_io_connPE_76_ready),
		.io_connPE_76_valid(_axis_stream_converters_in_76_io_dataOut_TVALID),
		.io_connPE_76_bits(_axis_stream_converters_in_76_io_dataOut_TDATA),
		.io_connPE_77_ready(_argSide_io_connPE_77_ready),
		.io_connPE_77_valid(_axis_stream_converters_in_77_io_dataOut_TVALID),
		.io_connPE_77_bits(_axis_stream_converters_in_77_io_dataOut_TDATA),
		.io_connPE_78_ready(_argSide_io_connPE_78_ready),
		.io_connPE_78_valid(_axis_stream_converters_in_78_io_dataOut_TVALID),
		.io_connPE_78_bits(_axis_stream_converters_in_78_io_dataOut_TDATA),
		.io_connPE_79_ready(_argSide_io_connPE_79_ready),
		.io_connPE_79_valid(_axis_stream_converters_in_79_io_dataOut_TVALID),
		.io_connPE_79_bits(_axis_stream_converters_in_79_io_dataOut_TDATA),
		.io_connPE_80_ready(_argSide_io_connPE_80_ready),
		.io_connPE_80_valid(_axis_stream_converters_in_80_io_dataOut_TVALID),
		.io_connPE_80_bits(_axis_stream_converters_in_80_io_dataOut_TDATA),
		.io_connPE_81_ready(_argSide_io_connPE_81_ready),
		.io_connPE_81_valid(_axis_stream_converters_in_81_io_dataOut_TVALID),
		.io_connPE_81_bits(_axis_stream_converters_in_81_io_dataOut_TDATA),
		.io_connPE_82_ready(_argSide_io_connPE_82_ready),
		.io_connPE_82_valid(_axis_stream_converters_in_82_io_dataOut_TVALID),
		.io_connPE_82_bits(_axis_stream_converters_in_82_io_dataOut_TDATA),
		.io_connPE_83_ready(_argSide_io_connPE_83_ready),
		.io_connPE_83_valid(_axis_stream_converters_in_83_io_dataOut_TVALID),
		.io_connPE_83_bits(_axis_stream_converters_in_83_io_dataOut_TDATA),
		.io_connPE_84_ready(_argSide_io_connPE_84_ready),
		.io_connPE_84_valid(_axis_stream_converters_in_84_io_dataOut_TVALID),
		.io_connPE_84_bits(_axis_stream_converters_in_84_io_dataOut_TDATA),
		.io_connPE_85_ready(_argSide_io_connPE_85_ready),
		.io_connPE_85_valid(_axis_stream_converters_in_85_io_dataOut_TVALID),
		.io_connPE_85_bits(_axis_stream_converters_in_85_io_dataOut_TDATA),
		.io_connPE_86_ready(_argSide_io_connPE_86_ready),
		.io_connPE_86_valid(_axis_stream_converters_in_86_io_dataOut_TVALID),
		.io_connPE_86_bits(_axis_stream_converters_in_86_io_dataOut_TDATA),
		.io_connPE_87_ready(_argSide_io_connPE_87_ready),
		.io_connPE_87_valid(_axis_stream_converters_in_87_io_dataOut_TVALID),
		.io_connPE_87_bits(_axis_stream_converters_in_87_io_dataOut_TDATA),
		.io_connPE_88_ready(_argSide_io_connPE_88_ready),
		.io_connPE_88_valid(_axis_stream_converters_in_88_io_dataOut_TVALID),
		.io_connPE_88_bits(_axis_stream_converters_in_88_io_dataOut_TDATA),
		.io_connPE_89_ready(_argSide_io_connPE_89_ready),
		.io_connPE_89_valid(_axis_stream_converters_in_89_io_dataOut_TVALID),
		.io_connPE_89_bits(_axis_stream_converters_in_89_io_dataOut_TDATA),
		.io_connPE_90_ready(_argSide_io_connPE_90_ready),
		.io_connPE_90_valid(_axis_stream_converters_in_90_io_dataOut_TVALID),
		.io_connPE_90_bits(_axis_stream_converters_in_90_io_dataOut_TDATA),
		.io_connPE_91_ready(_argSide_io_connPE_91_ready),
		.io_connPE_91_valid(_axis_stream_converters_in_91_io_dataOut_TVALID),
		.io_connPE_91_bits(_axis_stream_converters_in_91_io_dataOut_TDATA),
		.io_connPE_92_ready(_argSide_io_connPE_92_ready),
		.io_connPE_92_valid(_axis_stream_converters_in_92_io_dataOut_TVALID),
		.io_connPE_92_bits(_axis_stream_converters_in_92_io_dataOut_TDATA),
		.io_connPE_93_ready(_argSide_io_connPE_93_ready),
		.io_connPE_93_valid(_axis_stream_converters_in_93_io_dataOut_TVALID),
		.io_connPE_93_bits(_axis_stream_converters_in_93_io_dataOut_TDATA),
		.io_connPE_94_ready(_argSide_io_connPE_94_ready),
		.io_connPE_94_valid(_axis_stream_converters_in_94_io_dataOut_TVALID),
		.io_connPE_94_bits(_axis_stream_converters_in_94_io_dataOut_TDATA),
		.io_connPE_95_ready(_argSide_io_connPE_95_ready),
		.io_connPE_95_valid(_axis_stream_converters_in_95_io_dataOut_TVALID),
		.io_connPE_95_bits(_axis_stream_converters_in_95_io_dataOut_TDATA),
		.io_connPE_96_ready(_argSide_io_connPE_96_ready),
		.io_connPE_96_valid(_axis_stream_converters_in_96_io_dataOut_TVALID),
		.io_connPE_96_bits(_axis_stream_converters_in_96_io_dataOut_TDATA),
		.io_connPE_97_ready(_argSide_io_connPE_97_ready),
		.io_connPE_97_valid(_axis_stream_converters_in_97_io_dataOut_TVALID),
		.io_connPE_97_bits(_axis_stream_converters_in_97_io_dataOut_TDATA),
		.io_connPE_98_ready(_argSide_io_connPE_98_ready),
		.io_connPE_98_valid(_axis_stream_converters_in_98_io_dataOut_TVALID),
		.io_connPE_98_bits(_axis_stream_converters_in_98_io_dataOut_TDATA),
		.io_connPE_99_ready(_argSide_io_connPE_99_ready),
		.io_connPE_99_valid(_axis_stream_converters_in_99_io_dataOut_TVALID),
		.io_connPE_99_bits(_axis_stream_converters_in_99_io_dataOut_TDATA),
		.io_connPE_100_ready(_argSide_io_connPE_100_ready),
		.io_connPE_100_valid(_axis_stream_converters_in_100_io_dataOut_TVALID),
		.io_connPE_100_bits(_axis_stream_converters_in_100_io_dataOut_TDATA),
		.io_connPE_101_ready(_argSide_io_connPE_101_ready),
		.io_connPE_101_valid(_axis_stream_converters_in_101_io_dataOut_TVALID),
		.io_connPE_101_bits(_axis_stream_converters_in_101_io_dataOut_TDATA),
		.io_connPE_102_ready(_argSide_io_connPE_102_ready),
		.io_connPE_102_valid(_axis_stream_converters_in_102_io_dataOut_TVALID),
		.io_connPE_102_bits(_axis_stream_converters_in_102_io_dataOut_TDATA),
		.io_connPE_103_ready(_argSide_io_connPE_103_ready),
		.io_connPE_103_valid(_axis_stream_converters_in_103_io_dataOut_TVALID),
		.io_connPE_103_bits(_axis_stream_converters_in_103_io_dataOut_TDATA),
		.io_connPE_104_ready(_argSide_io_connPE_104_ready),
		.io_connPE_104_valid(_axis_stream_converters_in_104_io_dataOut_TVALID),
		.io_connPE_104_bits(_axis_stream_converters_in_104_io_dataOut_TDATA),
		.io_connPE_105_ready(_argSide_io_connPE_105_ready),
		.io_connPE_105_valid(_axis_stream_converters_in_105_io_dataOut_TVALID),
		.io_connPE_105_bits(_axis_stream_converters_in_105_io_dataOut_TDATA),
		.io_connPE_106_ready(_argSide_io_connPE_106_ready),
		.io_connPE_106_valid(_axis_stream_converters_in_106_io_dataOut_TVALID),
		.io_connPE_106_bits(_axis_stream_converters_in_106_io_dataOut_TDATA),
		.io_connPE_107_ready(_argSide_io_connPE_107_ready),
		.io_connPE_107_valid(_axis_stream_converters_in_107_io_dataOut_TVALID),
		.io_connPE_107_bits(_axis_stream_converters_in_107_io_dataOut_TDATA),
		.io_connPE_108_ready(_argSide_io_connPE_108_ready),
		.io_connPE_108_valid(_axis_stream_converters_in_108_io_dataOut_TVALID),
		.io_connPE_108_bits(_axis_stream_converters_in_108_io_dataOut_TDATA),
		.io_connPE_109_ready(_argSide_io_connPE_109_ready),
		.io_connPE_109_valid(_axis_stream_converters_in_109_io_dataOut_TVALID),
		.io_connPE_109_bits(_axis_stream_converters_in_109_io_dataOut_TDATA),
		.io_connPE_110_ready(_argSide_io_connPE_110_ready),
		.io_connPE_110_valid(_axis_stream_converters_in_110_io_dataOut_TVALID),
		.io_connPE_110_bits(_axis_stream_converters_in_110_io_dataOut_TDATA),
		.io_connPE_111_ready(_argSide_io_connPE_111_ready),
		.io_connPE_111_valid(_axis_stream_converters_in_111_io_dataOut_TVALID),
		.io_connPE_111_bits(_axis_stream_converters_in_111_io_dataOut_TDATA),
		.io_connPE_112_ready(_argSide_io_connPE_112_ready),
		.io_connPE_112_valid(_axis_stream_converters_in_112_io_dataOut_TVALID),
		.io_connPE_112_bits(_axis_stream_converters_in_112_io_dataOut_TDATA),
		.io_connPE_113_ready(_argSide_io_connPE_113_ready),
		.io_connPE_113_valid(_axis_stream_converters_in_113_io_dataOut_TVALID),
		.io_connPE_113_bits(_axis_stream_converters_in_113_io_dataOut_TDATA),
		.io_connPE_114_ready(_argSide_io_connPE_114_ready),
		.io_connPE_114_valid(_axis_stream_converters_in_114_io_dataOut_TVALID),
		.io_connPE_114_bits(_axis_stream_converters_in_114_io_dataOut_TDATA),
		.io_connPE_115_ready(_argSide_io_connPE_115_ready),
		.io_connPE_115_valid(_axis_stream_converters_in_115_io_dataOut_TVALID),
		.io_connPE_115_bits(_axis_stream_converters_in_115_io_dataOut_TDATA),
		.io_connPE_116_ready(_argSide_io_connPE_116_ready),
		.io_connPE_116_valid(_axis_stream_converters_in_116_io_dataOut_TVALID),
		.io_connPE_116_bits(_axis_stream_converters_in_116_io_dataOut_TDATA),
		.io_connPE_117_ready(_argSide_io_connPE_117_ready),
		.io_connPE_117_valid(_axis_stream_converters_in_117_io_dataOut_TVALID),
		.io_connPE_117_bits(_axis_stream_converters_in_117_io_dataOut_TDATA),
		.io_connPE_118_ready(_argSide_io_connPE_118_ready),
		.io_connPE_118_valid(_axis_stream_converters_in_118_io_dataOut_TVALID),
		.io_connPE_118_bits(_axis_stream_converters_in_118_io_dataOut_TDATA),
		.io_connPE_119_ready(_argSide_io_connPE_119_ready),
		.io_connPE_119_valid(_axis_stream_converters_in_119_io_dataOut_TVALID),
		.io_connPE_119_bits(_axis_stream_converters_in_119_io_dataOut_TDATA),
		.io_connPE_120_ready(_argSide_io_connPE_120_ready),
		.io_connPE_120_valid(_axis_stream_converters_in_120_io_dataOut_TVALID),
		.io_connPE_120_bits(_axis_stream_converters_in_120_io_dataOut_TDATA),
		.io_connPE_121_ready(_argSide_io_connPE_121_ready),
		.io_connPE_121_valid(_axis_stream_converters_in_121_io_dataOut_TVALID),
		.io_connPE_121_bits(_axis_stream_converters_in_121_io_dataOut_TDATA),
		.io_connPE_122_ready(_argSide_io_connPE_122_ready),
		.io_connPE_122_valid(_axis_stream_converters_in_122_io_dataOut_TVALID),
		.io_connPE_122_bits(_axis_stream_converters_in_122_io_dataOut_TDATA),
		.io_connPE_123_ready(_argSide_io_connPE_123_ready),
		.io_connPE_123_valid(_axis_stream_converters_in_123_io_dataOut_TVALID),
		.io_connPE_123_bits(_axis_stream_converters_in_123_io_dataOut_TDATA),
		.io_connPE_124_ready(_argSide_io_connPE_124_ready),
		.io_connPE_124_valid(_axis_stream_converters_in_124_io_dataOut_TVALID),
		.io_connPE_124_bits(_axis_stream_converters_in_124_io_dataOut_TDATA),
		.io_connPE_125_ready(_argSide_io_connPE_125_ready),
		.io_connPE_125_valid(_axis_stream_converters_in_125_io_dataOut_TVALID),
		.io_connPE_125_bits(_axis_stream_converters_in_125_io_dataOut_TDATA),
		.io_connPE_126_ready(_argSide_io_connPE_126_ready),
		.io_connPE_126_valid(_axis_stream_converters_in_126_io_dataOut_TVALID),
		.io_connPE_126_bits(_axis_stream_converters_in_126_io_dataOut_TDATA),
		.io_connPE_127_ready(_argSide_io_connPE_127_ready),
		.io_connPE_127_valid(_axis_stream_converters_in_127_io_dataOut_TVALID),
		.io_connPE_127_bits(_axis_stream_converters_in_127_io_dataOut_TDATA)
	);
	ArgumentServer argRouteServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_0_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_0_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_0_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_0_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_0_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_0_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_0_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_0_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_0_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_0_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_0_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_0_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_0_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_0_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_0_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_0_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_0_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_0_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_0_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_0_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_0_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_0_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_0_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_0_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_0_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_0_io_read_data_bits)
	);
	ArgumentServer argRouteServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_1_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_1_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_1_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_1_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_1_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_1_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_1_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_1_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_1_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_1_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_1_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_1_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_1_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_1_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_1_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_1_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_1_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_1_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_1_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_1_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_1_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_1_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_1_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_1_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_1_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_1_io_read_data_bits)
	);
	ArgumentServer argRouteServers_2(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_2_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_2_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_2_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_2_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_2_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_2_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_2_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_2_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_2_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_2_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_2_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_2_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_2_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_2_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_2_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_2_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_2_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_2_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_2_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_2_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_2_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_2_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_2_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_2_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_2_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_2_io_read_data_bits)
	);
	ArgumentServer argRouteServers_3(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_3_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_3_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_3_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_3_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_3_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_3_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_3_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_3_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_3_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_3_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_3_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_3_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_3_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_3_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_3_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_3_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_3_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_3_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_3_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_3_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_3_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_3_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_3_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_3_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_3_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_3_io_read_data_bits)
	);
	ArgumentServer argRouteServers_4(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_4_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_4_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_4_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_4_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_4_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_4_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_4_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_4_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_4_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_4_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_4_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_4_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_4_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_4_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_4_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_4_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_4_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_4_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_4_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_4_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_4_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_4_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_4_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_4_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_4_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_4_io_read_data_bits)
	);
	ArgumentServer argRouteServers_5(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_5_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_5_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_5_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_5_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_5_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_5_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_5_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_5_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_5_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_5_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_5_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_5_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_5_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_5_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_5_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_5_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_5_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_5_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_5_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_5_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_5_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_5_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_5_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_5_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_5_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_5_io_read_data_bits)
	);
	ArgumentServer argRouteServers_6(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_6_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_6_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_6_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_6_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_6_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_6_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_6_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_6_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_6_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_6_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_6_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_6_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_6_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_6_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_6_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_6_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_6_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_6_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_6_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_6_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_6_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_6_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_6_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_6_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_6_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_6_io_read_data_bits)
	);
	ArgumentServer argRouteServers_7(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_7_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_7_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_7_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_7_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_7_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_7_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_7_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_7_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_7_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_7_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_7_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_7_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_7_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_7_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_7_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_7_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_7_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_7_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_7_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_7_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_7_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_7_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_7_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_7_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_7_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_7_io_read_data_bits)
	);
	ArgumentServer argRouteServers_8(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_8_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_8_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_8_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_8_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_8_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_8_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_8_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_8_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_8_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_8_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_8_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_8_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_8_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_8_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_8_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_8_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_8_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_8_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_8_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_8_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_8_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_8_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_8_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_8_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_8_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_8_io_read_data_bits)
	);
	ArgumentServer argRouteServers_9(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_9_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_9_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_9_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_9_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_9_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_9_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_9_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_9_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_9_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_9_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_9_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_9_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_9_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_9_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_9_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_9_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_9_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_9_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_9_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_9_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_9_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_9_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_9_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_9_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_9_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_9_io_read_data_bits)
	);
	ArgumentServer argRouteServers_10(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_10_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_10_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_10_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_10_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_10_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_10_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_10_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_10_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_10_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_10_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_10_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_10_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_10_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_10_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_10_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_10_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_10_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_10_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_10_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_10_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_10_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_10_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_10_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_10_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_10_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_10_io_read_data_bits)
	);
	ArgumentServer argRouteServers_11(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_11_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_11_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_11_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_11_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_11_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_11_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_11_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_11_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_11_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_11_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_11_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_11_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_11_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_11_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_11_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_11_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_11_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_11_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_11_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_11_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_11_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_11_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_11_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_11_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_11_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_11_io_read_data_bits)
	);
	ArgumentServer argRouteServers_12(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_12_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_12_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_12_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_12_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_12_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_12_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_12_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_12_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_12_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_12_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_12_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_12_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_12_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_12_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_12_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_12_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_12_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_12_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_12_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_12_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_12_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_12_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_12_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_12_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_12_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_12_io_read_data_bits)
	);
	ArgumentServer argRouteServers_13(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_13_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_13_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_13_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_13_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_13_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_13_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_13_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_13_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_13_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_13_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_13_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_13_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_13_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_13_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_13_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_13_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_13_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_13_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_13_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_13_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_13_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_13_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_13_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_13_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_13_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_13_io_read_data_bits)
	);
	ArgumentServer argRouteServers_14(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_14_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_14_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_14_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_14_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_14_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_14_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_14_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_14_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_14_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_14_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_14_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_14_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_14_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_14_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_14_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_14_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_14_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_14_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_14_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_14_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_14_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_14_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_14_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_14_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_14_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_14_io_read_data_bits)
	);
	ArgumentServer argRouteServers_15(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_15_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_15_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_15_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_15_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_15_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_15_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_15_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_15_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_15_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_15_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_15_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_15_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_15_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_15_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_15_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_15_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_15_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_15_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_15_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_15_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_15_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_15_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_15_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_15_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_15_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_15_io_read_data_bits)
	);
	RVtoAXIBridge_8 argRouteRvm_0(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_0_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_0_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_0_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_0_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_0_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_0_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_0_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_0_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_0_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_0_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_0_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_0_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_0_ar_ready),
		.axi_ar_valid(_argRouteRvm_0_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_0_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_0_axi_r_ready),
		.axi_r_valid(_mux_s_axi_0_r_valid),
		.axi_r_bits_data(_mux_s_axi_0_r_bits_data),
		.axi_aw_ready(_mux_s_axi_0_aw_ready),
		.axi_aw_valid(_argRouteRvm_0_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_0_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_0_w_ready),
		.axi_w_valid(_argRouteRvm_0_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_0_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_0_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_1(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_1_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_1_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_1_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_1_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_1_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_1_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_1_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_1_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_1_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_1_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_1_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_1_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_1_ar_ready),
		.axi_ar_valid(_argRouteRvm_1_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_1_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_1_axi_r_ready),
		.axi_r_valid(_mux_s_axi_1_r_valid),
		.axi_r_bits_data(_mux_s_axi_1_r_bits_data),
		.axi_aw_ready(_mux_s_axi_1_aw_ready),
		.axi_aw_valid(_argRouteRvm_1_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_1_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_1_w_ready),
		.axi_w_valid(_argRouteRvm_1_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_1_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_1_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_2(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_2_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_2_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_2_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_2_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_2_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_2_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_2_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_2_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_2_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_2_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_2_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_2_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_2_ar_ready),
		.axi_ar_valid(_argRouteRvm_2_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_2_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_2_axi_r_ready),
		.axi_r_valid(_mux_s_axi_2_r_valid),
		.axi_r_bits_data(_mux_s_axi_2_r_bits_data),
		.axi_aw_ready(_mux_s_axi_2_aw_ready),
		.axi_aw_valid(_argRouteRvm_2_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_2_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_2_w_ready),
		.axi_w_valid(_argRouteRvm_2_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_2_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_2_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_3(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_3_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_3_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_3_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_3_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_3_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_3_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_3_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_3_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_3_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_3_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_3_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_3_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_3_ar_ready),
		.axi_ar_valid(_argRouteRvm_3_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_3_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_3_axi_r_ready),
		.axi_r_valid(_mux_s_axi_3_r_valid),
		.axi_r_bits_data(_mux_s_axi_3_r_bits_data),
		.axi_aw_ready(_mux_s_axi_3_aw_ready),
		.axi_aw_valid(_argRouteRvm_3_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_3_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_3_w_ready),
		.axi_w_valid(_argRouteRvm_3_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_3_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_3_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_4(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_4_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_4_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_4_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_4_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_4_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_4_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_4_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_4_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_4_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_4_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_4_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_4_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_4_ar_ready),
		.axi_ar_valid(_argRouteRvm_4_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_4_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_4_axi_r_ready),
		.axi_r_valid(_mux_s_axi_4_r_valid),
		.axi_r_bits_data(_mux_s_axi_4_r_bits_data),
		.axi_aw_ready(_mux_s_axi_4_aw_ready),
		.axi_aw_valid(_argRouteRvm_4_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_4_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_4_w_ready),
		.axi_w_valid(_argRouteRvm_4_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_4_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_4_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_5(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_5_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_5_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_5_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_5_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_5_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_5_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_5_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_5_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_5_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_5_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_5_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_5_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_5_ar_ready),
		.axi_ar_valid(_argRouteRvm_5_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_5_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_5_axi_r_ready),
		.axi_r_valid(_mux_s_axi_5_r_valid),
		.axi_r_bits_data(_mux_s_axi_5_r_bits_data),
		.axi_aw_ready(_mux_s_axi_5_aw_ready),
		.axi_aw_valid(_argRouteRvm_5_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_5_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_5_w_ready),
		.axi_w_valid(_argRouteRvm_5_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_5_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_5_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_6(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_6_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_6_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_6_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_6_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_6_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_6_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_6_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_6_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_6_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_6_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_6_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_6_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_6_ar_ready),
		.axi_ar_valid(_argRouteRvm_6_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_6_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_6_axi_r_ready),
		.axi_r_valid(_mux_s_axi_6_r_valid),
		.axi_r_bits_data(_mux_s_axi_6_r_bits_data),
		.axi_aw_ready(_mux_s_axi_6_aw_ready),
		.axi_aw_valid(_argRouteRvm_6_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_6_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_6_w_ready),
		.axi_w_valid(_argRouteRvm_6_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_6_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_6_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_7(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_7_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_7_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_7_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_7_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_7_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_7_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_7_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_7_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_7_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_7_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_7_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_7_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_7_ar_ready),
		.axi_ar_valid(_argRouteRvm_7_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_7_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_7_axi_r_ready),
		.axi_r_valid(_mux_s_axi_7_r_valid),
		.axi_r_bits_data(_mux_s_axi_7_r_bits_data),
		.axi_aw_ready(_mux_s_axi_7_aw_ready),
		.axi_aw_valid(_argRouteRvm_7_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_7_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_7_w_ready),
		.axi_w_valid(_argRouteRvm_7_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_7_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_7_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_8(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_8_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_8_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_8_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_8_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_8_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_8_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_8_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_8_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_8_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_8_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_8_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_8_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_8_ar_ready),
		.axi_ar_valid(_argRouteRvm_8_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_8_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_8_axi_r_ready),
		.axi_r_valid(_mux_s_axi_8_r_valid),
		.axi_r_bits_data(_mux_s_axi_8_r_bits_data),
		.axi_aw_ready(_mux_s_axi_8_aw_ready),
		.axi_aw_valid(_argRouteRvm_8_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_8_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_8_w_ready),
		.axi_w_valid(_argRouteRvm_8_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_8_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_8_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_9(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_9_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_9_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_9_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_9_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_9_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_9_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_9_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_9_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_9_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_9_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_9_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_9_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_9_ar_ready),
		.axi_ar_valid(_argRouteRvm_9_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_9_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_9_axi_r_ready),
		.axi_r_valid(_mux_s_axi_9_r_valid),
		.axi_r_bits_data(_mux_s_axi_9_r_bits_data),
		.axi_aw_ready(_mux_s_axi_9_aw_ready),
		.axi_aw_valid(_argRouteRvm_9_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_9_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_9_w_ready),
		.axi_w_valid(_argRouteRvm_9_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_9_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_9_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_10(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_10_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_10_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_10_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_10_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_10_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_10_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_10_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_10_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_10_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_10_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_10_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_10_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_10_ar_ready),
		.axi_ar_valid(_argRouteRvm_10_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_10_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_10_axi_r_ready),
		.axi_r_valid(_mux_s_axi_10_r_valid),
		.axi_r_bits_data(_mux_s_axi_10_r_bits_data),
		.axi_aw_ready(_mux_s_axi_10_aw_ready),
		.axi_aw_valid(_argRouteRvm_10_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_10_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_10_w_ready),
		.axi_w_valid(_argRouteRvm_10_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_10_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_10_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_11(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_11_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_11_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_11_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_11_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_11_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_11_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_11_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_11_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_11_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_11_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_11_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_11_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_11_ar_ready),
		.axi_ar_valid(_argRouteRvm_11_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_11_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_11_axi_r_ready),
		.axi_r_valid(_mux_s_axi_11_r_valid),
		.axi_r_bits_data(_mux_s_axi_11_r_bits_data),
		.axi_aw_ready(_mux_s_axi_11_aw_ready),
		.axi_aw_valid(_argRouteRvm_11_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_11_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_11_w_ready),
		.axi_w_valid(_argRouteRvm_11_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_11_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_11_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_12(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_12_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_12_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_12_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_12_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_12_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_12_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_12_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_12_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_12_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_12_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_12_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_12_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_12_ar_ready),
		.axi_ar_valid(_argRouteRvm_12_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_12_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_12_axi_r_ready),
		.axi_r_valid(_mux_s_axi_12_r_valid),
		.axi_r_bits_data(_mux_s_axi_12_r_bits_data),
		.axi_aw_ready(_mux_s_axi_12_aw_ready),
		.axi_aw_valid(_argRouteRvm_12_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_12_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_12_w_ready),
		.axi_w_valid(_argRouteRvm_12_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_12_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_12_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_13(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_13_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_13_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_13_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_13_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_13_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_13_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_13_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_13_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_13_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_13_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_13_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_13_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_13_ar_ready),
		.axi_ar_valid(_argRouteRvm_13_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_13_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_13_axi_r_ready),
		.axi_r_valid(_mux_s_axi_13_r_valid),
		.axi_r_bits_data(_mux_s_axi_13_r_bits_data),
		.axi_aw_ready(_mux_s_axi_13_aw_ready),
		.axi_aw_valid(_argRouteRvm_13_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_13_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_13_w_ready),
		.axi_w_valid(_argRouteRvm_13_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_13_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_13_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_14(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_14_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_14_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_14_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_14_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_14_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_14_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_14_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_14_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_14_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_14_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_14_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_14_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_14_ar_ready),
		.axi_ar_valid(_argRouteRvm_14_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_14_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_14_axi_r_ready),
		.axi_r_valid(_mux_s_axi_14_r_valid),
		.axi_r_bits_data(_mux_s_axi_14_r_bits_data),
		.axi_aw_ready(_mux_s_axi_14_aw_ready),
		.axi_aw_valid(_argRouteRvm_14_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_14_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_14_w_ready),
		.axi_w_valid(_argRouteRvm_14_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_14_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_14_b_valid)
	);
	RVtoAXIBridge_8 argRouteRvm_15(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_15_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_15_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_15_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_15_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_15_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_15_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_15_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_15_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_15_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_15_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_15_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_15_io_write_data_bits),
		.axi_ar_ready(_mux_s_axi_15_ar_ready),
		.axi_ar_valid(_argRouteRvm_15_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvm_15_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvm_15_axi_r_ready),
		.axi_r_valid(_mux_s_axi_15_r_valid),
		.axi_r_bits_data(_mux_s_axi_15_r_bits_data),
		.axi_aw_ready(_mux_s_axi_15_aw_ready),
		.axi_aw_valid(_argRouteRvm_15_axi_aw_valid),
		.axi_aw_bits_addr(_argRouteRvm_15_axi_aw_bits_addr),
		.axi_w_ready(_mux_s_axi_15_w_ready),
		.axi_w_valid(_argRouteRvm_15_axi_w_valid),
		.axi_w_bits_data(_argRouteRvm_15_axi_w_bits_data),
		.axi_b_valid(_mux_s_axi_15_b_valid)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_0(
		.io_read_address_ready(_argRouteRvmReadOnly_0_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_0_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_0_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_0_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_0_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_0_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_16_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_0_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_0_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_0_axi_r_ready),
		.axi_r_valid(_mux_s_axi_16_r_valid),
		.axi_r_bits_data(_mux_s_axi_16_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_1(
		.io_read_address_ready(_argRouteRvmReadOnly_1_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_1_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_1_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_1_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_1_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_1_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_17_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_1_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_1_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_1_axi_r_ready),
		.axi_r_valid(_mux_s_axi_17_r_valid),
		.axi_r_bits_data(_mux_s_axi_17_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_2(
		.io_read_address_ready(_argRouteRvmReadOnly_2_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_2_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_2_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_2_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_2_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_2_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_18_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_2_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_2_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_2_axi_r_ready),
		.axi_r_valid(_mux_s_axi_18_r_valid),
		.axi_r_bits_data(_mux_s_axi_18_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_3(
		.io_read_address_ready(_argRouteRvmReadOnly_3_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_3_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_3_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_3_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_3_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_3_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_19_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_3_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_3_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_3_axi_r_ready),
		.axi_r_valid(_mux_s_axi_19_r_valid),
		.axi_r_bits_data(_mux_s_axi_19_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_4(
		.io_read_address_ready(_argRouteRvmReadOnly_4_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_4_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_4_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_4_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_4_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_4_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_20_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_4_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_4_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_4_axi_r_ready),
		.axi_r_valid(_mux_s_axi_20_r_valid),
		.axi_r_bits_data(_mux_s_axi_20_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_5(
		.io_read_address_ready(_argRouteRvmReadOnly_5_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_5_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_5_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_5_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_5_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_5_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_21_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_5_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_5_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_5_axi_r_ready),
		.axi_r_valid(_mux_s_axi_21_r_valid),
		.axi_r_bits_data(_mux_s_axi_21_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_6(
		.io_read_address_ready(_argRouteRvmReadOnly_6_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_6_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_6_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_6_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_6_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_6_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_22_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_6_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_6_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_6_axi_r_ready),
		.axi_r_valid(_mux_s_axi_22_r_valid),
		.axi_r_bits_data(_mux_s_axi_22_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_7(
		.io_read_address_ready(_argRouteRvmReadOnly_7_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_7_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_7_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_7_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_7_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_7_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_23_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_7_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_7_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_7_axi_r_ready),
		.axi_r_valid(_mux_s_axi_23_r_valid),
		.axi_r_bits_data(_mux_s_axi_23_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_8(
		.io_read_address_ready(_argRouteRvmReadOnly_8_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_8_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_8_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_8_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_8_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_8_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_24_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_8_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_8_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_8_axi_r_ready),
		.axi_r_valid(_mux_s_axi_24_r_valid),
		.axi_r_bits_data(_mux_s_axi_24_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_9(
		.io_read_address_ready(_argRouteRvmReadOnly_9_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_9_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_9_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_9_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_9_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_9_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_25_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_9_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_9_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_9_axi_r_ready),
		.axi_r_valid(_mux_s_axi_25_r_valid),
		.axi_r_bits_data(_mux_s_axi_25_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_10(
		.io_read_address_ready(_argRouteRvmReadOnly_10_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_10_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_10_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_10_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_10_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_10_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_26_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_10_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_10_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_10_axi_r_ready),
		.axi_r_valid(_mux_s_axi_26_r_valid),
		.axi_r_bits_data(_mux_s_axi_26_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_11(
		.io_read_address_ready(_argRouteRvmReadOnly_11_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_11_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_11_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_11_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_11_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_11_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_27_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_11_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_11_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_11_axi_r_ready),
		.axi_r_valid(_mux_s_axi_27_r_valid),
		.axi_r_bits_data(_mux_s_axi_27_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_12(
		.io_read_address_ready(_argRouteRvmReadOnly_12_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_12_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_12_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_12_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_12_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_12_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_28_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_12_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_12_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_12_axi_r_ready),
		.axi_r_valid(_mux_s_axi_28_r_valid),
		.axi_r_bits_data(_mux_s_axi_28_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_13(
		.io_read_address_ready(_argRouteRvmReadOnly_13_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_13_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_13_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_13_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_13_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_13_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_29_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_13_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_13_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_13_axi_r_ready),
		.axi_r_valid(_mux_s_axi_29_r_valid),
		.axi_r_bits_data(_mux_s_axi_29_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_14(
		.io_read_address_ready(_argRouteRvmReadOnly_14_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_14_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_14_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_14_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_14_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_14_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_30_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_14_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_14_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_14_axi_r_ready),
		.axi_r_valid(_mux_s_axi_30_r_valid),
		.axi_r_bits_data(_mux_s_axi_30_r_bits_data)
	);
	RVtoAXIBridge_24 argRouteRvmReadOnly_15(
		.io_read_address_ready(_argRouteRvmReadOnly_15_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_15_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_15_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_15_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_15_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_15_io_read_data_bits),
		.axi_ar_ready(_mux_s_axi_31_ar_ready),
		.axi_ar_valid(_argRouteRvmReadOnly_15_axi_ar_valid),
		.axi_ar_bits_addr(_argRouteRvmReadOnly_15_axi_ar_bits_addr),
		.axi_r_ready(_argRouteRvmReadOnly_15_axi_r_ready),
		.axi_r_valid(_mux_s_axi_31_r_valid),
		.axi_r_bits_data(_mux_s_axi_31_r_bits_data)
	);
	axi4FullMux_3 mux(
		.clock(clock),
		.reset(reset),
		.s_axi_0_ar_ready(_mux_s_axi_0_ar_ready),
		.s_axi_0_ar_valid(_argRouteRvm_0_axi_ar_valid),
		.s_axi_0_ar_bits_addr(_argRouteRvm_0_axi_ar_bits_addr),
		.s_axi_0_r_ready(_argRouteRvm_0_axi_r_ready),
		.s_axi_0_r_valid(_mux_s_axi_0_r_valid),
		.s_axi_0_r_bits_data(_mux_s_axi_0_r_bits_data),
		.s_axi_0_aw_ready(_mux_s_axi_0_aw_ready),
		.s_axi_0_aw_valid(_argRouteRvm_0_axi_aw_valid),
		.s_axi_0_aw_bits_addr(_argRouteRvm_0_axi_aw_bits_addr),
		.s_axi_0_w_ready(_mux_s_axi_0_w_ready),
		.s_axi_0_w_valid(_argRouteRvm_0_axi_w_valid),
		.s_axi_0_w_bits_data(_argRouteRvm_0_axi_w_bits_data),
		.s_axi_0_b_valid(_mux_s_axi_0_b_valid),
		.s_axi_1_ar_ready(_mux_s_axi_1_ar_ready),
		.s_axi_1_ar_valid(_argRouteRvm_1_axi_ar_valid),
		.s_axi_1_ar_bits_addr(_argRouteRvm_1_axi_ar_bits_addr),
		.s_axi_1_r_ready(_argRouteRvm_1_axi_r_ready),
		.s_axi_1_r_valid(_mux_s_axi_1_r_valid),
		.s_axi_1_r_bits_data(_mux_s_axi_1_r_bits_data),
		.s_axi_1_aw_ready(_mux_s_axi_1_aw_ready),
		.s_axi_1_aw_valid(_argRouteRvm_1_axi_aw_valid),
		.s_axi_1_aw_bits_addr(_argRouteRvm_1_axi_aw_bits_addr),
		.s_axi_1_w_ready(_mux_s_axi_1_w_ready),
		.s_axi_1_w_valid(_argRouteRvm_1_axi_w_valid),
		.s_axi_1_w_bits_data(_argRouteRvm_1_axi_w_bits_data),
		.s_axi_1_b_valid(_mux_s_axi_1_b_valid),
		.s_axi_2_ar_ready(_mux_s_axi_2_ar_ready),
		.s_axi_2_ar_valid(_argRouteRvm_2_axi_ar_valid),
		.s_axi_2_ar_bits_addr(_argRouteRvm_2_axi_ar_bits_addr),
		.s_axi_2_r_ready(_argRouteRvm_2_axi_r_ready),
		.s_axi_2_r_valid(_mux_s_axi_2_r_valid),
		.s_axi_2_r_bits_data(_mux_s_axi_2_r_bits_data),
		.s_axi_2_aw_ready(_mux_s_axi_2_aw_ready),
		.s_axi_2_aw_valid(_argRouteRvm_2_axi_aw_valid),
		.s_axi_2_aw_bits_addr(_argRouteRvm_2_axi_aw_bits_addr),
		.s_axi_2_w_ready(_mux_s_axi_2_w_ready),
		.s_axi_2_w_valid(_argRouteRvm_2_axi_w_valid),
		.s_axi_2_w_bits_data(_argRouteRvm_2_axi_w_bits_data),
		.s_axi_2_b_valid(_mux_s_axi_2_b_valid),
		.s_axi_3_ar_ready(_mux_s_axi_3_ar_ready),
		.s_axi_3_ar_valid(_argRouteRvm_3_axi_ar_valid),
		.s_axi_3_ar_bits_addr(_argRouteRvm_3_axi_ar_bits_addr),
		.s_axi_3_r_ready(_argRouteRvm_3_axi_r_ready),
		.s_axi_3_r_valid(_mux_s_axi_3_r_valid),
		.s_axi_3_r_bits_data(_mux_s_axi_3_r_bits_data),
		.s_axi_3_aw_ready(_mux_s_axi_3_aw_ready),
		.s_axi_3_aw_valid(_argRouteRvm_3_axi_aw_valid),
		.s_axi_3_aw_bits_addr(_argRouteRvm_3_axi_aw_bits_addr),
		.s_axi_3_w_ready(_mux_s_axi_3_w_ready),
		.s_axi_3_w_valid(_argRouteRvm_3_axi_w_valid),
		.s_axi_3_w_bits_data(_argRouteRvm_3_axi_w_bits_data),
		.s_axi_3_b_valid(_mux_s_axi_3_b_valid),
		.s_axi_4_ar_ready(_mux_s_axi_4_ar_ready),
		.s_axi_4_ar_valid(_argRouteRvm_4_axi_ar_valid),
		.s_axi_4_ar_bits_addr(_argRouteRvm_4_axi_ar_bits_addr),
		.s_axi_4_r_ready(_argRouteRvm_4_axi_r_ready),
		.s_axi_4_r_valid(_mux_s_axi_4_r_valid),
		.s_axi_4_r_bits_data(_mux_s_axi_4_r_bits_data),
		.s_axi_4_aw_ready(_mux_s_axi_4_aw_ready),
		.s_axi_4_aw_valid(_argRouteRvm_4_axi_aw_valid),
		.s_axi_4_aw_bits_addr(_argRouteRvm_4_axi_aw_bits_addr),
		.s_axi_4_w_ready(_mux_s_axi_4_w_ready),
		.s_axi_4_w_valid(_argRouteRvm_4_axi_w_valid),
		.s_axi_4_w_bits_data(_argRouteRvm_4_axi_w_bits_data),
		.s_axi_4_b_valid(_mux_s_axi_4_b_valid),
		.s_axi_5_ar_ready(_mux_s_axi_5_ar_ready),
		.s_axi_5_ar_valid(_argRouteRvm_5_axi_ar_valid),
		.s_axi_5_ar_bits_addr(_argRouteRvm_5_axi_ar_bits_addr),
		.s_axi_5_r_ready(_argRouteRvm_5_axi_r_ready),
		.s_axi_5_r_valid(_mux_s_axi_5_r_valid),
		.s_axi_5_r_bits_data(_mux_s_axi_5_r_bits_data),
		.s_axi_5_aw_ready(_mux_s_axi_5_aw_ready),
		.s_axi_5_aw_valid(_argRouteRvm_5_axi_aw_valid),
		.s_axi_5_aw_bits_addr(_argRouteRvm_5_axi_aw_bits_addr),
		.s_axi_5_w_ready(_mux_s_axi_5_w_ready),
		.s_axi_5_w_valid(_argRouteRvm_5_axi_w_valid),
		.s_axi_5_w_bits_data(_argRouteRvm_5_axi_w_bits_data),
		.s_axi_5_b_valid(_mux_s_axi_5_b_valid),
		.s_axi_6_ar_ready(_mux_s_axi_6_ar_ready),
		.s_axi_6_ar_valid(_argRouteRvm_6_axi_ar_valid),
		.s_axi_6_ar_bits_addr(_argRouteRvm_6_axi_ar_bits_addr),
		.s_axi_6_r_ready(_argRouteRvm_6_axi_r_ready),
		.s_axi_6_r_valid(_mux_s_axi_6_r_valid),
		.s_axi_6_r_bits_data(_mux_s_axi_6_r_bits_data),
		.s_axi_6_aw_ready(_mux_s_axi_6_aw_ready),
		.s_axi_6_aw_valid(_argRouteRvm_6_axi_aw_valid),
		.s_axi_6_aw_bits_addr(_argRouteRvm_6_axi_aw_bits_addr),
		.s_axi_6_w_ready(_mux_s_axi_6_w_ready),
		.s_axi_6_w_valid(_argRouteRvm_6_axi_w_valid),
		.s_axi_6_w_bits_data(_argRouteRvm_6_axi_w_bits_data),
		.s_axi_6_b_valid(_mux_s_axi_6_b_valid),
		.s_axi_7_ar_ready(_mux_s_axi_7_ar_ready),
		.s_axi_7_ar_valid(_argRouteRvm_7_axi_ar_valid),
		.s_axi_7_ar_bits_addr(_argRouteRvm_7_axi_ar_bits_addr),
		.s_axi_7_r_ready(_argRouteRvm_7_axi_r_ready),
		.s_axi_7_r_valid(_mux_s_axi_7_r_valid),
		.s_axi_7_r_bits_data(_mux_s_axi_7_r_bits_data),
		.s_axi_7_aw_ready(_mux_s_axi_7_aw_ready),
		.s_axi_7_aw_valid(_argRouteRvm_7_axi_aw_valid),
		.s_axi_7_aw_bits_addr(_argRouteRvm_7_axi_aw_bits_addr),
		.s_axi_7_w_ready(_mux_s_axi_7_w_ready),
		.s_axi_7_w_valid(_argRouteRvm_7_axi_w_valid),
		.s_axi_7_w_bits_data(_argRouteRvm_7_axi_w_bits_data),
		.s_axi_7_b_valid(_mux_s_axi_7_b_valid),
		.s_axi_8_ar_ready(_mux_s_axi_8_ar_ready),
		.s_axi_8_ar_valid(_argRouteRvm_8_axi_ar_valid),
		.s_axi_8_ar_bits_addr(_argRouteRvm_8_axi_ar_bits_addr),
		.s_axi_8_r_ready(_argRouteRvm_8_axi_r_ready),
		.s_axi_8_r_valid(_mux_s_axi_8_r_valid),
		.s_axi_8_r_bits_data(_mux_s_axi_8_r_bits_data),
		.s_axi_8_aw_ready(_mux_s_axi_8_aw_ready),
		.s_axi_8_aw_valid(_argRouteRvm_8_axi_aw_valid),
		.s_axi_8_aw_bits_addr(_argRouteRvm_8_axi_aw_bits_addr),
		.s_axi_8_w_ready(_mux_s_axi_8_w_ready),
		.s_axi_8_w_valid(_argRouteRvm_8_axi_w_valid),
		.s_axi_8_w_bits_data(_argRouteRvm_8_axi_w_bits_data),
		.s_axi_8_b_valid(_mux_s_axi_8_b_valid),
		.s_axi_9_ar_ready(_mux_s_axi_9_ar_ready),
		.s_axi_9_ar_valid(_argRouteRvm_9_axi_ar_valid),
		.s_axi_9_ar_bits_addr(_argRouteRvm_9_axi_ar_bits_addr),
		.s_axi_9_r_ready(_argRouteRvm_9_axi_r_ready),
		.s_axi_9_r_valid(_mux_s_axi_9_r_valid),
		.s_axi_9_r_bits_data(_mux_s_axi_9_r_bits_data),
		.s_axi_9_aw_ready(_mux_s_axi_9_aw_ready),
		.s_axi_9_aw_valid(_argRouteRvm_9_axi_aw_valid),
		.s_axi_9_aw_bits_addr(_argRouteRvm_9_axi_aw_bits_addr),
		.s_axi_9_w_ready(_mux_s_axi_9_w_ready),
		.s_axi_9_w_valid(_argRouteRvm_9_axi_w_valid),
		.s_axi_9_w_bits_data(_argRouteRvm_9_axi_w_bits_data),
		.s_axi_9_b_valid(_mux_s_axi_9_b_valid),
		.s_axi_10_ar_ready(_mux_s_axi_10_ar_ready),
		.s_axi_10_ar_valid(_argRouteRvm_10_axi_ar_valid),
		.s_axi_10_ar_bits_addr(_argRouteRvm_10_axi_ar_bits_addr),
		.s_axi_10_r_ready(_argRouteRvm_10_axi_r_ready),
		.s_axi_10_r_valid(_mux_s_axi_10_r_valid),
		.s_axi_10_r_bits_data(_mux_s_axi_10_r_bits_data),
		.s_axi_10_aw_ready(_mux_s_axi_10_aw_ready),
		.s_axi_10_aw_valid(_argRouteRvm_10_axi_aw_valid),
		.s_axi_10_aw_bits_addr(_argRouteRvm_10_axi_aw_bits_addr),
		.s_axi_10_w_ready(_mux_s_axi_10_w_ready),
		.s_axi_10_w_valid(_argRouteRvm_10_axi_w_valid),
		.s_axi_10_w_bits_data(_argRouteRvm_10_axi_w_bits_data),
		.s_axi_10_b_valid(_mux_s_axi_10_b_valid),
		.s_axi_11_ar_ready(_mux_s_axi_11_ar_ready),
		.s_axi_11_ar_valid(_argRouteRvm_11_axi_ar_valid),
		.s_axi_11_ar_bits_addr(_argRouteRvm_11_axi_ar_bits_addr),
		.s_axi_11_r_ready(_argRouteRvm_11_axi_r_ready),
		.s_axi_11_r_valid(_mux_s_axi_11_r_valid),
		.s_axi_11_r_bits_data(_mux_s_axi_11_r_bits_data),
		.s_axi_11_aw_ready(_mux_s_axi_11_aw_ready),
		.s_axi_11_aw_valid(_argRouteRvm_11_axi_aw_valid),
		.s_axi_11_aw_bits_addr(_argRouteRvm_11_axi_aw_bits_addr),
		.s_axi_11_w_ready(_mux_s_axi_11_w_ready),
		.s_axi_11_w_valid(_argRouteRvm_11_axi_w_valid),
		.s_axi_11_w_bits_data(_argRouteRvm_11_axi_w_bits_data),
		.s_axi_11_b_valid(_mux_s_axi_11_b_valid),
		.s_axi_12_ar_ready(_mux_s_axi_12_ar_ready),
		.s_axi_12_ar_valid(_argRouteRvm_12_axi_ar_valid),
		.s_axi_12_ar_bits_addr(_argRouteRvm_12_axi_ar_bits_addr),
		.s_axi_12_r_ready(_argRouteRvm_12_axi_r_ready),
		.s_axi_12_r_valid(_mux_s_axi_12_r_valid),
		.s_axi_12_r_bits_data(_mux_s_axi_12_r_bits_data),
		.s_axi_12_aw_ready(_mux_s_axi_12_aw_ready),
		.s_axi_12_aw_valid(_argRouteRvm_12_axi_aw_valid),
		.s_axi_12_aw_bits_addr(_argRouteRvm_12_axi_aw_bits_addr),
		.s_axi_12_w_ready(_mux_s_axi_12_w_ready),
		.s_axi_12_w_valid(_argRouteRvm_12_axi_w_valid),
		.s_axi_12_w_bits_data(_argRouteRvm_12_axi_w_bits_data),
		.s_axi_12_b_valid(_mux_s_axi_12_b_valid),
		.s_axi_13_ar_ready(_mux_s_axi_13_ar_ready),
		.s_axi_13_ar_valid(_argRouteRvm_13_axi_ar_valid),
		.s_axi_13_ar_bits_addr(_argRouteRvm_13_axi_ar_bits_addr),
		.s_axi_13_r_ready(_argRouteRvm_13_axi_r_ready),
		.s_axi_13_r_valid(_mux_s_axi_13_r_valid),
		.s_axi_13_r_bits_data(_mux_s_axi_13_r_bits_data),
		.s_axi_13_aw_ready(_mux_s_axi_13_aw_ready),
		.s_axi_13_aw_valid(_argRouteRvm_13_axi_aw_valid),
		.s_axi_13_aw_bits_addr(_argRouteRvm_13_axi_aw_bits_addr),
		.s_axi_13_w_ready(_mux_s_axi_13_w_ready),
		.s_axi_13_w_valid(_argRouteRvm_13_axi_w_valid),
		.s_axi_13_w_bits_data(_argRouteRvm_13_axi_w_bits_data),
		.s_axi_13_b_valid(_mux_s_axi_13_b_valid),
		.s_axi_14_ar_ready(_mux_s_axi_14_ar_ready),
		.s_axi_14_ar_valid(_argRouteRvm_14_axi_ar_valid),
		.s_axi_14_ar_bits_addr(_argRouteRvm_14_axi_ar_bits_addr),
		.s_axi_14_r_ready(_argRouteRvm_14_axi_r_ready),
		.s_axi_14_r_valid(_mux_s_axi_14_r_valid),
		.s_axi_14_r_bits_data(_mux_s_axi_14_r_bits_data),
		.s_axi_14_aw_ready(_mux_s_axi_14_aw_ready),
		.s_axi_14_aw_valid(_argRouteRvm_14_axi_aw_valid),
		.s_axi_14_aw_bits_addr(_argRouteRvm_14_axi_aw_bits_addr),
		.s_axi_14_w_ready(_mux_s_axi_14_w_ready),
		.s_axi_14_w_valid(_argRouteRvm_14_axi_w_valid),
		.s_axi_14_w_bits_data(_argRouteRvm_14_axi_w_bits_data),
		.s_axi_14_b_valid(_mux_s_axi_14_b_valid),
		.s_axi_15_ar_ready(_mux_s_axi_15_ar_ready),
		.s_axi_15_ar_valid(_argRouteRvm_15_axi_ar_valid),
		.s_axi_15_ar_bits_addr(_argRouteRvm_15_axi_ar_bits_addr),
		.s_axi_15_r_ready(_argRouteRvm_15_axi_r_ready),
		.s_axi_15_r_valid(_mux_s_axi_15_r_valid),
		.s_axi_15_r_bits_data(_mux_s_axi_15_r_bits_data),
		.s_axi_15_aw_ready(_mux_s_axi_15_aw_ready),
		.s_axi_15_aw_valid(_argRouteRvm_15_axi_aw_valid),
		.s_axi_15_aw_bits_addr(_argRouteRvm_15_axi_aw_bits_addr),
		.s_axi_15_w_ready(_mux_s_axi_15_w_ready),
		.s_axi_15_w_valid(_argRouteRvm_15_axi_w_valid),
		.s_axi_15_w_bits_data(_argRouteRvm_15_axi_w_bits_data),
		.s_axi_15_b_valid(_mux_s_axi_15_b_valid),
		.s_axi_16_ar_ready(_mux_s_axi_16_ar_ready),
		.s_axi_16_ar_valid(_argRouteRvmReadOnly_0_axi_ar_valid),
		.s_axi_16_ar_bits_addr(_argRouteRvmReadOnly_0_axi_ar_bits_addr),
		.s_axi_16_r_ready(_argRouteRvmReadOnly_0_axi_r_ready),
		.s_axi_16_r_valid(_mux_s_axi_16_r_valid),
		.s_axi_16_r_bits_data(_mux_s_axi_16_r_bits_data),
		.s_axi_17_ar_ready(_mux_s_axi_17_ar_ready),
		.s_axi_17_ar_valid(_argRouteRvmReadOnly_1_axi_ar_valid),
		.s_axi_17_ar_bits_addr(_argRouteRvmReadOnly_1_axi_ar_bits_addr),
		.s_axi_17_r_ready(_argRouteRvmReadOnly_1_axi_r_ready),
		.s_axi_17_r_valid(_mux_s_axi_17_r_valid),
		.s_axi_17_r_bits_data(_mux_s_axi_17_r_bits_data),
		.s_axi_18_ar_ready(_mux_s_axi_18_ar_ready),
		.s_axi_18_ar_valid(_argRouteRvmReadOnly_2_axi_ar_valid),
		.s_axi_18_ar_bits_addr(_argRouteRvmReadOnly_2_axi_ar_bits_addr),
		.s_axi_18_r_ready(_argRouteRvmReadOnly_2_axi_r_ready),
		.s_axi_18_r_valid(_mux_s_axi_18_r_valid),
		.s_axi_18_r_bits_data(_mux_s_axi_18_r_bits_data),
		.s_axi_19_ar_ready(_mux_s_axi_19_ar_ready),
		.s_axi_19_ar_valid(_argRouteRvmReadOnly_3_axi_ar_valid),
		.s_axi_19_ar_bits_addr(_argRouteRvmReadOnly_3_axi_ar_bits_addr),
		.s_axi_19_r_ready(_argRouteRvmReadOnly_3_axi_r_ready),
		.s_axi_19_r_valid(_mux_s_axi_19_r_valid),
		.s_axi_19_r_bits_data(_mux_s_axi_19_r_bits_data),
		.s_axi_20_ar_ready(_mux_s_axi_20_ar_ready),
		.s_axi_20_ar_valid(_argRouteRvmReadOnly_4_axi_ar_valid),
		.s_axi_20_ar_bits_addr(_argRouteRvmReadOnly_4_axi_ar_bits_addr),
		.s_axi_20_r_ready(_argRouteRvmReadOnly_4_axi_r_ready),
		.s_axi_20_r_valid(_mux_s_axi_20_r_valid),
		.s_axi_20_r_bits_data(_mux_s_axi_20_r_bits_data),
		.s_axi_21_ar_ready(_mux_s_axi_21_ar_ready),
		.s_axi_21_ar_valid(_argRouteRvmReadOnly_5_axi_ar_valid),
		.s_axi_21_ar_bits_addr(_argRouteRvmReadOnly_5_axi_ar_bits_addr),
		.s_axi_21_r_ready(_argRouteRvmReadOnly_5_axi_r_ready),
		.s_axi_21_r_valid(_mux_s_axi_21_r_valid),
		.s_axi_21_r_bits_data(_mux_s_axi_21_r_bits_data),
		.s_axi_22_ar_ready(_mux_s_axi_22_ar_ready),
		.s_axi_22_ar_valid(_argRouteRvmReadOnly_6_axi_ar_valid),
		.s_axi_22_ar_bits_addr(_argRouteRvmReadOnly_6_axi_ar_bits_addr),
		.s_axi_22_r_ready(_argRouteRvmReadOnly_6_axi_r_ready),
		.s_axi_22_r_valid(_mux_s_axi_22_r_valid),
		.s_axi_22_r_bits_data(_mux_s_axi_22_r_bits_data),
		.s_axi_23_ar_ready(_mux_s_axi_23_ar_ready),
		.s_axi_23_ar_valid(_argRouteRvmReadOnly_7_axi_ar_valid),
		.s_axi_23_ar_bits_addr(_argRouteRvmReadOnly_7_axi_ar_bits_addr),
		.s_axi_23_r_ready(_argRouteRvmReadOnly_7_axi_r_ready),
		.s_axi_23_r_valid(_mux_s_axi_23_r_valid),
		.s_axi_23_r_bits_data(_mux_s_axi_23_r_bits_data),
		.s_axi_24_ar_ready(_mux_s_axi_24_ar_ready),
		.s_axi_24_ar_valid(_argRouteRvmReadOnly_8_axi_ar_valid),
		.s_axi_24_ar_bits_addr(_argRouteRvmReadOnly_8_axi_ar_bits_addr),
		.s_axi_24_r_ready(_argRouteRvmReadOnly_8_axi_r_ready),
		.s_axi_24_r_valid(_mux_s_axi_24_r_valid),
		.s_axi_24_r_bits_data(_mux_s_axi_24_r_bits_data),
		.s_axi_25_ar_ready(_mux_s_axi_25_ar_ready),
		.s_axi_25_ar_valid(_argRouteRvmReadOnly_9_axi_ar_valid),
		.s_axi_25_ar_bits_addr(_argRouteRvmReadOnly_9_axi_ar_bits_addr),
		.s_axi_25_r_ready(_argRouteRvmReadOnly_9_axi_r_ready),
		.s_axi_25_r_valid(_mux_s_axi_25_r_valid),
		.s_axi_25_r_bits_data(_mux_s_axi_25_r_bits_data),
		.s_axi_26_ar_ready(_mux_s_axi_26_ar_ready),
		.s_axi_26_ar_valid(_argRouteRvmReadOnly_10_axi_ar_valid),
		.s_axi_26_ar_bits_addr(_argRouteRvmReadOnly_10_axi_ar_bits_addr),
		.s_axi_26_r_ready(_argRouteRvmReadOnly_10_axi_r_ready),
		.s_axi_26_r_valid(_mux_s_axi_26_r_valid),
		.s_axi_26_r_bits_data(_mux_s_axi_26_r_bits_data),
		.s_axi_27_ar_ready(_mux_s_axi_27_ar_ready),
		.s_axi_27_ar_valid(_argRouteRvmReadOnly_11_axi_ar_valid),
		.s_axi_27_ar_bits_addr(_argRouteRvmReadOnly_11_axi_ar_bits_addr),
		.s_axi_27_r_ready(_argRouteRvmReadOnly_11_axi_r_ready),
		.s_axi_27_r_valid(_mux_s_axi_27_r_valid),
		.s_axi_27_r_bits_data(_mux_s_axi_27_r_bits_data),
		.s_axi_28_ar_ready(_mux_s_axi_28_ar_ready),
		.s_axi_28_ar_valid(_argRouteRvmReadOnly_12_axi_ar_valid),
		.s_axi_28_ar_bits_addr(_argRouteRvmReadOnly_12_axi_ar_bits_addr),
		.s_axi_28_r_ready(_argRouteRvmReadOnly_12_axi_r_ready),
		.s_axi_28_r_valid(_mux_s_axi_28_r_valid),
		.s_axi_28_r_bits_data(_mux_s_axi_28_r_bits_data),
		.s_axi_29_ar_ready(_mux_s_axi_29_ar_ready),
		.s_axi_29_ar_valid(_argRouteRvmReadOnly_13_axi_ar_valid),
		.s_axi_29_ar_bits_addr(_argRouteRvmReadOnly_13_axi_ar_bits_addr),
		.s_axi_29_r_ready(_argRouteRvmReadOnly_13_axi_r_ready),
		.s_axi_29_r_valid(_mux_s_axi_29_r_valid),
		.s_axi_29_r_bits_data(_mux_s_axi_29_r_bits_data),
		.s_axi_30_ar_ready(_mux_s_axi_30_ar_ready),
		.s_axi_30_ar_valid(_argRouteRvmReadOnly_14_axi_ar_valid),
		.s_axi_30_ar_bits_addr(_argRouteRvmReadOnly_14_axi_ar_bits_addr),
		.s_axi_30_r_ready(_argRouteRvmReadOnly_14_axi_r_ready),
		.s_axi_30_r_valid(_mux_s_axi_30_r_valid),
		.s_axi_30_r_bits_data(_mux_s_axi_30_r_bits_data),
		.s_axi_31_ar_ready(_mux_s_axi_31_ar_ready),
		.s_axi_31_ar_valid(_argRouteRvmReadOnly_15_axi_ar_valid),
		.s_axi_31_ar_bits_addr(_argRouteRvmReadOnly_15_axi_ar_bits_addr),
		.s_axi_31_r_ready(_argRouteRvmReadOnly_15_axi_r_ready),
		.s_axi_31_r_valid(_mux_s_axi_31_r_valid),
		.s_axi_31_r_bits_data(_mux_s_axi_31_r_bits_data),
		.m_axi_ar_ready(axi_full_argRoute_0_ar_ready),
		.m_axi_ar_valid(axi_full_argRoute_0_ar_valid),
		.m_axi_ar_bits_id(axi_full_argRoute_0_ar_bits_id),
		.m_axi_ar_bits_addr(axi_full_argRoute_0_ar_bits_addr),
		.m_axi_ar_bits_len(axi_full_argRoute_0_ar_bits_len),
		.m_axi_ar_bits_size(axi_full_argRoute_0_ar_bits_size),
		.m_axi_ar_bits_burst(axi_full_argRoute_0_ar_bits_burst),
		.m_axi_ar_bits_lock(axi_full_argRoute_0_ar_bits_lock),
		.m_axi_ar_bits_cache(axi_full_argRoute_0_ar_bits_cache),
		.m_axi_ar_bits_prot(axi_full_argRoute_0_ar_bits_prot),
		.m_axi_ar_bits_qos(axi_full_argRoute_0_ar_bits_qos),
		.m_axi_ar_bits_region(axi_full_argRoute_0_ar_bits_region),
		.m_axi_r_ready(axi_full_argRoute_0_r_ready),
		.m_axi_r_valid(axi_full_argRoute_0_r_valid),
		.m_axi_r_bits_id(axi_full_argRoute_0_r_bits_id),
		.m_axi_r_bits_data(axi_full_argRoute_0_r_bits_data),
		.m_axi_r_bits_resp(axi_full_argRoute_0_r_bits_resp),
		.m_axi_r_bits_last(axi_full_argRoute_0_r_bits_last),
		.m_axi_aw_ready(axi_full_argRoute_0_aw_ready),
		.m_axi_aw_valid(axi_full_argRoute_0_aw_valid),
		.m_axi_aw_bits_id(axi_full_argRoute_0_aw_bits_id),
		.m_axi_aw_bits_addr(axi_full_argRoute_0_aw_bits_addr),
		.m_axi_aw_bits_len(axi_full_argRoute_0_aw_bits_len),
		.m_axi_aw_bits_size(axi_full_argRoute_0_aw_bits_size),
		.m_axi_aw_bits_burst(axi_full_argRoute_0_aw_bits_burst),
		.m_axi_aw_bits_lock(axi_full_argRoute_0_aw_bits_lock),
		.m_axi_aw_bits_cache(axi_full_argRoute_0_aw_bits_cache),
		.m_axi_aw_bits_prot(axi_full_argRoute_0_aw_bits_prot),
		.m_axi_aw_bits_qos(axi_full_argRoute_0_aw_bits_qos),
		.m_axi_aw_bits_region(axi_full_argRoute_0_aw_bits_region),
		.m_axi_w_ready(axi_full_argRoute_0_w_ready),
		.m_axi_w_valid(axi_full_argRoute_0_w_valid),
		.m_axi_w_bits_data(axi_full_argRoute_0_w_bits_data),
		.m_axi_w_bits_strb(axi_full_argRoute_0_w_bits_strb),
		.m_axi_w_bits_last(axi_full_argRoute_0_w_bits_last),
		.m_axi_b_ready(axi_full_argRoute_0_b_ready),
		.m_axi_b_valid(axi_full_argRoute_0_b_valid),
		.m_axi_b_bits_id(axi_full_argRoute_0_b_bits_id),
		.m_axi_b_bits_resp(axi_full_argRoute_0_b_bits_resp)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_0(
		.io_dataIn_TREADY(_axis_stream_converters_in_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_0_TVALID),
		.io_dataIn_TDATA(io_export_argIn_0_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_0_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_0_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_1(
		.io_dataIn_TREADY(_axis_stream_converters_in_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_1_TVALID),
		.io_dataIn_TDATA(io_export_argIn_1_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_1_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_1_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_2(
		.io_dataIn_TREADY(_axis_stream_converters_in_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_2_TVALID),
		.io_dataIn_TDATA(io_export_argIn_2_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_2_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_2_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_3(
		.io_dataIn_TREADY(_axis_stream_converters_in_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_3_TVALID),
		.io_dataIn_TDATA(io_export_argIn_3_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_3_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_3_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_4(
		.io_dataIn_TREADY(_axis_stream_converters_in_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_4_TVALID),
		.io_dataIn_TDATA(io_export_argIn_4_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_4_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_4_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_5(
		.io_dataIn_TREADY(_axis_stream_converters_in_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_5_TVALID),
		.io_dataIn_TDATA(io_export_argIn_5_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_5_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_5_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_6(
		.io_dataIn_TREADY(_axis_stream_converters_in_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_6_TVALID),
		.io_dataIn_TDATA(io_export_argIn_6_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_6_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_6_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_7(
		.io_dataIn_TREADY(_axis_stream_converters_in_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_7_TVALID),
		.io_dataIn_TDATA(io_export_argIn_7_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_7_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_7_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_8(
		.io_dataIn_TREADY(_axis_stream_converters_in_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_8_TVALID),
		.io_dataIn_TDATA(io_export_argIn_8_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_8_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_8_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_9(
		.io_dataIn_TREADY(_axis_stream_converters_in_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_9_TVALID),
		.io_dataIn_TDATA(io_export_argIn_9_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_9_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_9_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_10(
		.io_dataIn_TREADY(_axis_stream_converters_in_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_10_TVALID),
		.io_dataIn_TDATA(io_export_argIn_10_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_10_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_10_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_11(
		.io_dataIn_TREADY(_axis_stream_converters_in_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_11_TVALID),
		.io_dataIn_TDATA(io_export_argIn_11_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_11_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_11_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_12(
		.io_dataIn_TREADY(_axis_stream_converters_in_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_12_TVALID),
		.io_dataIn_TDATA(io_export_argIn_12_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_12_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_12_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_13(
		.io_dataIn_TREADY(_axis_stream_converters_in_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_13_TVALID),
		.io_dataIn_TDATA(io_export_argIn_13_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_13_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_13_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_14(
		.io_dataIn_TREADY(_axis_stream_converters_in_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_14_TVALID),
		.io_dataIn_TDATA(io_export_argIn_14_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_14_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_14_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_15(
		.io_dataIn_TREADY(_axis_stream_converters_in_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_15_TVALID),
		.io_dataIn_TDATA(io_export_argIn_15_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_15_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_15_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_16(
		.io_dataIn_TREADY(_axis_stream_converters_in_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_16_TVALID),
		.io_dataIn_TDATA(io_export_argIn_16_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_16_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_16_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_17(
		.io_dataIn_TREADY(_axis_stream_converters_in_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_17_TVALID),
		.io_dataIn_TDATA(io_export_argIn_17_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_17_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_17_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_18(
		.io_dataIn_TREADY(_axis_stream_converters_in_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_18_TVALID),
		.io_dataIn_TDATA(io_export_argIn_18_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_18_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_18_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_19(
		.io_dataIn_TREADY(_axis_stream_converters_in_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_19_TVALID),
		.io_dataIn_TDATA(io_export_argIn_19_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_19_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_19_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_20(
		.io_dataIn_TREADY(_axis_stream_converters_in_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_20_TVALID),
		.io_dataIn_TDATA(io_export_argIn_20_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_20_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_20_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_21(
		.io_dataIn_TREADY(_axis_stream_converters_in_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_21_TVALID),
		.io_dataIn_TDATA(io_export_argIn_21_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_21_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_21_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_22(
		.io_dataIn_TREADY(_axis_stream_converters_in_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_22_TVALID),
		.io_dataIn_TDATA(io_export_argIn_22_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_22_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_22_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_23(
		.io_dataIn_TREADY(_axis_stream_converters_in_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_23_TVALID),
		.io_dataIn_TDATA(io_export_argIn_23_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_23_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_23_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_24(
		.io_dataIn_TREADY(_axis_stream_converters_in_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_24_TVALID),
		.io_dataIn_TDATA(io_export_argIn_24_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_24_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_24_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_25(
		.io_dataIn_TREADY(_axis_stream_converters_in_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_25_TVALID),
		.io_dataIn_TDATA(io_export_argIn_25_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_25_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_25_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_26(
		.io_dataIn_TREADY(_axis_stream_converters_in_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_26_TVALID),
		.io_dataIn_TDATA(io_export_argIn_26_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_26_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_26_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_27(
		.io_dataIn_TREADY(_axis_stream_converters_in_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_27_TVALID),
		.io_dataIn_TDATA(io_export_argIn_27_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_27_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_27_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_28(
		.io_dataIn_TREADY(_axis_stream_converters_in_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_28_TVALID),
		.io_dataIn_TDATA(io_export_argIn_28_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_28_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_28_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_29(
		.io_dataIn_TREADY(_axis_stream_converters_in_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_29_TVALID),
		.io_dataIn_TDATA(io_export_argIn_29_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_29_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_29_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_30(
		.io_dataIn_TREADY(_axis_stream_converters_in_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_30_TVALID),
		.io_dataIn_TDATA(io_export_argIn_30_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_30_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_30_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_31(
		.io_dataIn_TREADY(_axis_stream_converters_in_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_31_TVALID),
		.io_dataIn_TDATA(io_export_argIn_31_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_31_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_31_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_32(
		.io_dataIn_TREADY(_axis_stream_converters_in_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_32_TVALID),
		.io_dataIn_TDATA(io_export_argIn_32_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_32_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_32_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_33(
		.io_dataIn_TREADY(_axis_stream_converters_in_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_33_TVALID),
		.io_dataIn_TDATA(io_export_argIn_33_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_33_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_33_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_34(
		.io_dataIn_TREADY(_axis_stream_converters_in_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_34_TVALID),
		.io_dataIn_TDATA(io_export_argIn_34_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_34_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_34_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_35(
		.io_dataIn_TREADY(_axis_stream_converters_in_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_35_TVALID),
		.io_dataIn_TDATA(io_export_argIn_35_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_35_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_35_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_36(
		.io_dataIn_TREADY(_axis_stream_converters_in_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_36_TVALID),
		.io_dataIn_TDATA(io_export_argIn_36_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_36_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_36_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_37(
		.io_dataIn_TREADY(_axis_stream_converters_in_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_37_TVALID),
		.io_dataIn_TDATA(io_export_argIn_37_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_37_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_37_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_38(
		.io_dataIn_TREADY(_axis_stream_converters_in_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_38_TVALID),
		.io_dataIn_TDATA(io_export_argIn_38_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_38_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_38_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_39(
		.io_dataIn_TREADY(_axis_stream_converters_in_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_39_TVALID),
		.io_dataIn_TDATA(io_export_argIn_39_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_39_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_39_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_40(
		.io_dataIn_TREADY(_axis_stream_converters_in_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_40_TVALID),
		.io_dataIn_TDATA(io_export_argIn_40_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_40_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_40_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_41(
		.io_dataIn_TREADY(_axis_stream_converters_in_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_41_TVALID),
		.io_dataIn_TDATA(io_export_argIn_41_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_41_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_41_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_42(
		.io_dataIn_TREADY(_axis_stream_converters_in_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_42_TVALID),
		.io_dataIn_TDATA(io_export_argIn_42_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_42_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_42_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_43(
		.io_dataIn_TREADY(_axis_stream_converters_in_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_43_TVALID),
		.io_dataIn_TDATA(io_export_argIn_43_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_43_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_43_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_44(
		.io_dataIn_TREADY(_axis_stream_converters_in_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_44_TVALID),
		.io_dataIn_TDATA(io_export_argIn_44_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_44_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_44_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_45(
		.io_dataIn_TREADY(_axis_stream_converters_in_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_45_TVALID),
		.io_dataIn_TDATA(io_export_argIn_45_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_45_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_45_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_46(
		.io_dataIn_TREADY(_axis_stream_converters_in_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_46_TVALID),
		.io_dataIn_TDATA(io_export_argIn_46_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_46_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_46_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_47(
		.io_dataIn_TREADY(_axis_stream_converters_in_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_47_TVALID),
		.io_dataIn_TDATA(io_export_argIn_47_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_47_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_47_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_48(
		.io_dataIn_TREADY(_axis_stream_converters_in_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_48_TVALID),
		.io_dataIn_TDATA(io_export_argIn_48_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_48_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_48_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_49(
		.io_dataIn_TREADY(_axis_stream_converters_in_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_49_TVALID),
		.io_dataIn_TDATA(io_export_argIn_49_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_49_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_49_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_50(
		.io_dataIn_TREADY(_axis_stream_converters_in_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_50_TVALID),
		.io_dataIn_TDATA(io_export_argIn_50_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_50_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_50_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_51(
		.io_dataIn_TREADY(_axis_stream_converters_in_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_51_TVALID),
		.io_dataIn_TDATA(io_export_argIn_51_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_51_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_51_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_52(
		.io_dataIn_TREADY(_axis_stream_converters_in_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_52_TVALID),
		.io_dataIn_TDATA(io_export_argIn_52_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_52_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_52_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_53(
		.io_dataIn_TREADY(_axis_stream_converters_in_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_53_TVALID),
		.io_dataIn_TDATA(io_export_argIn_53_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_53_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_53_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_54(
		.io_dataIn_TREADY(_axis_stream_converters_in_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_54_TVALID),
		.io_dataIn_TDATA(io_export_argIn_54_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_54_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_54_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_55(
		.io_dataIn_TREADY(_axis_stream_converters_in_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_55_TVALID),
		.io_dataIn_TDATA(io_export_argIn_55_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_55_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_55_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_56(
		.io_dataIn_TREADY(_axis_stream_converters_in_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_56_TVALID),
		.io_dataIn_TDATA(io_export_argIn_56_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_56_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_56_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_57(
		.io_dataIn_TREADY(_axis_stream_converters_in_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_57_TVALID),
		.io_dataIn_TDATA(io_export_argIn_57_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_57_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_57_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_58(
		.io_dataIn_TREADY(_axis_stream_converters_in_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_58_TVALID),
		.io_dataIn_TDATA(io_export_argIn_58_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_58_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_58_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_59(
		.io_dataIn_TREADY(_axis_stream_converters_in_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_59_TVALID),
		.io_dataIn_TDATA(io_export_argIn_59_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_59_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_59_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_60(
		.io_dataIn_TREADY(_axis_stream_converters_in_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_60_TVALID),
		.io_dataIn_TDATA(io_export_argIn_60_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_60_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_60_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_61(
		.io_dataIn_TREADY(_axis_stream_converters_in_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_61_TVALID),
		.io_dataIn_TDATA(io_export_argIn_61_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_61_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_61_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_62(
		.io_dataIn_TREADY(_axis_stream_converters_in_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_62_TVALID),
		.io_dataIn_TDATA(io_export_argIn_62_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_62_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_62_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_63(
		.io_dataIn_TREADY(_axis_stream_converters_in_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_63_TVALID),
		.io_dataIn_TDATA(io_export_argIn_63_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_63_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_63_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_64(
		.io_dataIn_TREADY(_axis_stream_converters_in_64_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_64_TVALID),
		.io_dataIn_TDATA(io_export_argIn_64_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_64_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_64_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_64_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_65(
		.io_dataIn_TREADY(_axis_stream_converters_in_65_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_65_TVALID),
		.io_dataIn_TDATA(io_export_argIn_65_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_65_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_65_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_65_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_66(
		.io_dataIn_TREADY(_axis_stream_converters_in_66_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_66_TVALID),
		.io_dataIn_TDATA(io_export_argIn_66_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_66_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_66_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_66_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_67(
		.io_dataIn_TREADY(_axis_stream_converters_in_67_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_67_TVALID),
		.io_dataIn_TDATA(io_export_argIn_67_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_67_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_67_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_67_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_68(
		.io_dataIn_TREADY(_axis_stream_converters_in_68_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_68_TVALID),
		.io_dataIn_TDATA(io_export_argIn_68_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_68_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_68_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_68_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_69(
		.io_dataIn_TREADY(_axis_stream_converters_in_69_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_69_TVALID),
		.io_dataIn_TDATA(io_export_argIn_69_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_69_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_69_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_69_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_70(
		.io_dataIn_TREADY(_axis_stream_converters_in_70_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_70_TVALID),
		.io_dataIn_TDATA(io_export_argIn_70_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_70_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_70_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_70_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_71(
		.io_dataIn_TREADY(_axis_stream_converters_in_71_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_71_TVALID),
		.io_dataIn_TDATA(io_export_argIn_71_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_71_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_71_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_71_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_72(
		.io_dataIn_TREADY(_axis_stream_converters_in_72_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_72_TVALID),
		.io_dataIn_TDATA(io_export_argIn_72_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_72_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_72_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_72_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_73(
		.io_dataIn_TREADY(_axis_stream_converters_in_73_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_73_TVALID),
		.io_dataIn_TDATA(io_export_argIn_73_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_73_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_73_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_73_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_74(
		.io_dataIn_TREADY(_axis_stream_converters_in_74_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_74_TVALID),
		.io_dataIn_TDATA(io_export_argIn_74_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_74_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_74_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_74_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_75(
		.io_dataIn_TREADY(_axis_stream_converters_in_75_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_75_TVALID),
		.io_dataIn_TDATA(io_export_argIn_75_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_75_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_75_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_75_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_76(
		.io_dataIn_TREADY(_axis_stream_converters_in_76_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_76_TVALID),
		.io_dataIn_TDATA(io_export_argIn_76_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_76_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_76_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_76_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_77(
		.io_dataIn_TREADY(_axis_stream_converters_in_77_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_77_TVALID),
		.io_dataIn_TDATA(io_export_argIn_77_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_77_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_77_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_77_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_78(
		.io_dataIn_TREADY(_axis_stream_converters_in_78_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_78_TVALID),
		.io_dataIn_TDATA(io_export_argIn_78_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_78_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_78_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_78_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_79(
		.io_dataIn_TREADY(_axis_stream_converters_in_79_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_79_TVALID),
		.io_dataIn_TDATA(io_export_argIn_79_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_79_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_79_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_79_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_80(
		.io_dataIn_TREADY(_axis_stream_converters_in_80_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_80_TVALID),
		.io_dataIn_TDATA(io_export_argIn_80_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_80_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_80_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_80_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_81(
		.io_dataIn_TREADY(_axis_stream_converters_in_81_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_81_TVALID),
		.io_dataIn_TDATA(io_export_argIn_81_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_81_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_81_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_81_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_82(
		.io_dataIn_TREADY(_axis_stream_converters_in_82_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_82_TVALID),
		.io_dataIn_TDATA(io_export_argIn_82_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_82_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_82_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_82_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_83(
		.io_dataIn_TREADY(_axis_stream_converters_in_83_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_83_TVALID),
		.io_dataIn_TDATA(io_export_argIn_83_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_83_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_83_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_83_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_84(
		.io_dataIn_TREADY(_axis_stream_converters_in_84_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_84_TVALID),
		.io_dataIn_TDATA(io_export_argIn_84_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_84_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_84_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_84_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_85(
		.io_dataIn_TREADY(_axis_stream_converters_in_85_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_85_TVALID),
		.io_dataIn_TDATA(io_export_argIn_85_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_85_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_85_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_85_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_86(
		.io_dataIn_TREADY(_axis_stream_converters_in_86_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_86_TVALID),
		.io_dataIn_TDATA(io_export_argIn_86_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_86_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_86_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_86_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_87(
		.io_dataIn_TREADY(_axis_stream_converters_in_87_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_87_TVALID),
		.io_dataIn_TDATA(io_export_argIn_87_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_87_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_87_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_87_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_88(
		.io_dataIn_TREADY(_axis_stream_converters_in_88_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_88_TVALID),
		.io_dataIn_TDATA(io_export_argIn_88_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_88_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_88_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_88_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_89(
		.io_dataIn_TREADY(_axis_stream_converters_in_89_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_89_TVALID),
		.io_dataIn_TDATA(io_export_argIn_89_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_89_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_89_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_89_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_90(
		.io_dataIn_TREADY(_axis_stream_converters_in_90_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_90_TVALID),
		.io_dataIn_TDATA(io_export_argIn_90_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_90_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_90_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_90_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_91(
		.io_dataIn_TREADY(_axis_stream_converters_in_91_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_91_TVALID),
		.io_dataIn_TDATA(io_export_argIn_91_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_91_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_91_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_91_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_92(
		.io_dataIn_TREADY(_axis_stream_converters_in_92_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_92_TVALID),
		.io_dataIn_TDATA(io_export_argIn_92_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_92_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_92_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_92_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_93(
		.io_dataIn_TREADY(_axis_stream_converters_in_93_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_93_TVALID),
		.io_dataIn_TDATA(io_export_argIn_93_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_93_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_93_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_93_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_94(
		.io_dataIn_TREADY(_axis_stream_converters_in_94_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_94_TVALID),
		.io_dataIn_TDATA(io_export_argIn_94_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_94_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_94_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_94_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_95(
		.io_dataIn_TREADY(_axis_stream_converters_in_95_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_95_TVALID),
		.io_dataIn_TDATA(io_export_argIn_95_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_95_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_95_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_95_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_96(
		.io_dataIn_TREADY(_axis_stream_converters_in_96_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_96_TVALID),
		.io_dataIn_TDATA(io_export_argIn_96_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_96_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_96_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_96_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_97(
		.io_dataIn_TREADY(_axis_stream_converters_in_97_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_97_TVALID),
		.io_dataIn_TDATA(io_export_argIn_97_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_97_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_97_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_97_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_98(
		.io_dataIn_TREADY(_axis_stream_converters_in_98_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_98_TVALID),
		.io_dataIn_TDATA(io_export_argIn_98_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_98_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_98_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_98_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_99(
		.io_dataIn_TREADY(_axis_stream_converters_in_99_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_99_TVALID),
		.io_dataIn_TDATA(io_export_argIn_99_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_99_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_99_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_99_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_100(
		.io_dataIn_TREADY(_axis_stream_converters_in_100_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_100_TVALID),
		.io_dataIn_TDATA(io_export_argIn_100_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_100_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_100_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_100_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_101(
		.io_dataIn_TREADY(_axis_stream_converters_in_101_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_101_TVALID),
		.io_dataIn_TDATA(io_export_argIn_101_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_101_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_101_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_101_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_102(
		.io_dataIn_TREADY(_axis_stream_converters_in_102_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_102_TVALID),
		.io_dataIn_TDATA(io_export_argIn_102_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_102_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_102_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_102_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_103(
		.io_dataIn_TREADY(_axis_stream_converters_in_103_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_103_TVALID),
		.io_dataIn_TDATA(io_export_argIn_103_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_103_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_103_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_103_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_104(
		.io_dataIn_TREADY(_axis_stream_converters_in_104_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_104_TVALID),
		.io_dataIn_TDATA(io_export_argIn_104_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_104_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_104_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_104_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_105(
		.io_dataIn_TREADY(_axis_stream_converters_in_105_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_105_TVALID),
		.io_dataIn_TDATA(io_export_argIn_105_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_105_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_105_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_105_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_106(
		.io_dataIn_TREADY(_axis_stream_converters_in_106_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_106_TVALID),
		.io_dataIn_TDATA(io_export_argIn_106_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_106_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_106_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_106_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_107(
		.io_dataIn_TREADY(_axis_stream_converters_in_107_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_107_TVALID),
		.io_dataIn_TDATA(io_export_argIn_107_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_107_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_107_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_107_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_108(
		.io_dataIn_TREADY(_axis_stream_converters_in_108_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_108_TVALID),
		.io_dataIn_TDATA(io_export_argIn_108_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_108_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_108_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_108_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_109(
		.io_dataIn_TREADY(_axis_stream_converters_in_109_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_109_TVALID),
		.io_dataIn_TDATA(io_export_argIn_109_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_109_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_109_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_109_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_110(
		.io_dataIn_TREADY(_axis_stream_converters_in_110_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_110_TVALID),
		.io_dataIn_TDATA(io_export_argIn_110_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_110_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_110_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_110_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_111(
		.io_dataIn_TREADY(_axis_stream_converters_in_111_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_111_TVALID),
		.io_dataIn_TDATA(io_export_argIn_111_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_111_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_111_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_111_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_112(
		.io_dataIn_TREADY(_axis_stream_converters_in_112_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_112_TVALID),
		.io_dataIn_TDATA(io_export_argIn_112_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_112_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_112_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_112_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_113(
		.io_dataIn_TREADY(_axis_stream_converters_in_113_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_113_TVALID),
		.io_dataIn_TDATA(io_export_argIn_113_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_113_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_113_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_113_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_114(
		.io_dataIn_TREADY(_axis_stream_converters_in_114_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_114_TVALID),
		.io_dataIn_TDATA(io_export_argIn_114_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_114_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_114_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_114_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_115(
		.io_dataIn_TREADY(_axis_stream_converters_in_115_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_115_TVALID),
		.io_dataIn_TDATA(io_export_argIn_115_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_115_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_115_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_115_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_116(
		.io_dataIn_TREADY(_axis_stream_converters_in_116_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_116_TVALID),
		.io_dataIn_TDATA(io_export_argIn_116_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_116_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_116_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_116_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_117(
		.io_dataIn_TREADY(_axis_stream_converters_in_117_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_117_TVALID),
		.io_dataIn_TDATA(io_export_argIn_117_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_117_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_117_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_117_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_118(
		.io_dataIn_TREADY(_axis_stream_converters_in_118_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_118_TVALID),
		.io_dataIn_TDATA(io_export_argIn_118_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_118_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_118_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_118_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_119(
		.io_dataIn_TREADY(_axis_stream_converters_in_119_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_119_TVALID),
		.io_dataIn_TDATA(io_export_argIn_119_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_119_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_119_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_119_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_120(
		.io_dataIn_TREADY(_axis_stream_converters_in_120_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_120_TVALID),
		.io_dataIn_TDATA(io_export_argIn_120_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_120_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_120_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_120_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_121(
		.io_dataIn_TREADY(_axis_stream_converters_in_121_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_121_TVALID),
		.io_dataIn_TDATA(io_export_argIn_121_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_121_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_121_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_121_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_122(
		.io_dataIn_TREADY(_axis_stream_converters_in_122_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_122_TVALID),
		.io_dataIn_TDATA(io_export_argIn_122_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_122_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_122_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_122_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_123(
		.io_dataIn_TREADY(_axis_stream_converters_in_123_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_123_TVALID),
		.io_dataIn_TDATA(io_export_argIn_123_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_123_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_123_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_123_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_124(
		.io_dataIn_TREADY(_axis_stream_converters_in_124_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_124_TVALID),
		.io_dataIn_TDATA(io_export_argIn_124_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_124_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_124_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_124_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_125(
		.io_dataIn_TREADY(_axis_stream_converters_in_125_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_125_TVALID),
		.io_dataIn_TDATA(io_export_argIn_125_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_125_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_125_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_125_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_126(
		.io_dataIn_TREADY(_axis_stream_converters_in_126_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_126_TVALID),
		.io_dataIn_TDATA(io_export_argIn_126_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_126_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_126_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_126_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_192 axis_stream_converters_in_127(
		.io_dataIn_TREADY(_axis_stream_converters_in_127_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_127_TVALID),
		.io_dataIn_TDATA(io_export_argIn_127_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_127_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_127_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_127_io_dataOut_TDATA)
	);
	Counter64 argInCounter(
		.clock(clock),
		.reset(reset),
		.io_signals_0(io_export_argIn_0_TVALID & _axis_stream_converters_in_0_io_dataIn_TREADY),
		.io_signals_1(io_export_argIn_1_TVALID & _axis_stream_converters_in_1_io_dataIn_TREADY),
		.io_signals_2(io_export_argIn_2_TVALID & _axis_stream_converters_in_2_io_dataIn_TREADY),
		.io_signals_3(io_export_argIn_3_TVALID & _axis_stream_converters_in_3_io_dataIn_TREADY),
		.io_signals_4(io_export_argIn_4_TVALID & _axis_stream_converters_in_4_io_dataIn_TREADY),
		.io_signals_5(io_export_argIn_5_TVALID & _axis_stream_converters_in_5_io_dataIn_TREADY),
		.io_signals_6(io_export_argIn_6_TVALID & _axis_stream_converters_in_6_io_dataIn_TREADY),
		.io_signals_7(io_export_argIn_7_TVALID & _axis_stream_converters_in_7_io_dataIn_TREADY),
		.io_signals_8(io_export_argIn_8_TVALID & _axis_stream_converters_in_8_io_dataIn_TREADY),
		.io_signals_9(io_export_argIn_9_TVALID & _axis_stream_converters_in_9_io_dataIn_TREADY),
		.io_signals_10(io_export_argIn_10_TVALID & _axis_stream_converters_in_10_io_dataIn_TREADY),
		.io_signals_11(io_export_argIn_11_TVALID & _axis_stream_converters_in_11_io_dataIn_TREADY),
		.io_signals_12(io_export_argIn_12_TVALID & _axis_stream_converters_in_12_io_dataIn_TREADY),
		.io_signals_13(io_export_argIn_13_TVALID & _axis_stream_converters_in_13_io_dataIn_TREADY),
		.io_signals_14(io_export_argIn_14_TVALID & _axis_stream_converters_in_14_io_dataIn_TREADY),
		.io_signals_15(io_export_argIn_15_TVALID & _axis_stream_converters_in_15_io_dataIn_TREADY),
		.io_signals_16(io_export_argIn_16_TVALID & _axis_stream_converters_in_16_io_dataIn_TREADY),
		.io_signals_17(io_export_argIn_17_TVALID & _axis_stream_converters_in_17_io_dataIn_TREADY),
		.io_signals_18(io_export_argIn_18_TVALID & _axis_stream_converters_in_18_io_dataIn_TREADY),
		.io_signals_19(io_export_argIn_19_TVALID & _axis_stream_converters_in_19_io_dataIn_TREADY),
		.io_signals_20(io_export_argIn_20_TVALID & _axis_stream_converters_in_20_io_dataIn_TREADY),
		.io_signals_21(io_export_argIn_21_TVALID & _axis_stream_converters_in_21_io_dataIn_TREADY),
		.io_signals_22(io_export_argIn_22_TVALID & _axis_stream_converters_in_22_io_dataIn_TREADY),
		.io_signals_23(io_export_argIn_23_TVALID & _axis_stream_converters_in_23_io_dataIn_TREADY),
		.io_signals_24(io_export_argIn_24_TVALID & _axis_stream_converters_in_24_io_dataIn_TREADY),
		.io_signals_25(io_export_argIn_25_TVALID & _axis_stream_converters_in_25_io_dataIn_TREADY),
		.io_signals_26(io_export_argIn_26_TVALID & _axis_stream_converters_in_26_io_dataIn_TREADY),
		.io_signals_27(io_export_argIn_27_TVALID & _axis_stream_converters_in_27_io_dataIn_TREADY),
		.io_signals_28(io_export_argIn_28_TVALID & _axis_stream_converters_in_28_io_dataIn_TREADY),
		.io_signals_29(io_export_argIn_29_TVALID & _axis_stream_converters_in_29_io_dataIn_TREADY),
		.io_signals_30(io_export_argIn_30_TVALID & _axis_stream_converters_in_30_io_dataIn_TREADY),
		.io_signals_31(io_export_argIn_31_TVALID & _axis_stream_converters_in_31_io_dataIn_TREADY),
		.io_signals_32(io_export_argIn_32_TVALID & _axis_stream_converters_in_32_io_dataIn_TREADY),
		.io_signals_33(io_export_argIn_33_TVALID & _axis_stream_converters_in_33_io_dataIn_TREADY),
		.io_signals_34(io_export_argIn_34_TVALID & _axis_stream_converters_in_34_io_dataIn_TREADY),
		.io_signals_35(io_export_argIn_35_TVALID & _axis_stream_converters_in_35_io_dataIn_TREADY),
		.io_signals_36(io_export_argIn_36_TVALID & _axis_stream_converters_in_36_io_dataIn_TREADY),
		.io_signals_37(io_export_argIn_37_TVALID & _axis_stream_converters_in_37_io_dataIn_TREADY),
		.io_signals_38(io_export_argIn_38_TVALID & _axis_stream_converters_in_38_io_dataIn_TREADY),
		.io_signals_39(io_export_argIn_39_TVALID & _axis_stream_converters_in_39_io_dataIn_TREADY),
		.io_signals_40(io_export_argIn_40_TVALID & _axis_stream_converters_in_40_io_dataIn_TREADY),
		.io_signals_41(io_export_argIn_41_TVALID & _axis_stream_converters_in_41_io_dataIn_TREADY),
		.io_signals_42(io_export_argIn_42_TVALID & _axis_stream_converters_in_42_io_dataIn_TREADY),
		.io_signals_43(io_export_argIn_43_TVALID & _axis_stream_converters_in_43_io_dataIn_TREADY),
		.io_signals_44(io_export_argIn_44_TVALID & _axis_stream_converters_in_44_io_dataIn_TREADY),
		.io_signals_45(io_export_argIn_45_TVALID & _axis_stream_converters_in_45_io_dataIn_TREADY),
		.io_signals_46(io_export_argIn_46_TVALID & _axis_stream_converters_in_46_io_dataIn_TREADY),
		.io_signals_47(io_export_argIn_47_TVALID & _axis_stream_converters_in_47_io_dataIn_TREADY),
		.io_signals_48(io_export_argIn_48_TVALID & _axis_stream_converters_in_48_io_dataIn_TREADY),
		.io_signals_49(io_export_argIn_49_TVALID & _axis_stream_converters_in_49_io_dataIn_TREADY),
		.io_signals_50(io_export_argIn_50_TVALID & _axis_stream_converters_in_50_io_dataIn_TREADY),
		.io_signals_51(io_export_argIn_51_TVALID & _axis_stream_converters_in_51_io_dataIn_TREADY),
		.io_signals_52(io_export_argIn_52_TVALID & _axis_stream_converters_in_52_io_dataIn_TREADY),
		.io_signals_53(io_export_argIn_53_TVALID & _axis_stream_converters_in_53_io_dataIn_TREADY),
		.io_signals_54(io_export_argIn_54_TVALID & _axis_stream_converters_in_54_io_dataIn_TREADY),
		.io_signals_55(io_export_argIn_55_TVALID & _axis_stream_converters_in_55_io_dataIn_TREADY),
		.io_signals_56(io_export_argIn_56_TVALID & _axis_stream_converters_in_56_io_dataIn_TREADY),
		.io_signals_57(io_export_argIn_57_TVALID & _axis_stream_converters_in_57_io_dataIn_TREADY),
		.io_signals_58(io_export_argIn_58_TVALID & _axis_stream_converters_in_58_io_dataIn_TREADY),
		.io_signals_59(io_export_argIn_59_TVALID & _axis_stream_converters_in_59_io_dataIn_TREADY),
		.io_signals_60(io_export_argIn_60_TVALID & _axis_stream_converters_in_60_io_dataIn_TREADY),
		.io_signals_61(io_export_argIn_61_TVALID & _axis_stream_converters_in_61_io_dataIn_TREADY),
		.io_signals_62(io_export_argIn_62_TVALID & _axis_stream_converters_in_62_io_dataIn_TREADY),
		.io_signals_63(io_export_argIn_63_TVALID & _axis_stream_converters_in_63_io_dataIn_TREADY),
		.io_signals_64(io_export_argIn_64_TVALID & _axis_stream_converters_in_64_io_dataIn_TREADY),
		.io_signals_65(io_export_argIn_65_TVALID & _axis_stream_converters_in_65_io_dataIn_TREADY),
		.io_signals_66(io_export_argIn_66_TVALID & _axis_stream_converters_in_66_io_dataIn_TREADY),
		.io_signals_67(io_export_argIn_67_TVALID & _axis_stream_converters_in_67_io_dataIn_TREADY),
		.io_signals_68(io_export_argIn_68_TVALID & _axis_stream_converters_in_68_io_dataIn_TREADY),
		.io_signals_69(io_export_argIn_69_TVALID & _axis_stream_converters_in_69_io_dataIn_TREADY),
		.io_signals_70(io_export_argIn_70_TVALID & _axis_stream_converters_in_70_io_dataIn_TREADY),
		.io_signals_71(io_export_argIn_71_TVALID & _axis_stream_converters_in_71_io_dataIn_TREADY),
		.io_signals_72(io_export_argIn_72_TVALID & _axis_stream_converters_in_72_io_dataIn_TREADY),
		.io_signals_73(io_export_argIn_73_TVALID & _axis_stream_converters_in_73_io_dataIn_TREADY),
		.io_signals_74(io_export_argIn_74_TVALID & _axis_stream_converters_in_74_io_dataIn_TREADY),
		.io_signals_75(io_export_argIn_75_TVALID & _axis_stream_converters_in_75_io_dataIn_TREADY),
		.io_signals_76(io_export_argIn_76_TVALID & _axis_stream_converters_in_76_io_dataIn_TREADY),
		.io_signals_77(io_export_argIn_77_TVALID & _axis_stream_converters_in_77_io_dataIn_TREADY),
		.io_signals_78(io_export_argIn_78_TVALID & _axis_stream_converters_in_78_io_dataIn_TREADY),
		.io_signals_79(io_export_argIn_79_TVALID & _axis_stream_converters_in_79_io_dataIn_TREADY),
		.io_signals_80(io_export_argIn_80_TVALID & _axis_stream_converters_in_80_io_dataIn_TREADY),
		.io_signals_81(io_export_argIn_81_TVALID & _axis_stream_converters_in_81_io_dataIn_TREADY),
		.io_signals_82(io_export_argIn_82_TVALID & _axis_stream_converters_in_82_io_dataIn_TREADY),
		.io_signals_83(io_export_argIn_83_TVALID & _axis_stream_converters_in_83_io_dataIn_TREADY),
		.io_signals_84(io_export_argIn_84_TVALID & _axis_stream_converters_in_84_io_dataIn_TREADY),
		.io_signals_85(io_export_argIn_85_TVALID & _axis_stream_converters_in_85_io_dataIn_TREADY),
		.io_signals_86(io_export_argIn_86_TVALID & _axis_stream_converters_in_86_io_dataIn_TREADY),
		.io_signals_87(io_export_argIn_87_TVALID & _axis_stream_converters_in_87_io_dataIn_TREADY),
		.io_signals_88(io_export_argIn_88_TVALID & _axis_stream_converters_in_88_io_dataIn_TREADY),
		.io_signals_89(io_export_argIn_89_TVALID & _axis_stream_converters_in_89_io_dataIn_TREADY),
		.io_signals_90(io_export_argIn_90_TVALID & _axis_stream_converters_in_90_io_dataIn_TREADY),
		.io_signals_91(io_export_argIn_91_TVALID & _axis_stream_converters_in_91_io_dataIn_TREADY),
		.io_signals_92(io_export_argIn_92_TVALID & _axis_stream_converters_in_92_io_dataIn_TREADY),
		.io_signals_93(io_export_argIn_93_TVALID & _axis_stream_converters_in_93_io_dataIn_TREADY),
		.io_signals_94(io_export_argIn_94_TVALID & _axis_stream_converters_in_94_io_dataIn_TREADY),
		.io_signals_95(io_export_argIn_95_TVALID & _axis_stream_converters_in_95_io_dataIn_TREADY),
		.io_signals_96(io_export_argIn_96_TVALID & _axis_stream_converters_in_96_io_dataIn_TREADY),
		.io_signals_97(io_export_argIn_97_TVALID & _axis_stream_converters_in_97_io_dataIn_TREADY),
		.io_signals_98(io_export_argIn_98_TVALID & _axis_stream_converters_in_98_io_dataIn_TREADY),
		.io_signals_99(io_export_argIn_99_TVALID & _axis_stream_converters_in_99_io_dataIn_TREADY),
		.io_signals_100(io_export_argIn_100_TVALID & _axis_stream_converters_in_100_io_dataIn_TREADY),
		.io_signals_101(io_export_argIn_101_TVALID & _axis_stream_converters_in_101_io_dataIn_TREADY),
		.io_signals_102(io_export_argIn_102_TVALID & _axis_stream_converters_in_102_io_dataIn_TREADY),
		.io_signals_103(io_export_argIn_103_TVALID & _axis_stream_converters_in_103_io_dataIn_TREADY),
		.io_signals_104(io_export_argIn_104_TVALID & _axis_stream_converters_in_104_io_dataIn_TREADY),
		.io_signals_105(io_export_argIn_105_TVALID & _axis_stream_converters_in_105_io_dataIn_TREADY),
		.io_signals_106(io_export_argIn_106_TVALID & _axis_stream_converters_in_106_io_dataIn_TREADY),
		.io_signals_107(io_export_argIn_107_TVALID & _axis_stream_converters_in_107_io_dataIn_TREADY),
		.io_signals_108(io_export_argIn_108_TVALID & _axis_stream_converters_in_108_io_dataIn_TREADY),
		.io_signals_109(io_export_argIn_109_TVALID & _axis_stream_converters_in_109_io_dataIn_TREADY),
		.io_signals_110(io_export_argIn_110_TVALID & _axis_stream_converters_in_110_io_dataIn_TREADY),
		.io_signals_111(io_export_argIn_111_TVALID & _axis_stream_converters_in_111_io_dataIn_TREADY),
		.io_signals_112(io_export_argIn_112_TVALID & _axis_stream_converters_in_112_io_dataIn_TREADY),
		.io_signals_113(io_export_argIn_113_TVALID & _axis_stream_converters_in_113_io_dataIn_TREADY),
		.io_signals_114(io_export_argIn_114_TVALID & _axis_stream_converters_in_114_io_dataIn_TREADY),
		.io_signals_115(io_export_argIn_115_TVALID & _axis_stream_converters_in_115_io_dataIn_TREADY),
		.io_signals_116(io_export_argIn_116_TVALID & _axis_stream_converters_in_116_io_dataIn_TREADY),
		.io_signals_117(io_export_argIn_117_TVALID & _axis_stream_converters_in_117_io_dataIn_TREADY),
		.io_signals_118(io_export_argIn_118_TVALID & _axis_stream_converters_in_118_io_dataIn_TREADY),
		.io_signals_119(io_export_argIn_119_TVALID & _axis_stream_converters_in_119_io_dataIn_TREADY),
		.io_signals_120(io_export_argIn_120_TVALID & _axis_stream_converters_in_120_io_dataIn_TREADY),
		.io_signals_121(io_export_argIn_121_TVALID & _axis_stream_converters_in_121_io_dataIn_TREADY),
		.io_signals_122(io_export_argIn_122_TVALID & _axis_stream_converters_in_122_io_dataIn_TREADY),
		.io_signals_123(io_export_argIn_123_TVALID & _axis_stream_converters_in_123_io_dataIn_TREADY),
		.io_signals_124(io_export_argIn_124_TVALID & _axis_stream_converters_in_124_io_dataIn_TREADY),
		.io_signals_125(io_export_argIn_125_TVALID & _axis_stream_converters_in_125_io_dataIn_TREADY),
		.io_signals_126(io_export_argIn_126_TVALID & _axis_stream_converters_in_126_io_dataIn_TREADY),
		.io_signals_127(io_export_argIn_127_TVALID & _axis_stream_converters_in_127_io_dataIn_TREADY),
		.io_counter()
	);
	assign io_export_argIn_0_TREADY = _axis_stream_converters_in_0_io_dataIn_TREADY;
	assign io_export_argIn_1_TREADY = _axis_stream_converters_in_1_io_dataIn_TREADY;
	assign io_export_argIn_2_TREADY = _axis_stream_converters_in_2_io_dataIn_TREADY;
	assign io_export_argIn_3_TREADY = _axis_stream_converters_in_3_io_dataIn_TREADY;
	assign io_export_argIn_4_TREADY = _axis_stream_converters_in_4_io_dataIn_TREADY;
	assign io_export_argIn_5_TREADY = _axis_stream_converters_in_5_io_dataIn_TREADY;
	assign io_export_argIn_6_TREADY = _axis_stream_converters_in_6_io_dataIn_TREADY;
	assign io_export_argIn_7_TREADY = _axis_stream_converters_in_7_io_dataIn_TREADY;
	assign io_export_argIn_8_TREADY = _axis_stream_converters_in_8_io_dataIn_TREADY;
	assign io_export_argIn_9_TREADY = _axis_stream_converters_in_9_io_dataIn_TREADY;
	assign io_export_argIn_10_TREADY = _axis_stream_converters_in_10_io_dataIn_TREADY;
	assign io_export_argIn_11_TREADY = _axis_stream_converters_in_11_io_dataIn_TREADY;
	assign io_export_argIn_12_TREADY = _axis_stream_converters_in_12_io_dataIn_TREADY;
	assign io_export_argIn_13_TREADY = _axis_stream_converters_in_13_io_dataIn_TREADY;
	assign io_export_argIn_14_TREADY = _axis_stream_converters_in_14_io_dataIn_TREADY;
	assign io_export_argIn_15_TREADY = _axis_stream_converters_in_15_io_dataIn_TREADY;
	assign io_export_argIn_16_TREADY = _axis_stream_converters_in_16_io_dataIn_TREADY;
	assign io_export_argIn_17_TREADY = _axis_stream_converters_in_17_io_dataIn_TREADY;
	assign io_export_argIn_18_TREADY = _axis_stream_converters_in_18_io_dataIn_TREADY;
	assign io_export_argIn_19_TREADY = _axis_stream_converters_in_19_io_dataIn_TREADY;
	assign io_export_argIn_20_TREADY = _axis_stream_converters_in_20_io_dataIn_TREADY;
	assign io_export_argIn_21_TREADY = _axis_stream_converters_in_21_io_dataIn_TREADY;
	assign io_export_argIn_22_TREADY = _axis_stream_converters_in_22_io_dataIn_TREADY;
	assign io_export_argIn_23_TREADY = _axis_stream_converters_in_23_io_dataIn_TREADY;
	assign io_export_argIn_24_TREADY = _axis_stream_converters_in_24_io_dataIn_TREADY;
	assign io_export_argIn_25_TREADY = _axis_stream_converters_in_25_io_dataIn_TREADY;
	assign io_export_argIn_26_TREADY = _axis_stream_converters_in_26_io_dataIn_TREADY;
	assign io_export_argIn_27_TREADY = _axis_stream_converters_in_27_io_dataIn_TREADY;
	assign io_export_argIn_28_TREADY = _axis_stream_converters_in_28_io_dataIn_TREADY;
	assign io_export_argIn_29_TREADY = _axis_stream_converters_in_29_io_dataIn_TREADY;
	assign io_export_argIn_30_TREADY = _axis_stream_converters_in_30_io_dataIn_TREADY;
	assign io_export_argIn_31_TREADY = _axis_stream_converters_in_31_io_dataIn_TREADY;
	assign io_export_argIn_32_TREADY = _axis_stream_converters_in_32_io_dataIn_TREADY;
	assign io_export_argIn_33_TREADY = _axis_stream_converters_in_33_io_dataIn_TREADY;
	assign io_export_argIn_34_TREADY = _axis_stream_converters_in_34_io_dataIn_TREADY;
	assign io_export_argIn_35_TREADY = _axis_stream_converters_in_35_io_dataIn_TREADY;
	assign io_export_argIn_36_TREADY = _axis_stream_converters_in_36_io_dataIn_TREADY;
	assign io_export_argIn_37_TREADY = _axis_stream_converters_in_37_io_dataIn_TREADY;
	assign io_export_argIn_38_TREADY = _axis_stream_converters_in_38_io_dataIn_TREADY;
	assign io_export_argIn_39_TREADY = _axis_stream_converters_in_39_io_dataIn_TREADY;
	assign io_export_argIn_40_TREADY = _axis_stream_converters_in_40_io_dataIn_TREADY;
	assign io_export_argIn_41_TREADY = _axis_stream_converters_in_41_io_dataIn_TREADY;
	assign io_export_argIn_42_TREADY = _axis_stream_converters_in_42_io_dataIn_TREADY;
	assign io_export_argIn_43_TREADY = _axis_stream_converters_in_43_io_dataIn_TREADY;
	assign io_export_argIn_44_TREADY = _axis_stream_converters_in_44_io_dataIn_TREADY;
	assign io_export_argIn_45_TREADY = _axis_stream_converters_in_45_io_dataIn_TREADY;
	assign io_export_argIn_46_TREADY = _axis_stream_converters_in_46_io_dataIn_TREADY;
	assign io_export_argIn_47_TREADY = _axis_stream_converters_in_47_io_dataIn_TREADY;
	assign io_export_argIn_48_TREADY = _axis_stream_converters_in_48_io_dataIn_TREADY;
	assign io_export_argIn_49_TREADY = _axis_stream_converters_in_49_io_dataIn_TREADY;
	assign io_export_argIn_50_TREADY = _axis_stream_converters_in_50_io_dataIn_TREADY;
	assign io_export_argIn_51_TREADY = _axis_stream_converters_in_51_io_dataIn_TREADY;
	assign io_export_argIn_52_TREADY = _axis_stream_converters_in_52_io_dataIn_TREADY;
	assign io_export_argIn_53_TREADY = _axis_stream_converters_in_53_io_dataIn_TREADY;
	assign io_export_argIn_54_TREADY = _axis_stream_converters_in_54_io_dataIn_TREADY;
	assign io_export_argIn_55_TREADY = _axis_stream_converters_in_55_io_dataIn_TREADY;
	assign io_export_argIn_56_TREADY = _axis_stream_converters_in_56_io_dataIn_TREADY;
	assign io_export_argIn_57_TREADY = _axis_stream_converters_in_57_io_dataIn_TREADY;
	assign io_export_argIn_58_TREADY = _axis_stream_converters_in_58_io_dataIn_TREADY;
	assign io_export_argIn_59_TREADY = _axis_stream_converters_in_59_io_dataIn_TREADY;
	assign io_export_argIn_60_TREADY = _axis_stream_converters_in_60_io_dataIn_TREADY;
	assign io_export_argIn_61_TREADY = _axis_stream_converters_in_61_io_dataIn_TREADY;
	assign io_export_argIn_62_TREADY = _axis_stream_converters_in_62_io_dataIn_TREADY;
	assign io_export_argIn_63_TREADY = _axis_stream_converters_in_63_io_dataIn_TREADY;
	assign io_export_argIn_64_TREADY = _axis_stream_converters_in_64_io_dataIn_TREADY;
	assign io_export_argIn_65_TREADY = _axis_stream_converters_in_65_io_dataIn_TREADY;
	assign io_export_argIn_66_TREADY = _axis_stream_converters_in_66_io_dataIn_TREADY;
	assign io_export_argIn_67_TREADY = _axis_stream_converters_in_67_io_dataIn_TREADY;
	assign io_export_argIn_68_TREADY = _axis_stream_converters_in_68_io_dataIn_TREADY;
	assign io_export_argIn_69_TREADY = _axis_stream_converters_in_69_io_dataIn_TREADY;
	assign io_export_argIn_70_TREADY = _axis_stream_converters_in_70_io_dataIn_TREADY;
	assign io_export_argIn_71_TREADY = _axis_stream_converters_in_71_io_dataIn_TREADY;
	assign io_export_argIn_72_TREADY = _axis_stream_converters_in_72_io_dataIn_TREADY;
	assign io_export_argIn_73_TREADY = _axis_stream_converters_in_73_io_dataIn_TREADY;
	assign io_export_argIn_74_TREADY = _axis_stream_converters_in_74_io_dataIn_TREADY;
	assign io_export_argIn_75_TREADY = _axis_stream_converters_in_75_io_dataIn_TREADY;
	assign io_export_argIn_76_TREADY = _axis_stream_converters_in_76_io_dataIn_TREADY;
	assign io_export_argIn_77_TREADY = _axis_stream_converters_in_77_io_dataIn_TREADY;
	assign io_export_argIn_78_TREADY = _axis_stream_converters_in_78_io_dataIn_TREADY;
	assign io_export_argIn_79_TREADY = _axis_stream_converters_in_79_io_dataIn_TREADY;
	assign io_export_argIn_80_TREADY = _axis_stream_converters_in_80_io_dataIn_TREADY;
	assign io_export_argIn_81_TREADY = _axis_stream_converters_in_81_io_dataIn_TREADY;
	assign io_export_argIn_82_TREADY = _axis_stream_converters_in_82_io_dataIn_TREADY;
	assign io_export_argIn_83_TREADY = _axis_stream_converters_in_83_io_dataIn_TREADY;
	assign io_export_argIn_84_TREADY = _axis_stream_converters_in_84_io_dataIn_TREADY;
	assign io_export_argIn_85_TREADY = _axis_stream_converters_in_85_io_dataIn_TREADY;
	assign io_export_argIn_86_TREADY = _axis_stream_converters_in_86_io_dataIn_TREADY;
	assign io_export_argIn_87_TREADY = _axis_stream_converters_in_87_io_dataIn_TREADY;
	assign io_export_argIn_88_TREADY = _axis_stream_converters_in_88_io_dataIn_TREADY;
	assign io_export_argIn_89_TREADY = _axis_stream_converters_in_89_io_dataIn_TREADY;
	assign io_export_argIn_90_TREADY = _axis_stream_converters_in_90_io_dataIn_TREADY;
	assign io_export_argIn_91_TREADY = _axis_stream_converters_in_91_io_dataIn_TREADY;
	assign io_export_argIn_92_TREADY = _axis_stream_converters_in_92_io_dataIn_TREADY;
	assign io_export_argIn_93_TREADY = _axis_stream_converters_in_93_io_dataIn_TREADY;
	assign io_export_argIn_94_TREADY = _axis_stream_converters_in_94_io_dataIn_TREADY;
	assign io_export_argIn_95_TREADY = _axis_stream_converters_in_95_io_dataIn_TREADY;
	assign io_export_argIn_96_TREADY = _axis_stream_converters_in_96_io_dataIn_TREADY;
	assign io_export_argIn_97_TREADY = _axis_stream_converters_in_97_io_dataIn_TREADY;
	assign io_export_argIn_98_TREADY = _axis_stream_converters_in_98_io_dataIn_TREADY;
	assign io_export_argIn_99_TREADY = _axis_stream_converters_in_99_io_dataIn_TREADY;
	assign io_export_argIn_100_TREADY = _axis_stream_converters_in_100_io_dataIn_TREADY;
	assign io_export_argIn_101_TREADY = _axis_stream_converters_in_101_io_dataIn_TREADY;
	assign io_export_argIn_102_TREADY = _axis_stream_converters_in_102_io_dataIn_TREADY;
	assign io_export_argIn_103_TREADY = _axis_stream_converters_in_103_io_dataIn_TREADY;
	assign io_export_argIn_104_TREADY = _axis_stream_converters_in_104_io_dataIn_TREADY;
	assign io_export_argIn_105_TREADY = _axis_stream_converters_in_105_io_dataIn_TREADY;
	assign io_export_argIn_106_TREADY = _axis_stream_converters_in_106_io_dataIn_TREADY;
	assign io_export_argIn_107_TREADY = _axis_stream_converters_in_107_io_dataIn_TREADY;
	assign io_export_argIn_108_TREADY = _axis_stream_converters_in_108_io_dataIn_TREADY;
	assign io_export_argIn_109_TREADY = _axis_stream_converters_in_109_io_dataIn_TREADY;
	assign io_export_argIn_110_TREADY = _axis_stream_converters_in_110_io_dataIn_TREADY;
	assign io_export_argIn_111_TREADY = _axis_stream_converters_in_111_io_dataIn_TREADY;
	assign io_export_argIn_112_TREADY = _axis_stream_converters_in_112_io_dataIn_TREADY;
	assign io_export_argIn_113_TREADY = _axis_stream_converters_in_113_io_dataIn_TREADY;
	assign io_export_argIn_114_TREADY = _axis_stream_converters_in_114_io_dataIn_TREADY;
	assign io_export_argIn_115_TREADY = _axis_stream_converters_in_115_io_dataIn_TREADY;
	assign io_export_argIn_116_TREADY = _axis_stream_converters_in_116_io_dataIn_TREADY;
	assign io_export_argIn_117_TREADY = _axis_stream_converters_in_117_io_dataIn_TREADY;
	assign io_export_argIn_118_TREADY = _axis_stream_converters_in_118_io_dataIn_TREADY;
	assign io_export_argIn_119_TREADY = _axis_stream_converters_in_119_io_dataIn_TREADY;
	assign io_export_argIn_120_TREADY = _axis_stream_converters_in_120_io_dataIn_TREADY;
	assign io_export_argIn_121_TREADY = _axis_stream_converters_in_121_io_dataIn_TREADY;
	assign io_export_argIn_122_TREADY = _axis_stream_converters_in_122_io_dataIn_TREADY;
	assign io_export_argIn_123_TREADY = _axis_stream_converters_in_123_io_dataIn_TREADY;
	assign io_export_argIn_124_TREADY = _axis_stream_converters_in_124_io_dataIn_TREADY;
	assign io_export_argIn_125_TREADY = _axis_stream_converters_in_125_io_dataIn_TREADY;
	assign io_export_argIn_126_TREADY = _axis_stream_converters_in_126_io_dataIn_TREADY;
	assign io_export_argIn_127_TREADY = _axis_stream_converters_in_127_io_dataIn_TREADY;
endmodule
module fibonacci (
	clock,
	reset,
	s_axil_mgmt_hardcilk_ARREADY,
	s_axil_mgmt_hardcilk_ARVALID,
	s_axil_mgmt_hardcilk_ARADDR,
	s_axil_mgmt_hardcilk_ARPROT,
	s_axil_mgmt_hardcilk_RREADY,
	s_axil_mgmt_hardcilk_RVALID,
	s_axil_mgmt_hardcilk_RDATA,
	s_axil_mgmt_hardcilk_RRESP,
	s_axil_mgmt_hardcilk_AWREADY,
	s_axil_mgmt_hardcilk_AWVALID,
	s_axil_mgmt_hardcilk_AWADDR,
	s_axil_mgmt_hardcilk_AWPROT,
	s_axil_mgmt_hardcilk_WREADY,
	s_axil_mgmt_hardcilk_WVALID,
	s_axil_mgmt_hardcilk_WDATA,
	s_axil_mgmt_hardcilk_WSTRB,
	s_axil_mgmt_hardcilk_BREADY,
	s_axil_mgmt_hardcilk_BVALID,
	s_axil_mgmt_hardcilk_BRESP,
	fib_0_m_axi_gmem_ARREADY,
	fib_0_m_axi_gmem_ARVALID,
	fib_0_m_axi_gmem_ARID,
	fib_0_m_axi_gmem_ARADDR,
	fib_0_m_axi_gmem_ARLEN,
	fib_0_m_axi_gmem_ARSIZE,
	fib_0_m_axi_gmem_ARBURST,
	fib_0_m_axi_gmem_ARLOCK,
	fib_0_m_axi_gmem_ARCACHE,
	fib_0_m_axi_gmem_ARPROT,
	fib_0_m_axi_gmem_ARQOS,
	fib_0_m_axi_gmem_ARREGION,
	fib_0_m_axi_gmem_ARUSER,
	fib_0_m_axi_gmem_RREADY,
	fib_0_m_axi_gmem_RVALID,
	fib_0_m_axi_gmem_RID,
	fib_0_m_axi_gmem_RDATA,
	fib_0_m_axi_gmem_RRESP,
	fib_0_m_axi_gmem_RLAST,
	fib_0_m_axi_gmem_RUSER,
	fib_0_m_axi_gmem_AWREADY,
	fib_0_m_axi_gmem_AWVALID,
	fib_0_m_axi_gmem_AWID,
	fib_0_m_axi_gmem_AWADDR,
	fib_0_m_axi_gmem_AWLEN,
	fib_0_m_axi_gmem_AWSIZE,
	fib_0_m_axi_gmem_AWBURST,
	fib_0_m_axi_gmem_AWLOCK,
	fib_0_m_axi_gmem_AWCACHE,
	fib_0_m_axi_gmem_AWPROT,
	fib_0_m_axi_gmem_AWQOS,
	fib_0_m_axi_gmem_AWREGION,
	fib_0_m_axi_gmem_AWUSER,
	fib_0_m_axi_gmem_WREADY,
	fib_0_m_axi_gmem_WVALID,
	fib_0_m_axi_gmem_WDATA,
	fib_0_m_axi_gmem_WSTRB,
	fib_0_m_axi_gmem_WLAST,
	fib_0_m_axi_gmem_WUSER,
	fib_0_m_axi_gmem_BREADY,
	fib_0_m_axi_gmem_BVALID,
	fib_0_m_axi_gmem_BID,
	fib_0_m_axi_gmem_BRESP,
	fib_0_m_axi_gmem_BUSER,
	fib_0_s_axi_control_ARREADY,
	fib_0_s_axi_control_ARVALID,
	fib_0_s_axi_control_ARADDR,
	fib_0_s_axi_control_RREADY,
	fib_0_s_axi_control_RVALID,
	fib_0_s_axi_control_RDATA,
	fib_0_s_axi_control_RRESP,
	fib_0_s_axi_control_AWREADY,
	fib_0_s_axi_control_AWVALID,
	fib_0_s_axi_control_AWADDR,
	fib_0_s_axi_control_WREADY,
	fib_0_s_axi_control_WVALID,
	fib_0_s_axi_control_WDATA,
	fib_0_s_axi_control_WSTRB,
	fib_0_s_axi_control_BREADY,
	fib_0_s_axi_control_BVALID,
	fib_0_s_axi_control_BRESP,
	fib_1_m_axi_gmem_ARREADY,
	fib_1_m_axi_gmem_ARVALID,
	fib_1_m_axi_gmem_ARID,
	fib_1_m_axi_gmem_ARADDR,
	fib_1_m_axi_gmem_ARLEN,
	fib_1_m_axi_gmem_ARSIZE,
	fib_1_m_axi_gmem_ARBURST,
	fib_1_m_axi_gmem_ARLOCK,
	fib_1_m_axi_gmem_ARCACHE,
	fib_1_m_axi_gmem_ARPROT,
	fib_1_m_axi_gmem_ARQOS,
	fib_1_m_axi_gmem_ARREGION,
	fib_1_m_axi_gmem_ARUSER,
	fib_1_m_axi_gmem_RREADY,
	fib_1_m_axi_gmem_RVALID,
	fib_1_m_axi_gmem_RID,
	fib_1_m_axi_gmem_RDATA,
	fib_1_m_axi_gmem_RRESP,
	fib_1_m_axi_gmem_RLAST,
	fib_1_m_axi_gmem_RUSER,
	fib_1_m_axi_gmem_AWREADY,
	fib_1_m_axi_gmem_AWVALID,
	fib_1_m_axi_gmem_AWID,
	fib_1_m_axi_gmem_AWADDR,
	fib_1_m_axi_gmem_AWLEN,
	fib_1_m_axi_gmem_AWSIZE,
	fib_1_m_axi_gmem_AWBURST,
	fib_1_m_axi_gmem_AWLOCK,
	fib_1_m_axi_gmem_AWCACHE,
	fib_1_m_axi_gmem_AWPROT,
	fib_1_m_axi_gmem_AWQOS,
	fib_1_m_axi_gmem_AWREGION,
	fib_1_m_axi_gmem_AWUSER,
	fib_1_m_axi_gmem_WREADY,
	fib_1_m_axi_gmem_WVALID,
	fib_1_m_axi_gmem_WDATA,
	fib_1_m_axi_gmem_WSTRB,
	fib_1_m_axi_gmem_WLAST,
	fib_1_m_axi_gmem_WUSER,
	fib_1_m_axi_gmem_BREADY,
	fib_1_m_axi_gmem_BVALID,
	fib_1_m_axi_gmem_BID,
	fib_1_m_axi_gmem_BRESP,
	fib_1_m_axi_gmem_BUSER,
	fib_1_s_axi_control_ARREADY,
	fib_1_s_axi_control_ARVALID,
	fib_1_s_axi_control_ARADDR,
	fib_1_s_axi_control_RREADY,
	fib_1_s_axi_control_RVALID,
	fib_1_s_axi_control_RDATA,
	fib_1_s_axi_control_RRESP,
	fib_1_s_axi_control_AWREADY,
	fib_1_s_axi_control_AWVALID,
	fib_1_s_axi_control_AWADDR,
	fib_1_s_axi_control_WREADY,
	fib_1_s_axi_control_WVALID,
	fib_1_s_axi_control_WDATA,
	fib_1_s_axi_control_WSTRB,
	fib_1_s_axi_control_BREADY,
	fib_1_s_axi_control_BVALID,
	fib_1_s_axi_control_BRESP,
	fib_2_m_axi_gmem_ARREADY,
	fib_2_m_axi_gmem_ARVALID,
	fib_2_m_axi_gmem_ARID,
	fib_2_m_axi_gmem_ARADDR,
	fib_2_m_axi_gmem_ARLEN,
	fib_2_m_axi_gmem_ARSIZE,
	fib_2_m_axi_gmem_ARBURST,
	fib_2_m_axi_gmem_ARLOCK,
	fib_2_m_axi_gmem_ARCACHE,
	fib_2_m_axi_gmem_ARPROT,
	fib_2_m_axi_gmem_ARQOS,
	fib_2_m_axi_gmem_ARREGION,
	fib_2_m_axi_gmem_ARUSER,
	fib_2_m_axi_gmem_RREADY,
	fib_2_m_axi_gmem_RVALID,
	fib_2_m_axi_gmem_RID,
	fib_2_m_axi_gmem_RDATA,
	fib_2_m_axi_gmem_RRESP,
	fib_2_m_axi_gmem_RLAST,
	fib_2_m_axi_gmem_RUSER,
	fib_2_m_axi_gmem_AWREADY,
	fib_2_m_axi_gmem_AWVALID,
	fib_2_m_axi_gmem_AWID,
	fib_2_m_axi_gmem_AWADDR,
	fib_2_m_axi_gmem_AWLEN,
	fib_2_m_axi_gmem_AWSIZE,
	fib_2_m_axi_gmem_AWBURST,
	fib_2_m_axi_gmem_AWLOCK,
	fib_2_m_axi_gmem_AWCACHE,
	fib_2_m_axi_gmem_AWPROT,
	fib_2_m_axi_gmem_AWQOS,
	fib_2_m_axi_gmem_AWREGION,
	fib_2_m_axi_gmem_AWUSER,
	fib_2_m_axi_gmem_WREADY,
	fib_2_m_axi_gmem_WVALID,
	fib_2_m_axi_gmem_WDATA,
	fib_2_m_axi_gmem_WSTRB,
	fib_2_m_axi_gmem_WLAST,
	fib_2_m_axi_gmem_WUSER,
	fib_2_m_axi_gmem_BREADY,
	fib_2_m_axi_gmem_BVALID,
	fib_2_m_axi_gmem_BID,
	fib_2_m_axi_gmem_BRESP,
	fib_2_m_axi_gmem_BUSER,
	fib_2_s_axi_control_ARREADY,
	fib_2_s_axi_control_ARVALID,
	fib_2_s_axi_control_ARADDR,
	fib_2_s_axi_control_RREADY,
	fib_2_s_axi_control_RVALID,
	fib_2_s_axi_control_RDATA,
	fib_2_s_axi_control_RRESP,
	fib_2_s_axi_control_AWREADY,
	fib_2_s_axi_control_AWVALID,
	fib_2_s_axi_control_AWADDR,
	fib_2_s_axi_control_WREADY,
	fib_2_s_axi_control_WVALID,
	fib_2_s_axi_control_WDATA,
	fib_2_s_axi_control_WSTRB,
	fib_2_s_axi_control_BREADY,
	fib_2_s_axi_control_BVALID,
	fib_2_s_axi_control_BRESP,
	fib_3_m_axi_gmem_ARREADY,
	fib_3_m_axi_gmem_ARVALID,
	fib_3_m_axi_gmem_ARID,
	fib_3_m_axi_gmem_ARADDR,
	fib_3_m_axi_gmem_ARLEN,
	fib_3_m_axi_gmem_ARSIZE,
	fib_3_m_axi_gmem_ARBURST,
	fib_3_m_axi_gmem_ARLOCK,
	fib_3_m_axi_gmem_ARCACHE,
	fib_3_m_axi_gmem_ARPROT,
	fib_3_m_axi_gmem_ARQOS,
	fib_3_m_axi_gmem_ARREGION,
	fib_3_m_axi_gmem_ARUSER,
	fib_3_m_axi_gmem_RREADY,
	fib_3_m_axi_gmem_RVALID,
	fib_3_m_axi_gmem_RID,
	fib_3_m_axi_gmem_RDATA,
	fib_3_m_axi_gmem_RRESP,
	fib_3_m_axi_gmem_RLAST,
	fib_3_m_axi_gmem_RUSER,
	fib_3_m_axi_gmem_AWREADY,
	fib_3_m_axi_gmem_AWVALID,
	fib_3_m_axi_gmem_AWID,
	fib_3_m_axi_gmem_AWADDR,
	fib_3_m_axi_gmem_AWLEN,
	fib_3_m_axi_gmem_AWSIZE,
	fib_3_m_axi_gmem_AWBURST,
	fib_3_m_axi_gmem_AWLOCK,
	fib_3_m_axi_gmem_AWCACHE,
	fib_3_m_axi_gmem_AWPROT,
	fib_3_m_axi_gmem_AWQOS,
	fib_3_m_axi_gmem_AWREGION,
	fib_3_m_axi_gmem_AWUSER,
	fib_3_m_axi_gmem_WREADY,
	fib_3_m_axi_gmem_WVALID,
	fib_3_m_axi_gmem_WDATA,
	fib_3_m_axi_gmem_WSTRB,
	fib_3_m_axi_gmem_WLAST,
	fib_3_m_axi_gmem_WUSER,
	fib_3_m_axi_gmem_BREADY,
	fib_3_m_axi_gmem_BVALID,
	fib_3_m_axi_gmem_BID,
	fib_3_m_axi_gmem_BRESP,
	fib_3_m_axi_gmem_BUSER,
	fib_3_s_axi_control_ARREADY,
	fib_3_s_axi_control_ARVALID,
	fib_3_s_axi_control_ARADDR,
	fib_3_s_axi_control_RREADY,
	fib_3_s_axi_control_RVALID,
	fib_3_s_axi_control_RDATA,
	fib_3_s_axi_control_RRESP,
	fib_3_s_axi_control_AWREADY,
	fib_3_s_axi_control_AWVALID,
	fib_3_s_axi_control_AWADDR,
	fib_3_s_axi_control_WREADY,
	fib_3_s_axi_control_WVALID,
	fib_3_s_axi_control_WDATA,
	fib_3_s_axi_control_WSTRB,
	fib_3_s_axi_control_BREADY,
	fib_3_s_axi_control_BVALID,
	fib_3_s_axi_control_BRESP,
	fib_4_m_axi_gmem_ARREADY,
	fib_4_m_axi_gmem_ARVALID,
	fib_4_m_axi_gmem_ARID,
	fib_4_m_axi_gmem_ARADDR,
	fib_4_m_axi_gmem_ARLEN,
	fib_4_m_axi_gmem_ARSIZE,
	fib_4_m_axi_gmem_ARBURST,
	fib_4_m_axi_gmem_ARLOCK,
	fib_4_m_axi_gmem_ARCACHE,
	fib_4_m_axi_gmem_ARPROT,
	fib_4_m_axi_gmem_ARQOS,
	fib_4_m_axi_gmem_ARREGION,
	fib_4_m_axi_gmem_ARUSER,
	fib_4_m_axi_gmem_RREADY,
	fib_4_m_axi_gmem_RVALID,
	fib_4_m_axi_gmem_RID,
	fib_4_m_axi_gmem_RDATA,
	fib_4_m_axi_gmem_RRESP,
	fib_4_m_axi_gmem_RLAST,
	fib_4_m_axi_gmem_RUSER,
	fib_4_m_axi_gmem_AWREADY,
	fib_4_m_axi_gmem_AWVALID,
	fib_4_m_axi_gmem_AWID,
	fib_4_m_axi_gmem_AWADDR,
	fib_4_m_axi_gmem_AWLEN,
	fib_4_m_axi_gmem_AWSIZE,
	fib_4_m_axi_gmem_AWBURST,
	fib_4_m_axi_gmem_AWLOCK,
	fib_4_m_axi_gmem_AWCACHE,
	fib_4_m_axi_gmem_AWPROT,
	fib_4_m_axi_gmem_AWQOS,
	fib_4_m_axi_gmem_AWREGION,
	fib_4_m_axi_gmem_AWUSER,
	fib_4_m_axi_gmem_WREADY,
	fib_4_m_axi_gmem_WVALID,
	fib_4_m_axi_gmem_WDATA,
	fib_4_m_axi_gmem_WSTRB,
	fib_4_m_axi_gmem_WLAST,
	fib_4_m_axi_gmem_WUSER,
	fib_4_m_axi_gmem_BREADY,
	fib_4_m_axi_gmem_BVALID,
	fib_4_m_axi_gmem_BID,
	fib_4_m_axi_gmem_BRESP,
	fib_4_m_axi_gmem_BUSER,
	fib_4_s_axi_control_ARREADY,
	fib_4_s_axi_control_ARVALID,
	fib_4_s_axi_control_ARADDR,
	fib_4_s_axi_control_RREADY,
	fib_4_s_axi_control_RVALID,
	fib_4_s_axi_control_RDATA,
	fib_4_s_axi_control_RRESP,
	fib_4_s_axi_control_AWREADY,
	fib_4_s_axi_control_AWVALID,
	fib_4_s_axi_control_AWADDR,
	fib_4_s_axi_control_WREADY,
	fib_4_s_axi_control_WVALID,
	fib_4_s_axi_control_WDATA,
	fib_4_s_axi_control_WSTRB,
	fib_4_s_axi_control_BREADY,
	fib_4_s_axi_control_BVALID,
	fib_4_s_axi_control_BRESP,
	fib_5_m_axi_gmem_ARREADY,
	fib_5_m_axi_gmem_ARVALID,
	fib_5_m_axi_gmem_ARID,
	fib_5_m_axi_gmem_ARADDR,
	fib_5_m_axi_gmem_ARLEN,
	fib_5_m_axi_gmem_ARSIZE,
	fib_5_m_axi_gmem_ARBURST,
	fib_5_m_axi_gmem_ARLOCK,
	fib_5_m_axi_gmem_ARCACHE,
	fib_5_m_axi_gmem_ARPROT,
	fib_5_m_axi_gmem_ARQOS,
	fib_5_m_axi_gmem_ARREGION,
	fib_5_m_axi_gmem_ARUSER,
	fib_5_m_axi_gmem_RREADY,
	fib_5_m_axi_gmem_RVALID,
	fib_5_m_axi_gmem_RID,
	fib_5_m_axi_gmem_RDATA,
	fib_5_m_axi_gmem_RRESP,
	fib_5_m_axi_gmem_RLAST,
	fib_5_m_axi_gmem_RUSER,
	fib_5_m_axi_gmem_AWREADY,
	fib_5_m_axi_gmem_AWVALID,
	fib_5_m_axi_gmem_AWID,
	fib_5_m_axi_gmem_AWADDR,
	fib_5_m_axi_gmem_AWLEN,
	fib_5_m_axi_gmem_AWSIZE,
	fib_5_m_axi_gmem_AWBURST,
	fib_5_m_axi_gmem_AWLOCK,
	fib_5_m_axi_gmem_AWCACHE,
	fib_5_m_axi_gmem_AWPROT,
	fib_5_m_axi_gmem_AWQOS,
	fib_5_m_axi_gmem_AWREGION,
	fib_5_m_axi_gmem_AWUSER,
	fib_5_m_axi_gmem_WREADY,
	fib_5_m_axi_gmem_WVALID,
	fib_5_m_axi_gmem_WDATA,
	fib_5_m_axi_gmem_WSTRB,
	fib_5_m_axi_gmem_WLAST,
	fib_5_m_axi_gmem_WUSER,
	fib_5_m_axi_gmem_BREADY,
	fib_5_m_axi_gmem_BVALID,
	fib_5_m_axi_gmem_BID,
	fib_5_m_axi_gmem_BRESP,
	fib_5_m_axi_gmem_BUSER,
	fib_5_s_axi_control_ARREADY,
	fib_5_s_axi_control_ARVALID,
	fib_5_s_axi_control_ARADDR,
	fib_5_s_axi_control_RREADY,
	fib_5_s_axi_control_RVALID,
	fib_5_s_axi_control_RDATA,
	fib_5_s_axi_control_RRESP,
	fib_5_s_axi_control_AWREADY,
	fib_5_s_axi_control_AWVALID,
	fib_5_s_axi_control_AWADDR,
	fib_5_s_axi_control_WREADY,
	fib_5_s_axi_control_WVALID,
	fib_5_s_axi_control_WDATA,
	fib_5_s_axi_control_WSTRB,
	fib_5_s_axi_control_BREADY,
	fib_5_s_axi_control_BVALID,
	fib_5_s_axi_control_BRESP,
	fib_6_m_axi_gmem_ARREADY,
	fib_6_m_axi_gmem_ARVALID,
	fib_6_m_axi_gmem_ARID,
	fib_6_m_axi_gmem_ARADDR,
	fib_6_m_axi_gmem_ARLEN,
	fib_6_m_axi_gmem_ARSIZE,
	fib_6_m_axi_gmem_ARBURST,
	fib_6_m_axi_gmem_ARLOCK,
	fib_6_m_axi_gmem_ARCACHE,
	fib_6_m_axi_gmem_ARPROT,
	fib_6_m_axi_gmem_ARQOS,
	fib_6_m_axi_gmem_ARREGION,
	fib_6_m_axi_gmem_ARUSER,
	fib_6_m_axi_gmem_RREADY,
	fib_6_m_axi_gmem_RVALID,
	fib_6_m_axi_gmem_RID,
	fib_6_m_axi_gmem_RDATA,
	fib_6_m_axi_gmem_RRESP,
	fib_6_m_axi_gmem_RLAST,
	fib_6_m_axi_gmem_RUSER,
	fib_6_m_axi_gmem_AWREADY,
	fib_6_m_axi_gmem_AWVALID,
	fib_6_m_axi_gmem_AWID,
	fib_6_m_axi_gmem_AWADDR,
	fib_6_m_axi_gmem_AWLEN,
	fib_6_m_axi_gmem_AWSIZE,
	fib_6_m_axi_gmem_AWBURST,
	fib_6_m_axi_gmem_AWLOCK,
	fib_6_m_axi_gmem_AWCACHE,
	fib_6_m_axi_gmem_AWPROT,
	fib_6_m_axi_gmem_AWQOS,
	fib_6_m_axi_gmem_AWREGION,
	fib_6_m_axi_gmem_AWUSER,
	fib_6_m_axi_gmem_WREADY,
	fib_6_m_axi_gmem_WVALID,
	fib_6_m_axi_gmem_WDATA,
	fib_6_m_axi_gmem_WSTRB,
	fib_6_m_axi_gmem_WLAST,
	fib_6_m_axi_gmem_WUSER,
	fib_6_m_axi_gmem_BREADY,
	fib_6_m_axi_gmem_BVALID,
	fib_6_m_axi_gmem_BID,
	fib_6_m_axi_gmem_BRESP,
	fib_6_m_axi_gmem_BUSER,
	fib_6_s_axi_control_ARREADY,
	fib_6_s_axi_control_ARVALID,
	fib_6_s_axi_control_ARADDR,
	fib_6_s_axi_control_RREADY,
	fib_6_s_axi_control_RVALID,
	fib_6_s_axi_control_RDATA,
	fib_6_s_axi_control_RRESP,
	fib_6_s_axi_control_AWREADY,
	fib_6_s_axi_control_AWVALID,
	fib_6_s_axi_control_AWADDR,
	fib_6_s_axi_control_WREADY,
	fib_6_s_axi_control_WVALID,
	fib_6_s_axi_control_WDATA,
	fib_6_s_axi_control_WSTRB,
	fib_6_s_axi_control_BREADY,
	fib_6_s_axi_control_BVALID,
	fib_6_s_axi_control_BRESP,
	fib_7_m_axi_gmem_ARREADY,
	fib_7_m_axi_gmem_ARVALID,
	fib_7_m_axi_gmem_ARID,
	fib_7_m_axi_gmem_ARADDR,
	fib_7_m_axi_gmem_ARLEN,
	fib_7_m_axi_gmem_ARSIZE,
	fib_7_m_axi_gmem_ARBURST,
	fib_7_m_axi_gmem_ARLOCK,
	fib_7_m_axi_gmem_ARCACHE,
	fib_7_m_axi_gmem_ARPROT,
	fib_7_m_axi_gmem_ARQOS,
	fib_7_m_axi_gmem_ARREGION,
	fib_7_m_axi_gmem_ARUSER,
	fib_7_m_axi_gmem_RREADY,
	fib_7_m_axi_gmem_RVALID,
	fib_7_m_axi_gmem_RID,
	fib_7_m_axi_gmem_RDATA,
	fib_7_m_axi_gmem_RRESP,
	fib_7_m_axi_gmem_RLAST,
	fib_7_m_axi_gmem_RUSER,
	fib_7_m_axi_gmem_AWREADY,
	fib_7_m_axi_gmem_AWVALID,
	fib_7_m_axi_gmem_AWID,
	fib_7_m_axi_gmem_AWADDR,
	fib_7_m_axi_gmem_AWLEN,
	fib_7_m_axi_gmem_AWSIZE,
	fib_7_m_axi_gmem_AWBURST,
	fib_7_m_axi_gmem_AWLOCK,
	fib_7_m_axi_gmem_AWCACHE,
	fib_7_m_axi_gmem_AWPROT,
	fib_7_m_axi_gmem_AWQOS,
	fib_7_m_axi_gmem_AWREGION,
	fib_7_m_axi_gmem_AWUSER,
	fib_7_m_axi_gmem_WREADY,
	fib_7_m_axi_gmem_WVALID,
	fib_7_m_axi_gmem_WDATA,
	fib_7_m_axi_gmem_WSTRB,
	fib_7_m_axi_gmem_WLAST,
	fib_7_m_axi_gmem_WUSER,
	fib_7_m_axi_gmem_BREADY,
	fib_7_m_axi_gmem_BVALID,
	fib_7_m_axi_gmem_BID,
	fib_7_m_axi_gmem_BRESP,
	fib_7_m_axi_gmem_BUSER,
	fib_7_s_axi_control_ARREADY,
	fib_7_s_axi_control_ARVALID,
	fib_7_s_axi_control_ARADDR,
	fib_7_s_axi_control_RREADY,
	fib_7_s_axi_control_RVALID,
	fib_7_s_axi_control_RDATA,
	fib_7_s_axi_control_RRESP,
	fib_7_s_axi_control_AWREADY,
	fib_7_s_axi_control_AWVALID,
	fib_7_s_axi_control_AWADDR,
	fib_7_s_axi_control_WREADY,
	fib_7_s_axi_control_WVALID,
	fib_7_s_axi_control_WDATA,
	fib_7_s_axi_control_WSTRB,
	fib_7_s_axi_control_BREADY,
	fib_7_s_axi_control_BVALID,
	fib_7_s_axi_control_BRESP,
	fib_8_m_axi_gmem_ARREADY,
	fib_8_m_axi_gmem_ARVALID,
	fib_8_m_axi_gmem_ARID,
	fib_8_m_axi_gmem_ARADDR,
	fib_8_m_axi_gmem_ARLEN,
	fib_8_m_axi_gmem_ARSIZE,
	fib_8_m_axi_gmem_ARBURST,
	fib_8_m_axi_gmem_ARLOCK,
	fib_8_m_axi_gmem_ARCACHE,
	fib_8_m_axi_gmem_ARPROT,
	fib_8_m_axi_gmem_ARQOS,
	fib_8_m_axi_gmem_ARREGION,
	fib_8_m_axi_gmem_ARUSER,
	fib_8_m_axi_gmem_RREADY,
	fib_8_m_axi_gmem_RVALID,
	fib_8_m_axi_gmem_RID,
	fib_8_m_axi_gmem_RDATA,
	fib_8_m_axi_gmem_RRESP,
	fib_8_m_axi_gmem_RLAST,
	fib_8_m_axi_gmem_RUSER,
	fib_8_m_axi_gmem_AWREADY,
	fib_8_m_axi_gmem_AWVALID,
	fib_8_m_axi_gmem_AWID,
	fib_8_m_axi_gmem_AWADDR,
	fib_8_m_axi_gmem_AWLEN,
	fib_8_m_axi_gmem_AWSIZE,
	fib_8_m_axi_gmem_AWBURST,
	fib_8_m_axi_gmem_AWLOCK,
	fib_8_m_axi_gmem_AWCACHE,
	fib_8_m_axi_gmem_AWPROT,
	fib_8_m_axi_gmem_AWQOS,
	fib_8_m_axi_gmem_AWREGION,
	fib_8_m_axi_gmem_AWUSER,
	fib_8_m_axi_gmem_WREADY,
	fib_8_m_axi_gmem_WVALID,
	fib_8_m_axi_gmem_WDATA,
	fib_8_m_axi_gmem_WSTRB,
	fib_8_m_axi_gmem_WLAST,
	fib_8_m_axi_gmem_WUSER,
	fib_8_m_axi_gmem_BREADY,
	fib_8_m_axi_gmem_BVALID,
	fib_8_m_axi_gmem_BID,
	fib_8_m_axi_gmem_BRESP,
	fib_8_m_axi_gmem_BUSER,
	fib_8_s_axi_control_ARREADY,
	fib_8_s_axi_control_ARVALID,
	fib_8_s_axi_control_ARADDR,
	fib_8_s_axi_control_RREADY,
	fib_8_s_axi_control_RVALID,
	fib_8_s_axi_control_RDATA,
	fib_8_s_axi_control_RRESP,
	fib_8_s_axi_control_AWREADY,
	fib_8_s_axi_control_AWVALID,
	fib_8_s_axi_control_AWADDR,
	fib_8_s_axi_control_WREADY,
	fib_8_s_axi_control_WVALID,
	fib_8_s_axi_control_WDATA,
	fib_8_s_axi_control_WSTRB,
	fib_8_s_axi_control_BREADY,
	fib_8_s_axi_control_BVALID,
	fib_8_s_axi_control_BRESP,
	fib_9_m_axi_gmem_ARREADY,
	fib_9_m_axi_gmem_ARVALID,
	fib_9_m_axi_gmem_ARID,
	fib_9_m_axi_gmem_ARADDR,
	fib_9_m_axi_gmem_ARLEN,
	fib_9_m_axi_gmem_ARSIZE,
	fib_9_m_axi_gmem_ARBURST,
	fib_9_m_axi_gmem_ARLOCK,
	fib_9_m_axi_gmem_ARCACHE,
	fib_9_m_axi_gmem_ARPROT,
	fib_9_m_axi_gmem_ARQOS,
	fib_9_m_axi_gmem_ARREGION,
	fib_9_m_axi_gmem_ARUSER,
	fib_9_m_axi_gmem_RREADY,
	fib_9_m_axi_gmem_RVALID,
	fib_9_m_axi_gmem_RID,
	fib_9_m_axi_gmem_RDATA,
	fib_9_m_axi_gmem_RRESP,
	fib_9_m_axi_gmem_RLAST,
	fib_9_m_axi_gmem_RUSER,
	fib_9_m_axi_gmem_AWREADY,
	fib_9_m_axi_gmem_AWVALID,
	fib_9_m_axi_gmem_AWID,
	fib_9_m_axi_gmem_AWADDR,
	fib_9_m_axi_gmem_AWLEN,
	fib_9_m_axi_gmem_AWSIZE,
	fib_9_m_axi_gmem_AWBURST,
	fib_9_m_axi_gmem_AWLOCK,
	fib_9_m_axi_gmem_AWCACHE,
	fib_9_m_axi_gmem_AWPROT,
	fib_9_m_axi_gmem_AWQOS,
	fib_9_m_axi_gmem_AWREGION,
	fib_9_m_axi_gmem_AWUSER,
	fib_9_m_axi_gmem_WREADY,
	fib_9_m_axi_gmem_WVALID,
	fib_9_m_axi_gmem_WDATA,
	fib_9_m_axi_gmem_WSTRB,
	fib_9_m_axi_gmem_WLAST,
	fib_9_m_axi_gmem_WUSER,
	fib_9_m_axi_gmem_BREADY,
	fib_9_m_axi_gmem_BVALID,
	fib_9_m_axi_gmem_BID,
	fib_9_m_axi_gmem_BRESP,
	fib_9_m_axi_gmem_BUSER,
	fib_9_s_axi_control_ARREADY,
	fib_9_s_axi_control_ARVALID,
	fib_9_s_axi_control_ARADDR,
	fib_9_s_axi_control_RREADY,
	fib_9_s_axi_control_RVALID,
	fib_9_s_axi_control_RDATA,
	fib_9_s_axi_control_RRESP,
	fib_9_s_axi_control_AWREADY,
	fib_9_s_axi_control_AWVALID,
	fib_9_s_axi_control_AWADDR,
	fib_9_s_axi_control_WREADY,
	fib_9_s_axi_control_WVALID,
	fib_9_s_axi_control_WDATA,
	fib_9_s_axi_control_WSTRB,
	fib_9_s_axi_control_BREADY,
	fib_9_s_axi_control_BVALID,
	fib_9_s_axi_control_BRESP,
	fib_10_m_axi_gmem_ARREADY,
	fib_10_m_axi_gmem_ARVALID,
	fib_10_m_axi_gmem_ARID,
	fib_10_m_axi_gmem_ARADDR,
	fib_10_m_axi_gmem_ARLEN,
	fib_10_m_axi_gmem_ARSIZE,
	fib_10_m_axi_gmem_ARBURST,
	fib_10_m_axi_gmem_ARLOCK,
	fib_10_m_axi_gmem_ARCACHE,
	fib_10_m_axi_gmem_ARPROT,
	fib_10_m_axi_gmem_ARQOS,
	fib_10_m_axi_gmem_ARREGION,
	fib_10_m_axi_gmem_ARUSER,
	fib_10_m_axi_gmem_RREADY,
	fib_10_m_axi_gmem_RVALID,
	fib_10_m_axi_gmem_RID,
	fib_10_m_axi_gmem_RDATA,
	fib_10_m_axi_gmem_RRESP,
	fib_10_m_axi_gmem_RLAST,
	fib_10_m_axi_gmem_RUSER,
	fib_10_m_axi_gmem_AWREADY,
	fib_10_m_axi_gmem_AWVALID,
	fib_10_m_axi_gmem_AWID,
	fib_10_m_axi_gmem_AWADDR,
	fib_10_m_axi_gmem_AWLEN,
	fib_10_m_axi_gmem_AWSIZE,
	fib_10_m_axi_gmem_AWBURST,
	fib_10_m_axi_gmem_AWLOCK,
	fib_10_m_axi_gmem_AWCACHE,
	fib_10_m_axi_gmem_AWPROT,
	fib_10_m_axi_gmem_AWQOS,
	fib_10_m_axi_gmem_AWREGION,
	fib_10_m_axi_gmem_AWUSER,
	fib_10_m_axi_gmem_WREADY,
	fib_10_m_axi_gmem_WVALID,
	fib_10_m_axi_gmem_WDATA,
	fib_10_m_axi_gmem_WSTRB,
	fib_10_m_axi_gmem_WLAST,
	fib_10_m_axi_gmem_WUSER,
	fib_10_m_axi_gmem_BREADY,
	fib_10_m_axi_gmem_BVALID,
	fib_10_m_axi_gmem_BID,
	fib_10_m_axi_gmem_BRESP,
	fib_10_m_axi_gmem_BUSER,
	fib_10_s_axi_control_ARREADY,
	fib_10_s_axi_control_ARVALID,
	fib_10_s_axi_control_ARADDR,
	fib_10_s_axi_control_RREADY,
	fib_10_s_axi_control_RVALID,
	fib_10_s_axi_control_RDATA,
	fib_10_s_axi_control_RRESP,
	fib_10_s_axi_control_AWREADY,
	fib_10_s_axi_control_AWVALID,
	fib_10_s_axi_control_AWADDR,
	fib_10_s_axi_control_WREADY,
	fib_10_s_axi_control_WVALID,
	fib_10_s_axi_control_WDATA,
	fib_10_s_axi_control_WSTRB,
	fib_10_s_axi_control_BREADY,
	fib_10_s_axi_control_BVALID,
	fib_10_s_axi_control_BRESP,
	fib_11_m_axi_gmem_ARREADY,
	fib_11_m_axi_gmem_ARVALID,
	fib_11_m_axi_gmem_ARID,
	fib_11_m_axi_gmem_ARADDR,
	fib_11_m_axi_gmem_ARLEN,
	fib_11_m_axi_gmem_ARSIZE,
	fib_11_m_axi_gmem_ARBURST,
	fib_11_m_axi_gmem_ARLOCK,
	fib_11_m_axi_gmem_ARCACHE,
	fib_11_m_axi_gmem_ARPROT,
	fib_11_m_axi_gmem_ARQOS,
	fib_11_m_axi_gmem_ARREGION,
	fib_11_m_axi_gmem_ARUSER,
	fib_11_m_axi_gmem_RREADY,
	fib_11_m_axi_gmem_RVALID,
	fib_11_m_axi_gmem_RID,
	fib_11_m_axi_gmem_RDATA,
	fib_11_m_axi_gmem_RRESP,
	fib_11_m_axi_gmem_RLAST,
	fib_11_m_axi_gmem_RUSER,
	fib_11_m_axi_gmem_AWREADY,
	fib_11_m_axi_gmem_AWVALID,
	fib_11_m_axi_gmem_AWID,
	fib_11_m_axi_gmem_AWADDR,
	fib_11_m_axi_gmem_AWLEN,
	fib_11_m_axi_gmem_AWSIZE,
	fib_11_m_axi_gmem_AWBURST,
	fib_11_m_axi_gmem_AWLOCK,
	fib_11_m_axi_gmem_AWCACHE,
	fib_11_m_axi_gmem_AWPROT,
	fib_11_m_axi_gmem_AWQOS,
	fib_11_m_axi_gmem_AWREGION,
	fib_11_m_axi_gmem_AWUSER,
	fib_11_m_axi_gmem_WREADY,
	fib_11_m_axi_gmem_WVALID,
	fib_11_m_axi_gmem_WDATA,
	fib_11_m_axi_gmem_WSTRB,
	fib_11_m_axi_gmem_WLAST,
	fib_11_m_axi_gmem_WUSER,
	fib_11_m_axi_gmem_BREADY,
	fib_11_m_axi_gmem_BVALID,
	fib_11_m_axi_gmem_BID,
	fib_11_m_axi_gmem_BRESP,
	fib_11_m_axi_gmem_BUSER,
	fib_11_s_axi_control_ARREADY,
	fib_11_s_axi_control_ARVALID,
	fib_11_s_axi_control_ARADDR,
	fib_11_s_axi_control_RREADY,
	fib_11_s_axi_control_RVALID,
	fib_11_s_axi_control_RDATA,
	fib_11_s_axi_control_RRESP,
	fib_11_s_axi_control_AWREADY,
	fib_11_s_axi_control_AWVALID,
	fib_11_s_axi_control_AWADDR,
	fib_11_s_axi_control_WREADY,
	fib_11_s_axi_control_WVALID,
	fib_11_s_axi_control_WDATA,
	fib_11_s_axi_control_WSTRB,
	fib_11_s_axi_control_BREADY,
	fib_11_s_axi_control_BVALID,
	fib_11_s_axi_control_BRESP,
	fib_12_m_axi_gmem_ARREADY,
	fib_12_m_axi_gmem_ARVALID,
	fib_12_m_axi_gmem_ARID,
	fib_12_m_axi_gmem_ARADDR,
	fib_12_m_axi_gmem_ARLEN,
	fib_12_m_axi_gmem_ARSIZE,
	fib_12_m_axi_gmem_ARBURST,
	fib_12_m_axi_gmem_ARLOCK,
	fib_12_m_axi_gmem_ARCACHE,
	fib_12_m_axi_gmem_ARPROT,
	fib_12_m_axi_gmem_ARQOS,
	fib_12_m_axi_gmem_ARREGION,
	fib_12_m_axi_gmem_ARUSER,
	fib_12_m_axi_gmem_RREADY,
	fib_12_m_axi_gmem_RVALID,
	fib_12_m_axi_gmem_RID,
	fib_12_m_axi_gmem_RDATA,
	fib_12_m_axi_gmem_RRESP,
	fib_12_m_axi_gmem_RLAST,
	fib_12_m_axi_gmem_RUSER,
	fib_12_m_axi_gmem_AWREADY,
	fib_12_m_axi_gmem_AWVALID,
	fib_12_m_axi_gmem_AWID,
	fib_12_m_axi_gmem_AWADDR,
	fib_12_m_axi_gmem_AWLEN,
	fib_12_m_axi_gmem_AWSIZE,
	fib_12_m_axi_gmem_AWBURST,
	fib_12_m_axi_gmem_AWLOCK,
	fib_12_m_axi_gmem_AWCACHE,
	fib_12_m_axi_gmem_AWPROT,
	fib_12_m_axi_gmem_AWQOS,
	fib_12_m_axi_gmem_AWREGION,
	fib_12_m_axi_gmem_AWUSER,
	fib_12_m_axi_gmem_WREADY,
	fib_12_m_axi_gmem_WVALID,
	fib_12_m_axi_gmem_WDATA,
	fib_12_m_axi_gmem_WSTRB,
	fib_12_m_axi_gmem_WLAST,
	fib_12_m_axi_gmem_WUSER,
	fib_12_m_axi_gmem_BREADY,
	fib_12_m_axi_gmem_BVALID,
	fib_12_m_axi_gmem_BID,
	fib_12_m_axi_gmem_BRESP,
	fib_12_m_axi_gmem_BUSER,
	fib_12_s_axi_control_ARREADY,
	fib_12_s_axi_control_ARVALID,
	fib_12_s_axi_control_ARADDR,
	fib_12_s_axi_control_RREADY,
	fib_12_s_axi_control_RVALID,
	fib_12_s_axi_control_RDATA,
	fib_12_s_axi_control_RRESP,
	fib_12_s_axi_control_AWREADY,
	fib_12_s_axi_control_AWVALID,
	fib_12_s_axi_control_AWADDR,
	fib_12_s_axi_control_WREADY,
	fib_12_s_axi_control_WVALID,
	fib_12_s_axi_control_WDATA,
	fib_12_s_axi_control_WSTRB,
	fib_12_s_axi_control_BREADY,
	fib_12_s_axi_control_BVALID,
	fib_12_s_axi_control_BRESP,
	fib_13_m_axi_gmem_ARREADY,
	fib_13_m_axi_gmem_ARVALID,
	fib_13_m_axi_gmem_ARID,
	fib_13_m_axi_gmem_ARADDR,
	fib_13_m_axi_gmem_ARLEN,
	fib_13_m_axi_gmem_ARSIZE,
	fib_13_m_axi_gmem_ARBURST,
	fib_13_m_axi_gmem_ARLOCK,
	fib_13_m_axi_gmem_ARCACHE,
	fib_13_m_axi_gmem_ARPROT,
	fib_13_m_axi_gmem_ARQOS,
	fib_13_m_axi_gmem_ARREGION,
	fib_13_m_axi_gmem_ARUSER,
	fib_13_m_axi_gmem_RREADY,
	fib_13_m_axi_gmem_RVALID,
	fib_13_m_axi_gmem_RID,
	fib_13_m_axi_gmem_RDATA,
	fib_13_m_axi_gmem_RRESP,
	fib_13_m_axi_gmem_RLAST,
	fib_13_m_axi_gmem_RUSER,
	fib_13_m_axi_gmem_AWREADY,
	fib_13_m_axi_gmem_AWVALID,
	fib_13_m_axi_gmem_AWID,
	fib_13_m_axi_gmem_AWADDR,
	fib_13_m_axi_gmem_AWLEN,
	fib_13_m_axi_gmem_AWSIZE,
	fib_13_m_axi_gmem_AWBURST,
	fib_13_m_axi_gmem_AWLOCK,
	fib_13_m_axi_gmem_AWCACHE,
	fib_13_m_axi_gmem_AWPROT,
	fib_13_m_axi_gmem_AWQOS,
	fib_13_m_axi_gmem_AWREGION,
	fib_13_m_axi_gmem_AWUSER,
	fib_13_m_axi_gmem_WREADY,
	fib_13_m_axi_gmem_WVALID,
	fib_13_m_axi_gmem_WDATA,
	fib_13_m_axi_gmem_WSTRB,
	fib_13_m_axi_gmem_WLAST,
	fib_13_m_axi_gmem_WUSER,
	fib_13_m_axi_gmem_BREADY,
	fib_13_m_axi_gmem_BVALID,
	fib_13_m_axi_gmem_BID,
	fib_13_m_axi_gmem_BRESP,
	fib_13_m_axi_gmem_BUSER,
	fib_13_s_axi_control_ARREADY,
	fib_13_s_axi_control_ARVALID,
	fib_13_s_axi_control_ARADDR,
	fib_13_s_axi_control_RREADY,
	fib_13_s_axi_control_RVALID,
	fib_13_s_axi_control_RDATA,
	fib_13_s_axi_control_RRESP,
	fib_13_s_axi_control_AWREADY,
	fib_13_s_axi_control_AWVALID,
	fib_13_s_axi_control_AWADDR,
	fib_13_s_axi_control_WREADY,
	fib_13_s_axi_control_WVALID,
	fib_13_s_axi_control_WDATA,
	fib_13_s_axi_control_WSTRB,
	fib_13_s_axi_control_BREADY,
	fib_13_s_axi_control_BVALID,
	fib_13_s_axi_control_BRESP,
	fib_14_m_axi_gmem_ARREADY,
	fib_14_m_axi_gmem_ARVALID,
	fib_14_m_axi_gmem_ARID,
	fib_14_m_axi_gmem_ARADDR,
	fib_14_m_axi_gmem_ARLEN,
	fib_14_m_axi_gmem_ARSIZE,
	fib_14_m_axi_gmem_ARBURST,
	fib_14_m_axi_gmem_ARLOCK,
	fib_14_m_axi_gmem_ARCACHE,
	fib_14_m_axi_gmem_ARPROT,
	fib_14_m_axi_gmem_ARQOS,
	fib_14_m_axi_gmem_ARREGION,
	fib_14_m_axi_gmem_ARUSER,
	fib_14_m_axi_gmem_RREADY,
	fib_14_m_axi_gmem_RVALID,
	fib_14_m_axi_gmem_RID,
	fib_14_m_axi_gmem_RDATA,
	fib_14_m_axi_gmem_RRESP,
	fib_14_m_axi_gmem_RLAST,
	fib_14_m_axi_gmem_RUSER,
	fib_14_m_axi_gmem_AWREADY,
	fib_14_m_axi_gmem_AWVALID,
	fib_14_m_axi_gmem_AWID,
	fib_14_m_axi_gmem_AWADDR,
	fib_14_m_axi_gmem_AWLEN,
	fib_14_m_axi_gmem_AWSIZE,
	fib_14_m_axi_gmem_AWBURST,
	fib_14_m_axi_gmem_AWLOCK,
	fib_14_m_axi_gmem_AWCACHE,
	fib_14_m_axi_gmem_AWPROT,
	fib_14_m_axi_gmem_AWQOS,
	fib_14_m_axi_gmem_AWREGION,
	fib_14_m_axi_gmem_AWUSER,
	fib_14_m_axi_gmem_WREADY,
	fib_14_m_axi_gmem_WVALID,
	fib_14_m_axi_gmem_WDATA,
	fib_14_m_axi_gmem_WSTRB,
	fib_14_m_axi_gmem_WLAST,
	fib_14_m_axi_gmem_WUSER,
	fib_14_m_axi_gmem_BREADY,
	fib_14_m_axi_gmem_BVALID,
	fib_14_m_axi_gmem_BID,
	fib_14_m_axi_gmem_BRESP,
	fib_14_m_axi_gmem_BUSER,
	fib_14_s_axi_control_ARREADY,
	fib_14_s_axi_control_ARVALID,
	fib_14_s_axi_control_ARADDR,
	fib_14_s_axi_control_RREADY,
	fib_14_s_axi_control_RVALID,
	fib_14_s_axi_control_RDATA,
	fib_14_s_axi_control_RRESP,
	fib_14_s_axi_control_AWREADY,
	fib_14_s_axi_control_AWVALID,
	fib_14_s_axi_control_AWADDR,
	fib_14_s_axi_control_WREADY,
	fib_14_s_axi_control_WVALID,
	fib_14_s_axi_control_WDATA,
	fib_14_s_axi_control_WSTRB,
	fib_14_s_axi_control_BREADY,
	fib_14_s_axi_control_BVALID,
	fib_14_s_axi_control_BRESP,
	fib_15_m_axi_gmem_ARREADY,
	fib_15_m_axi_gmem_ARVALID,
	fib_15_m_axi_gmem_ARID,
	fib_15_m_axi_gmem_ARADDR,
	fib_15_m_axi_gmem_ARLEN,
	fib_15_m_axi_gmem_ARSIZE,
	fib_15_m_axi_gmem_ARBURST,
	fib_15_m_axi_gmem_ARLOCK,
	fib_15_m_axi_gmem_ARCACHE,
	fib_15_m_axi_gmem_ARPROT,
	fib_15_m_axi_gmem_ARQOS,
	fib_15_m_axi_gmem_ARREGION,
	fib_15_m_axi_gmem_ARUSER,
	fib_15_m_axi_gmem_RREADY,
	fib_15_m_axi_gmem_RVALID,
	fib_15_m_axi_gmem_RID,
	fib_15_m_axi_gmem_RDATA,
	fib_15_m_axi_gmem_RRESP,
	fib_15_m_axi_gmem_RLAST,
	fib_15_m_axi_gmem_RUSER,
	fib_15_m_axi_gmem_AWREADY,
	fib_15_m_axi_gmem_AWVALID,
	fib_15_m_axi_gmem_AWID,
	fib_15_m_axi_gmem_AWADDR,
	fib_15_m_axi_gmem_AWLEN,
	fib_15_m_axi_gmem_AWSIZE,
	fib_15_m_axi_gmem_AWBURST,
	fib_15_m_axi_gmem_AWLOCK,
	fib_15_m_axi_gmem_AWCACHE,
	fib_15_m_axi_gmem_AWPROT,
	fib_15_m_axi_gmem_AWQOS,
	fib_15_m_axi_gmem_AWREGION,
	fib_15_m_axi_gmem_AWUSER,
	fib_15_m_axi_gmem_WREADY,
	fib_15_m_axi_gmem_WVALID,
	fib_15_m_axi_gmem_WDATA,
	fib_15_m_axi_gmem_WSTRB,
	fib_15_m_axi_gmem_WLAST,
	fib_15_m_axi_gmem_WUSER,
	fib_15_m_axi_gmem_BREADY,
	fib_15_m_axi_gmem_BVALID,
	fib_15_m_axi_gmem_BID,
	fib_15_m_axi_gmem_BRESP,
	fib_15_m_axi_gmem_BUSER,
	fib_15_s_axi_control_ARREADY,
	fib_15_s_axi_control_ARVALID,
	fib_15_s_axi_control_ARADDR,
	fib_15_s_axi_control_RREADY,
	fib_15_s_axi_control_RVALID,
	fib_15_s_axi_control_RDATA,
	fib_15_s_axi_control_RRESP,
	fib_15_s_axi_control_AWREADY,
	fib_15_s_axi_control_AWVALID,
	fib_15_s_axi_control_AWADDR,
	fib_15_s_axi_control_WREADY,
	fib_15_s_axi_control_WVALID,
	fib_15_s_axi_control_WDATA,
	fib_15_s_axi_control_WSTRB,
	fib_15_s_axi_control_BREADY,
	fib_15_s_axi_control_BVALID,
	fib_15_s_axi_control_BRESP,
	fib_16_m_axi_gmem_ARREADY,
	fib_16_m_axi_gmem_ARVALID,
	fib_16_m_axi_gmem_ARID,
	fib_16_m_axi_gmem_ARADDR,
	fib_16_m_axi_gmem_ARLEN,
	fib_16_m_axi_gmem_ARSIZE,
	fib_16_m_axi_gmem_ARBURST,
	fib_16_m_axi_gmem_ARLOCK,
	fib_16_m_axi_gmem_ARCACHE,
	fib_16_m_axi_gmem_ARPROT,
	fib_16_m_axi_gmem_ARQOS,
	fib_16_m_axi_gmem_ARREGION,
	fib_16_m_axi_gmem_ARUSER,
	fib_16_m_axi_gmem_RREADY,
	fib_16_m_axi_gmem_RVALID,
	fib_16_m_axi_gmem_RID,
	fib_16_m_axi_gmem_RDATA,
	fib_16_m_axi_gmem_RRESP,
	fib_16_m_axi_gmem_RLAST,
	fib_16_m_axi_gmem_RUSER,
	fib_16_m_axi_gmem_AWREADY,
	fib_16_m_axi_gmem_AWVALID,
	fib_16_m_axi_gmem_AWID,
	fib_16_m_axi_gmem_AWADDR,
	fib_16_m_axi_gmem_AWLEN,
	fib_16_m_axi_gmem_AWSIZE,
	fib_16_m_axi_gmem_AWBURST,
	fib_16_m_axi_gmem_AWLOCK,
	fib_16_m_axi_gmem_AWCACHE,
	fib_16_m_axi_gmem_AWPROT,
	fib_16_m_axi_gmem_AWQOS,
	fib_16_m_axi_gmem_AWREGION,
	fib_16_m_axi_gmem_AWUSER,
	fib_16_m_axi_gmem_WREADY,
	fib_16_m_axi_gmem_WVALID,
	fib_16_m_axi_gmem_WDATA,
	fib_16_m_axi_gmem_WSTRB,
	fib_16_m_axi_gmem_WLAST,
	fib_16_m_axi_gmem_WUSER,
	fib_16_m_axi_gmem_BREADY,
	fib_16_m_axi_gmem_BVALID,
	fib_16_m_axi_gmem_BID,
	fib_16_m_axi_gmem_BRESP,
	fib_16_m_axi_gmem_BUSER,
	fib_16_s_axi_control_ARREADY,
	fib_16_s_axi_control_ARVALID,
	fib_16_s_axi_control_ARADDR,
	fib_16_s_axi_control_RREADY,
	fib_16_s_axi_control_RVALID,
	fib_16_s_axi_control_RDATA,
	fib_16_s_axi_control_RRESP,
	fib_16_s_axi_control_AWREADY,
	fib_16_s_axi_control_AWVALID,
	fib_16_s_axi_control_AWADDR,
	fib_16_s_axi_control_WREADY,
	fib_16_s_axi_control_WVALID,
	fib_16_s_axi_control_WDATA,
	fib_16_s_axi_control_WSTRB,
	fib_16_s_axi_control_BREADY,
	fib_16_s_axi_control_BVALID,
	fib_16_s_axi_control_BRESP,
	fib_17_m_axi_gmem_ARREADY,
	fib_17_m_axi_gmem_ARVALID,
	fib_17_m_axi_gmem_ARID,
	fib_17_m_axi_gmem_ARADDR,
	fib_17_m_axi_gmem_ARLEN,
	fib_17_m_axi_gmem_ARSIZE,
	fib_17_m_axi_gmem_ARBURST,
	fib_17_m_axi_gmem_ARLOCK,
	fib_17_m_axi_gmem_ARCACHE,
	fib_17_m_axi_gmem_ARPROT,
	fib_17_m_axi_gmem_ARQOS,
	fib_17_m_axi_gmem_ARREGION,
	fib_17_m_axi_gmem_ARUSER,
	fib_17_m_axi_gmem_RREADY,
	fib_17_m_axi_gmem_RVALID,
	fib_17_m_axi_gmem_RID,
	fib_17_m_axi_gmem_RDATA,
	fib_17_m_axi_gmem_RRESP,
	fib_17_m_axi_gmem_RLAST,
	fib_17_m_axi_gmem_RUSER,
	fib_17_m_axi_gmem_AWREADY,
	fib_17_m_axi_gmem_AWVALID,
	fib_17_m_axi_gmem_AWID,
	fib_17_m_axi_gmem_AWADDR,
	fib_17_m_axi_gmem_AWLEN,
	fib_17_m_axi_gmem_AWSIZE,
	fib_17_m_axi_gmem_AWBURST,
	fib_17_m_axi_gmem_AWLOCK,
	fib_17_m_axi_gmem_AWCACHE,
	fib_17_m_axi_gmem_AWPROT,
	fib_17_m_axi_gmem_AWQOS,
	fib_17_m_axi_gmem_AWREGION,
	fib_17_m_axi_gmem_AWUSER,
	fib_17_m_axi_gmem_WREADY,
	fib_17_m_axi_gmem_WVALID,
	fib_17_m_axi_gmem_WDATA,
	fib_17_m_axi_gmem_WSTRB,
	fib_17_m_axi_gmem_WLAST,
	fib_17_m_axi_gmem_WUSER,
	fib_17_m_axi_gmem_BREADY,
	fib_17_m_axi_gmem_BVALID,
	fib_17_m_axi_gmem_BID,
	fib_17_m_axi_gmem_BRESP,
	fib_17_m_axi_gmem_BUSER,
	fib_17_s_axi_control_ARREADY,
	fib_17_s_axi_control_ARVALID,
	fib_17_s_axi_control_ARADDR,
	fib_17_s_axi_control_RREADY,
	fib_17_s_axi_control_RVALID,
	fib_17_s_axi_control_RDATA,
	fib_17_s_axi_control_RRESP,
	fib_17_s_axi_control_AWREADY,
	fib_17_s_axi_control_AWVALID,
	fib_17_s_axi_control_AWADDR,
	fib_17_s_axi_control_WREADY,
	fib_17_s_axi_control_WVALID,
	fib_17_s_axi_control_WDATA,
	fib_17_s_axi_control_WSTRB,
	fib_17_s_axi_control_BREADY,
	fib_17_s_axi_control_BVALID,
	fib_17_s_axi_control_BRESP,
	fib_18_m_axi_gmem_ARREADY,
	fib_18_m_axi_gmem_ARVALID,
	fib_18_m_axi_gmem_ARID,
	fib_18_m_axi_gmem_ARADDR,
	fib_18_m_axi_gmem_ARLEN,
	fib_18_m_axi_gmem_ARSIZE,
	fib_18_m_axi_gmem_ARBURST,
	fib_18_m_axi_gmem_ARLOCK,
	fib_18_m_axi_gmem_ARCACHE,
	fib_18_m_axi_gmem_ARPROT,
	fib_18_m_axi_gmem_ARQOS,
	fib_18_m_axi_gmem_ARREGION,
	fib_18_m_axi_gmem_ARUSER,
	fib_18_m_axi_gmem_RREADY,
	fib_18_m_axi_gmem_RVALID,
	fib_18_m_axi_gmem_RID,
	fib_18_m_axi_gmem_RDATA,
	fib_18_m_axi_gmem_RRESP,
	fib_18_m_axi_gmem_RLAST,
	fib_18_m_axi_gmem_RUSER,
	fib_18_m_axi_gmem_AWREADY,
	fib_18_m_axi_gmem_AWVALID,
	fib_18_m_axi_gmem_AWID,
	fib_18_m_axi_gmem_AWADDR,
	fib_18_m_axi_gmem_AWLEN,
	fib_18_m_axi_gmem_AWSIZE,
	fib_18_m_axi_gmem_AWBURST,
	fib_18_m_axi_gmem_AWLOCK,
	fib_18_m_axi_gmem_AWCACHE,
	fib_18_m_axi_gmem_AWPROT,
	fib_18_m_axi_gmem_AWQOS,
	fib_18_m_axi_gmem_AWREGION,
	fib_18_m_axi_gmem_AWUSER,
	fib_18_m_axi_gmem_WREADY,
	fib_18_m_axi_gmem_WVALID,
	fib_18_m_axi_gmem_WDATA,
	fib_18_m_axi_gmem_WSTRB,
	fib_18_m_axi_gmem_WLAST,
	fib_18_m_axi_gmem_WUSER,
	fib_18_m_axi_gmem_BREADY,
	fib_18_m_axi_gmem_BVALID,
	fib_18_m_axi_gmem_BID,
	fib_18_m_axi_gmem_BRESP,
	fib_18_m_axi_gmem_BUSER,
	fib_18_s_axi_control_ARREADY,
	fib_18_s_axi_control_ARVALID,
	fib_18_s_axi_control_ARADDR,
	fib_18_s_axi_control_RREADY,
	fib_18_s_axi_control_RVALID,
	fib_18_s_axi_control_RDATA,
	fib_18_s_axi_control_RRESP,
	fib_18_s_axi_control_AWREADY,
	fib_18_s_axi_control_AWVALID,
	fib_18_s_axi_control_AWADDR,
	fib_18_s_axi_control_WREADY,
	fib_18_s_axi_control_WVALID,
	fib_18_s_axi_control_WDATA,
	fib_18_s_axi_control_WSTRB,
	fib_18_s_axi_control_BREADY,
	fib_18_s_axi_control_BVALID,
	fib_18_s_axi_control_BRESP,
	fib_19_m_axi_gmem_ARREADY,
	fib_19_m_axi_gmem_ARVALID,
	fib_19_m_axi_gmem_ARID,
	fib_19_m_axi_gmem_ARADDR,
	fib_19_m_axi_gmem_ARLEN,
	fib_19_m_axi_gmem_ARSIZE,
	fib_19_m_axi_gmem_ARBURST,
	fib_19_m_axi_gmem_ARLOCK,
	fib_19_m_axi_gmem_ARCACHE,
	fib_19_m_axi_gmem_ARPROT,
	fib_19_m_axi_gmem_ARQOS,
	fib_19_m_axi_gmem_ARREGION,
	fib_19_m_axi_gmem_ARUSER,
	fib_19_m_axi_gmem_RREADY,
	fib_19_m_axi_gmem_RVALID,
	fib_19_m_axi_gmem_RID,
	fib_19_m_axi_gmem_RDATA,
	fib_19_m_axi_gmem_RRESP,
	fib_19_m_axi_gmem_RLAST,
	fib_19_m_axi_gmem_RUSER,
	fib_19_m_axi_gmem_AWREADY,
	fib_19_m_axi_gmem_AWVALID,
	fib_19_m_axi_gmem_AWID,
	fib_19_m_axi_gmem_AWADDR,
	fib_19_m_axi_gmem_AWLEN,
	fib_19_m_axi_gmem_AWSIZE,
	fib_19_m_axi_gmem_AWBURST,
	fib_19_m_axi_gmem_AWLOCK,
	fib_19_m_axi_gmem_AWCACHE,
	fib_19_m_axi_gmem_AWPROT,
	fib_19_m_axi_gmem_AWQOS,
	fib_19_m_axi_gmem_AWREGION,
	fib_19_m_axi_gmem_AWUSER,
	fib_19_m_axi_gmem_WREADY,
	fib_19_m_axi_gmem_WVALID,
	fib_19_m_axi_gmem_WDATA,
	fib_19_m_axi_gmem_WSTRB,
	fib_19_m_axi_gmem_WLAST,
	fib_19_m_axi_gmem_WUSER,
	fib_19_m_axi_gmem_BREADY,
	fib_19_m_axi_gmem_BVALID,
	fib_19_m_axi_gmem_BID,
	fib_19_m_axi_gmem_BRESP,
	fib_19_m_axi_gmem_BUSER,
	fib_19_s_axi_control_ARREADY,
	fib_19_s_axi_control_ARVALID,
	fib_19_s_axi_control_ARADDR,
	fib_19_s_axi_control_RREADY,
	fib_19_s_axi_control_RVALID,
	fib_19_s_axi_control_RDATA,
	fib_19_s_axi_control_RRESP,
	fib_19_s_axi_control_AWREADY,
	fib_19_s_axi_control_AWVALID,
	fib_19_s_axi_control_AWADDR,
	fib_19_s_axi_control_WREADY,
	fib_19_s_axi_control_WVALID,
	fib_19_s_axi_control_WDATA,
	fib_19_s_axi_control_WSTRB,
	fib_19_s_axi_control_BREADY,
	fib_19_s_axi_control_BVALID,
	fib_19_s_axi_control_BRESP,
	fib_20_m_axi_gmem_ARREADY,
	fib_20_m_axi_gmem_ARVALID,
	fib_20_m_axi_gmem_ARID,
	fib_20_m_axi_gmem_ARADDR,
	fib_20_m_axi_gmem_ARLEN,
	fib_20_m_axi_gmem_ARSIZE,
	fib_20_m_axi_gmem_ARBURST,
	fib_20_m_axi_gmem_ARLOCK,
	fib_20_m_axi_gmem_ARCACHE,
	fib_20_m_axi_gmem_ARPROT,
	fib_20_m_axi_gmem_ARQOS,
	fib_20_m_axi_gmem_ARREGION,
	fib_20_m_axi_gmem_ARUSER,
	fib_20_m_axi_gmem_RREADY,
	fib_20_m_axi_gmem_RVALID,
	fib_20_m_axi_gmem_RID,
	fib_20_m_axi_gmem_RDATA,
	fib_20_m_axi_gmem_RRESP,
	fib_20_m_axi_gmem_RLAST,
	fib_20_m_axi_gmem_RUSER,
	fib_20_m_axi_gmem_AWREADY,
	fib_20_m_axi_gmem_AWVALID,
	fib_20_m_axi_gmem_AWID,
	fib_20_m_axi_gmem_AWADDR,
	fib_20_m_axi_gmem_AWLEN,
	fib_20_m_axi_gmem_AWSIZE,
	fib_20_m_axi_gmem_AWBURST,
	fib_20_m_axi_gmem_AWLOCK,
	fib_20_m_axi_gmem_AWCACHE,
	fib_20_m_axi_gmem_AWPROT,
	fib_20_m_axi_gmem_AWQOS,
	fib_20_m_axi_gmem_AWREGION,
	fib_20_m_axi_gmem_AWUSER,
	fib_20_m_axi_gmem_WREADY,
	fib_20_m_axi_gmem_WVALID,
	fib_20_m_axi_gmem_WDATA,
	fib_20_m_axi_gmem_WSTRB,
	fib_20_m_axi_gmem_WLAST,
	fib_20_m_axi_gmem_WUSER,
	fib_20_m_axi_gmem_BREADY,
	fib_20_m_axi_gmem_BVALID,
	fib_20_m_axi_gmem_BID,
	fib_20_m_axi_gmem_BRESP,
	fib_20_m_axi_gmem_BUSER,
	fib_20_s_axi_control_ARREADY,
	fib_20_s_axi_control_ARVALID,
	fib_20_s_axi_control_ARADDR,
	fib_20_s_axi_control_RREADY,
	fib_20_s_axi_control_RVALID,
	fib_20_s_axi_control_RDATA,
	fib_20_s_axi_control_RRESP,
	fib_20_s_axi_control_AWREADY,
	fib_20_s_axi_control_AWVALID,
	fib_20_s_axi_control_AWADDR,
	fib_20_s_axi_control_WREADY,
	fib_20_s_axi_control_WVALID,
	fib_20_s_axi_control_WDATA,
	fib_20_s_axi_control_WSTRB,
	fib_20_s_axi_control_BREADY,
	fib_20_s_axi_control_BVALID,
	fib_20_s_axi_control_BRESP,
	fib_21_m_axi_gmem_ARREADY,
	fib_21_m_axi_gmem_ARVALID,
	fib_21_m_axi_gmem_ARID,
	fib_21_m_axi_gmem_ARADDR,
	fib_21_m_axi_gmem_ARLEN,
	fib_21_m_axi_gmem_ARSIZE,
	fib_21_m_axi_gmem_ARBURST,
	fib_21_m_axi_gmem_ARLOCK,
	fib_21_m_axi_gmem_ARCACHE,
	fib_21_m_axi_gmem_ARPROT,
	fib_21_m_axi_gmem_ARQOS,
	fib_21_m_axi_gmem_ARREGION,
	fib_21_m_axi_gmem_ARUSER,
	fib_21_m_axi_gmem_RREADY,
	fib_21_m_axi_gmem_RVALID,
	fib_21_m_axi_gmem_RID,
	fib_21_m_axi_gmem_RDATA,
	fib_21_m_axi_gmem_RRESP,
	fib_21_m_axi_gmem_RLAST,
	fib_21_m_axi_gmem_RUSER,
	fib_21_m_axi_gmem_AWREADY,
	fib_21_m_axi_gmem_AWVALID,
	fib_21_m_axi_gmem_AWID,
	fib_21_m_axi_gmem_AWADDR,
	fib_21_m_axi_gmem_AWLEN,
	fib_21_m_axi_gmem_AWSIZE,
	fib_21_m_axi_gmem_AWBURST,
	fib_21_m_axi_gmem_AWLOCK,
	fib_21_m_axi_gmem_AWCACHE,
	fib_21_m_axi_gmem_AWPROT,
	fib_21_m_axi_gmem_AWQOS,
	fib_21_m_axi_gmem_AWREGION,
	fib_21_m_axi_gmem_AWUSER,
	fib_21_m_axi_gmem_WREADY,
	fib_21_m_axi_gmem_WVALID,
	fib_21_m_axi_gmem_WDATA,
	fib_21_m_axi_gmem_WSTRB,
	fib_21_m_axi_gmem_WLAST,
	fib_21_m_axi_gmem_WUSER,
	fib_21_m_axi_gmem_BREADY,
	fib_21_m_axi_gmem_BVALID,
	fib_21_m_axi_gmem_BID,
	fib_21_m_axi_gmem_BRESP,
	fib_21_m_axi_gmem_BUSER,
	fib_21_s_axi_control_ARREADY,
	fib_21_s_axi_control_ARVALID,
	fib_21_s_axi_control_ARADDR,
	fib_21_s_axi_control_RREADY,
	fib_21_s_axi_control_RVALID,
	fib_21_s_axi_control_RDATA,
	fib_21_s_axi_control_RRESP,
	fib_21_s_axi_control_AWREADY,
	fib_21_s_axi_control_AWVALID,
	fib_21_s_axi_control_AWADDR,
	fib_21_s_axi_control_WREADY,
	fib_21_s_axi_control_WVALID,
	fib_21_s_axi_control_WDATA,
	fib_21_s_axi_control_WSTRB,
	fib_21_s_axi_control_BREADY,
	fib_21_s_axi_control_BVALID,
	fib_21_s_axi_control_BRESP,
	fib_22_m_axi_gmem_ARREADY,
	fib_22_m_axi_gmem_ARVALID,
	fib_22_m_axi_gmem_ARID,
	fib_22_m_axi_gmem_ARADDR,
	fib_22_m_axi_gmem_ARLEN,
	fib_22_m_axi_gmem_ARSIZE,
	fib_22_m_axi_gmem_ARBURST,
	fib_22_m_axi_gmem_ARLOCK,
	fib_22_m_axi_gmem_ARCACHE,
	fib_22_m_axi_gmem_ARPROT,
	fib_22_m_axi_gmem_ARQOS,
	fib_22_m_axi_gmem_ARREGION,
	fib_22_m_axi_gmem_ARUSER,
	fib_22_m_axi_gmem_RREADY,
	fib_22_m_axi_gmem_RVALID,
	fib_22_m_axi_gmem_RID,
	fib_22_m_axi_gmem_RDATA,
	fib_22_m_axi_gmem_RRESP,
	fib_22_m_axi_gmem_RLAST,
	fib_22_m_axi_gmem_RUSER,
	fib_22_m_axi_gmem_AWREADY,
	fib_22_m_axi_gmem_AWVALID,
	fib_22_m_axi_gmem_AWID,
	fib_22_m_axi_gmem_AWADDR,
	fib_22_m_axi_gmem_AWLEN,
	fib_22_m_axi_gmem_AWSIZE,
	fib_22_m_axi_gmem_AWBURST,
	fib_22_m_axi_gmem_AWLOCK,
	fib_22_m_axi_gmem_AWCACHE,
	fib_22_m_axi_gmem_AWPROT,
	fib_22_m_axi_gmem_AWQOS,
	fib_22_m_axi_gmem_AWREGION,
	fib_22_m_axi_gmem_AWUSER,
	fib_22_m_axi_gmem_WREADY,
	fib_22_m_axi_gmem_WVALID,
	fib_22_m_axi_gmem_WDATA,
	fib_22_m_axi_gmem_WSTRB,
	fib_22_m_axi_gmem_WLAST,
	fib_22_m_axi_gmem_WUSER,
	fib_22_m_axi_gmem_BREADY,
	fib_22_m_axi_gmem_BVALID,
	fib_22_m_axi_gmem_BID,
	fib_22_m_axi_gmem_BRESP,
	fib_22_m_axi_gmem_BUSER,
	fib_22_s_axi_control_ARREADY,
	fib_22_s_axi_control_ARVALID,
	fib_22_s_axi_control_ARADDR,
	fib_22_s_axi_control_RREADY,
	fib_22_s_axi_control_RVALID,
	fib_22_s_axi_control_RDATA,
	fib_22_s_axi_control_RRESP,
	fib_22_s_axi_control_AWREADY,
	fib_22_s_axi_control_AWVALID,
	fib_22_s_axi_control_AWADDR,
	fib_22_s_axi_control_WREADY,
	fib_22_s_axi_control_WVALID,
	fib_22_s_axi_control_WDATA,
	fib_22_s_axi_control_WSTRB,
	fib_22_s_axi_control_BREADY,
	fib_22_s_axi_control_BVALID,
	fib_22_s_axi_control_BRESP,
	fib_23_m_axi_gmem_ARREADY,
	fib_23_m_axi_gmem_ARVALID,
	fib_23_m_axi_gmem_ARID,
	fib_23_m_axi_gmem_ARADDR,
	fib_23_m_axi_gmem_ARLEN,
	fib_23_m_axi_gmem_ARSIZE,
	fib_23_m_axi_gmem_ARBURST,
	fib_23_m_axi_gmem_ARLOCK,
	fib_23_m_axi_gmem_ARCACHE,
	fib_23_m_axi_gmem_ARPROT,
	fib_23_m_axi_gmem_ARQOS,
	fib_23_m_axi_gmem_ARREGION,
	fib_23_m_axi_gmem_ARUSER,
	fib_23_m_axi_gmem_RREADY,
	fib_23_m_axi_gmem_RVALID,
	fib_23_m_axi_gmem_RID,
	fib_23_m_axi_gmem_RDATA,
	fib_23_m_axi_gmem_RRESP,
	fib_23_m_axi_gmem_RLAST,
	fib_23_m_axi_gmem_RUSER,
	fib_23_m_axi_gmem_AWREADY,
	fib_23_m_axi_gmem_AWVALID,
	fib_23_m_axi_gmem_AWID,
	fib_23_m_axi_gmem_AWADDR,
	fib_23_m_axi_gmem_AWLEN,
	fib_23_m_axi_gmem_AWSIZE,
	fib_23_m_axi_gmem_AWBURST,
	fib_23_m_axi_gmem_AWLOCK,
	fib_23_m_axi_gmem_AWCACHE,
	fib_23_m_axi_gmem_AWPROT,
	fib_23_m_axi_gmem_AWQOS,
	fib_23_m_axi_gmem_AWREGION,
	fib_23_m_axi_gmem_AWUSER,
	fib_23_m_axi_gmem_WREADY,
	fib_23_m_axi_gmem_WVALID,
	fib_23_m_axi_gmem_WDATA,
	fib_23_m_axi_gmem_WSTRB,
	fib_23_m_axi_gmem_WLAST,
	fib_23_m_axi_gmem_WUSER,
	fib_23_m_axi_gmem_BREADY,
	fib_23_m_axi_gmem_BVALID,
	fib_23_m_axi_gmem_BID,
	fib_23_m_axi_gmem_BRESP,
	fib_23_m_axi_gmem_BUSER,
	fib_23_s_axi_control_ARREADY,
	fib_23_s_axi_control_ARVALID,
	fib_23_s_axi_control_ARADDR,
	fib_23_s_axi_control_RREADY,
	fib_23_s_axi_control_RVALID,
	fib_23_s_axi_control_RDATA,
	fib_23_s_axi_control_RRESP,
	fib_23_s_axi_control_AWREADY,
	fib_23_s_axi_control_AWVALID,
	fib_23_s_axi_control_AWADDR,
	fib_23_s_axi_control_WREADY,
	fib_23_s_axi_control_WVALID,
	fib_23_s_axi_control_WDATA,
	fib_23_s_axi_control_WSTRB,
	fib_23_s_axi_control_BREADY,
	fib_23_s_axi_control_BVALID,
	fib_23_s_axi_control_BRESP,
	fib_24_m_axi_gmem_ARREADY,
	fib_24_m_axi_gmem_ARVALID,
	fib_24_m_axi_gmem_ARID,
	fib_24_m_axi_gmem_ARADDR,
	fib_24_m_axi_gmem_ARLEN,
	fib_24_m_axi_gmem_ARSIZE,
	fib_24_m_axi_gmem_ARBURST,
	fib_24_m_axi_gmem_ARLOCK,
	fib_24_m_axi_gmem_ARCACHE,
	fib_24_m_axi_gmem_ARPROT,
	fib_24_m_axi_gmem_ARQOS,
	fib_24_m_axi_gmem_ARREGION,
	fib_24_m_axi_gmem_ARUSER,
	fib_24_m_axi_gmem_RREADY,
	fib_24_m_axi_gmem_RVALID,
	fib_24_m_axi_gmem_RID,
	fib_24_m_axi_gmem_RDATA,
	fib_24_m_axi_gmem_RRESP,
	fib_24_m_axi_gmem_RLAST,
	fib_24_m_axi_gmem_RUSER,
	fib_24_m_axi_gmem_AWREADY,
	fib_24_m_axi_gmem_AWVALID,
	fib_24_m_axi_gmem_AWID,
	fib_24_m_axi_gmem_AWADDR,
	fib_24_m_axi_gmem_AWLEN,
	fib_24_m_axi_gmem_AWSIZE,
	fib_24_m_axi_gmem_AWBURST,
	fib_24_m_axi_gmem_AWLOCK,
	fib_24_m_axi_gmem_AWCACHE,
	fib_24_m_axi_gmem_AWPROT,
	fib_24_m_axi_gmem_AWQOS,
	fib_24_m_axi_gmem_AWREGION,
	fib_24_m_axi_gmem_AWUSER,
	fib_24_m_axi_gmem_WREADY,
	fib_24_m_axi_gmem_WVALID,
	fib_24_m_axi_gmem_WDATA,
	fib_24_m_axi_gmem_WSTRB,
	fib_24_m_axi_gmem_WLAST,
	fib_24_m_axi_gmem_WUSER,
	fib_24_m_axi_gmem_BREADY,
	fib_24_m_axi_gmem_BVALID,
	fib_24_m_axi_gmem_BID,
	fib_24_m_axi_gmem_BRESP,
	fib_24_m_axi_gmem_BUSER,
	fib_24_s_axi_control_ARREADY,
	fib_24_s_axi_control_ARVALID,
	fib_24_s_axi_control_ARADDR,
	fib_24_s_axi_control_RREADY,
	fib_24_s_axi_control_RVALID,
	fib_24_s_axi_control_RDATA,
	fib_24_s_axi_control_RRESP,
	fib_24_s_axi_control_AWREADY,
	fib_24_s_axi_control_AWVALID,
	fib_24_s_axi_control_AWADDR,
	fib_24_s_axi_control_WREADY,
	fib_24_s_axi_control_WVALID,
	fib_24_s_axi_control_WDATA,
	fib_24_s_axi_control_WSTRB,
	fib_24_s_axi_control_BREADY,
	fib_24_s_axi_control_BVALID,
	fib_24_s_axi_control_BRESP,
	fib_25_m_axi_gmem_ARREADY,
	fib_25_m_axi_gmem_ARVALID,
	fib_25_m_axi_gmem_ARID,
	fib_25_m_axi_gmem_ARADDR,
	fib_25_m_axi_gmem_ARLEN,
	fib_25_m_axi_gmem_ARSIZE,
	fib_25_m_axi_gmem_ARBURST,
	fib_25_m_axi_gmem_ARLOCK,
	fib_25_m_axi_gmem_ARCACHE,
	fib_25_m_axi_gmem_ARPROT,
	fib_25_m_axi_gmem_ARQOS,
	fib_25_m_axi_gmem_ARREGION,
	fib_25_m_axi_gmem_ARUSER,
	fib_25_m_axi_gmem_RREADY,
	fib_25_m_axi_gmem_RVALID,
	fib_25_m_axi_gmem_RID,
	fib_25_m_axi_gmem_RDATA,
	fib_25_m_axi_gmem_RRESP,
	fib_25_m_axi_gmem_RLAST,
	fib_25_m_axi_gmem_RUSER,
	fib_25_m_axi_gmem_AWREADY,
	fib_25_m_axi_gmem_AWVALID,
	fib_25_m_axi_gmem_AWID,
	fib_25_m_axi_gmem_AWADDR,
	fib_25_m_axi_gmem_AWLEN,
	fib_25_m_axi_gmem_AWSIZE,
	fib_25_m_axi_gmem_AWBURST,
	fib_25_m_axi_gmem_AWLOCK,
	fib_25_m_axi_gmem_AWCACHE,
	fib_25_m_axi_gmem_AWPROT,
	fib_25_m_axi_gmem_AWQOS,
	fib_25_m_axi_gmem_AWREGION,
	fib_25_m_axi_gmem_AWUSER,
	fib_25_m_axi_gmem_WREADY,
	fib_25_m_axi_gmem_WVALID,
	fib_25_m_axi_gmem_WDATA,
	fib_25_m_axi_gmem_WSTRB,
	fib_25_m_axi_gmem_WLAST,
	fib_25_m_axi_gmem_WUSER,
	fib_25_m_axi_gmem_BREADY,
	fib_25_m_axi_gmem_BVALID,
	fib_25_m_axi_gmem_BID,
	fib_25_m_axi_gmem_BRESP,
	fib_25_m_axi_gmem_BUSER,
	fib_25_s_axi_control_ARREADY,
	fib_25_s_axi_control_ARVALID,
	fib_25_s_axi_control_ARADDR,
	fib_25_s_axi_control_RREADY,
	fib_25_s_axi_control_RVALID,
	fib_25_s_axi_control_RDATA,
	fib_25_s_axi_control_RRESP,
	fib_25_s_axi_control_AWREADY,
	fib_25_s_axi_control_AWVALID,
	fib_25_s_axi_control_AWADDR,
	fib_25_s_axi_control_WREADY,
	fib_25_s_axi_control_WVALID,
	fib_25_s_axi_control_WDATA,
	fib_25_s_axi_control_WSTRB,
	fib_25_s_axi_control_BREADY,
	fib_25_s_axi_control_BVALID,
	fib_25_s_axi_control_BRESP,
	fib_26_m_axi_gmem_ARREADY,
	fib_26_m_axi_gmem_ARVALID,
	fib_26_m_axi_gmem_ARID,
	fib_26_m_axi_gmem_ARADDR,
	fib_26_m_axi_gmem_ARLEN,
	fib_26_m_axi_gmem_ARSIZE,
	fib_26_m_axi_gmem_ARBURST,
	fib_26_m_axi_gmem_ARLOCK,
	fib_26_m_axi_gmem_ARCACHE,
	fib_26_m_axi_gmem_ARPROT,
	fib_26_m_axi_gmem_ARQOS,
	fib_26_m_axi_gmem_ARREGION,
	fib_26_m_axi_gmem_ARUSER,
	fib_26_m_axi_gmem_RREADY,
	fib_26_m_axi_gmem_RVALID,
	fib_26_m_axi_gmem_RID,
	fib_26_m_axi_gmem_RDATA,
	fib_26_m_axi_gmem_RRESP,
	fib_26_m_axi_gmem_RLAST,
	fib_26_m_axi_gmem_RUSER,
	fib_26_m_axi_gmem_AWREADY,
	fib_26_m_axi_gmem_AWVALID,
	fib_26_m_axi_gmem_AWID,
	fib_26_m_axi_gmem_AWADDR,
	fib_26_m_axi_gmem_AWLEN,
	fib_26_m_axi_gmem_AWSIZE,
	fib_26_m_axi_gmem_AWBURST,
	fib_26_m_axi_gmem_AWLOCK,
	fib_26_m_axi_gmem_AWCACHE,
	fib_26_m_axi_gmem_AWPROT,
	fib_26_m_axi_gmem_AWQOS,
	fib_26_m_axi_gmem_AWREGION,
	fib_26_m_axi_gmem_AWUSER,
	fib_26_m_axi_gmem_WREADY,
	fib_26_m_axi_gmem_WVALID,
	fib_26_m_axi_gmem_WDATA,
	fib_26_m_axi_gmem_WSTRB,
	fib_26_m_axi_gmem_WLAST,
	fib_26_m_axi_gmem_WUSER,
	fib_26_m_axi_gmem_BREADY,
	fib_26_m_axi_gmem_BVALID,
	fib_26_m_axi_gmem_BID,
	fib_26_m_axi_gmem_BRESP,
	fib_26_m_axi_gmem_BUSER,
	fib_26_s_axi_control_ARREADY,
	fib_26_s_axi_control_ARVALID,
	fib_26_s_axi_control_ARADDR,
	fib_26_s_axi_control_RREADY,
	fib_26_s_axi_control_RVALID,
	fib_26_s_axi_control_RDATA,
	fib_26_s_axi_control_RRESP,
	fib_26_s_axi_control_AWREADY,
	fib_26_s_axi_control_AWVALID,
	fib_26_s_axi_control_AWADDR,
	fib_26_s_axi_control_WREADY,
	fib_26_s_axi_control_WVALID,
	fib_26_s_axi_control_WDATA,
	fib_26_s_axi_control_WSTRB,
	fib_26_s_axi_control_BREADY,
	fib_26_s_axi_control_BVALID,
	fib_26_s_axi_control_BRESP,
	fib_27_m_axi_gmem_ARREADY,
	fib_27_m_axi_gmem_ARVALID,
	fib_27_m_axi_gmem_ARID,
	fib_27_m_axi_gmem_ARADDR,
	fib_27_m_axi_gmem_ARLEN,
	fib_27_m_axi_gmem_ARSIZE,
	fib_27_m_axi_gmem_ARBURST,
	fib_27_m_axi_gmem_ARLOCK,
	fib_27_m_axi_gmem_ARCACHE,
	fib_27_m_axi_gmem_ARPROT,
	fib_27_m_axi_gmem_ARQOS,
	fib_27_m_axi_gmem_ARREGION,
	fib_27_m_axi_gmem_ARUSER,
	fib_27_m_axi_gmem_RREADY,
	fib_27_m_axi_gmem_RVALID,
	fib_27_m_axi_gmem_RID,
	fib_27_m_axi_gmem_RDATA,
	fib_27_m_axi_gmem_RRESP,
	fib_27_m_axi_gmem_RLAST,
	fib_27_m_axi_gmem_RUSER,
	fib_27_m_axi_gmem_AWREADY,
	fib_27_m_axi_gmem_AWVALID,
	fib_27_m_axi_gmem_AWID,
	fib_27_m_axi_gmem_AWADDR,
	fib_27_m_axi_gmem_AWLEN,
	fib_27_m_axi_gmem_AWSIZE,
	fib_27_m_axi_gmem_AWBURST,
	fib_27_m_axi_gmem_AWLOCK,
	fib_27_m_axi_gmem_AWCACHE,
	fib_27_m_axi_gmem_AWPROT,
	fib_27_m_axi_gmem_AWQOS,
	fib_27_m_axi_gmem_AWREGION,
	fib_27_m_axi_gmem_AWUSER,
	fib_27_m_axi_gmem_WREADY,
	fib_27_m_axi_gmem_WVALID,
	fib_27_m_axi_gmem_WDATA,
	fib_27_m_axi_gmem_WSTRB,
	fib_27_m_axi_gmem_WLAST,
	fib_27_m_axi_gmem_WUSER,
	fib_27_m_axi_gmem_BREADY,
	fib_27_m_axi_gmem_BVALID,
	fib_27_m_axi_gmem_BID,
	fib_27_m_axi_gmem_BRESP,
	fib_27_m_axi_gmem_BUSER,
	fib_27_s_axi_control_ARREADY,
	fib_27_s_axi_control_ARVALID,
	fib_27_s_axi_control_ARADDR,
	fib_27_s_axi_control_RREADY,
	fib_27_s_axi_control_RVALID,
	fib_27_s_axi_control_RDATA,
	fib_27_s_axi_control_RRESP,
	fib_27_s_axi_control_AWREADY,
	fib_27_s_axi_control_AWVALID,
	fib_27_s_axi_control_AWADDR,
	fib_27_s_axi_control_WREADY,
	fib_27_s_axi_control_WVALID,
	fib_27_s_axi_control_WDATA,
	fib_27_s_axi_control_WSTRB,
	fib_27_s_axi_control_BREADY,
	fib_27_s_axi_control_BVALID,
	fib_27_s_axi_control_BRESP,
	fib_28_m_axi_gmem_ARREADY,
	fib_28_m_axi_gmem_ARVALID,
	fib_28_m_axi_gmem_ARID,
	fib_28_m_axi_gmem_ARADDR,
	fib_28_m_axi_gmem_ARLEN,
	fib_28_m_axi_gmem_ARSIZE,
	fib_28_m_axi_gmem_ARBURST,
	fib_28_m_axi_gmem_ARLOCK,
	fib_28_m_axi_gmem_ARCACHE,
	fib_28_m_axi_gmem_ARPROT,
	fib_28_m_axi_gmem_ARQOS,
	fib_28_m_axi_gmem_ARREGION,
	fib_28_m_axi_gmem_ARUSER,
	fib_28_m_axi_gmem_RREADY,
	fib_28_m_axi_gmem_RVALID,
	fib_28_m_axi_gmem_RID,
	fib_28_m_axi_gmem_RDATA,
	fib_28_m_axi_gmem_RRESP,
	fib_28_m_axi_gmem_RLAST,
	fib_28_m_axi_gmem_RUSER,
	fib_28_m_axi_gmem_AWREADY,
	fib_28_m_axi_gmem_AWVALID,
	fib_28_m_axi_gmem_AWID,
	fib_28_m_axi_gmem_AWADDR,
	fib_28_m_axi_gmem_AWLEN,
	fib_28_m_axi_gmem_AWSIZE,
	fib_28_m_axi_gmem_AWBURST,
	fib_28_m_axi_gmem_AWLOCK,
	fib_28_m_axi_gmem_AWCACHE,
	fib_28_m_axi_gmem_AWPROT,
	fib_28_m_axi_gmem_AWQOS,
	fib_28_m_axi_gmem_AWREGION,
	fib_28_m_axi_gmem_AWUSER,
	fib_28_m_axi_gmem_WREADY,
	fib_28_m_axi_gmem_WVALID,
	fib_28_m_axi_gmem_WDATA,
	fib_28_m_axi_gmem_WSTRB,
	fib_28_m_axi_gmem_WLAST,
	fib_28_m_axi_gmem_WUSER,
	fib_28_m_axi_gmem_BREADY,
	fib_28_m_axi_gmem_BVALID,
	fib_28_m_axi_gmem_BID,
	fib_28_m_axi_gmem_BRESP,
	fib_28_m_axi_gmem_BUSER,
	fib_28_s_axi_control_ARREADY,
	fib_28_s_axi_control_ARVALID,
	fib_28_s_axi_control_ARADDR,
	fib_28_s_axi_control_RREADY,
	fib_28_s_axi_control_RVALID,
	fib_28_s_axi_control_RDATA,
	fib_28_s_axi_control_RRESP,
	fib_28_s_axi_control_AWREADY,
	fib_28_s_axi_control_AWVALID,
	fib_28_s_axi_control_AWADDR,
	fib_28_s_axi_control_WREADY,
	fib_28_s_axi_control_WVALID,
	fib_28_s_axi_control_WDATA,
	fib_28_s_axi_control_WSTRB,
	fib_28_s_axi_control_BREADY,
	fib_28_s_axi_control_BVALID,
	fib_28_s_axi_control_BRESP,
	fib_29_m_axi_gmem_ARREADY,
	fib_29_m_axi_gmem_ARVALID,
	fib_29_m_axi_gmem_ARID,
	fib_29_m_axi_gmem_ARADDR,
	fib_29_m_axi_gmem_ARLEN,
	fib_29_m_axi_gmem_ARSIZE,
	fib_29_m_axi_gmem_ARBURST,
	fib_29_m_axi_gmem_ARLOCK,
	fib_29_m_axi_gmem_ARCACHE,
	fib_29_m_axi_gmem_ARPROT,
	fib_29_m_axi_gmem_ARQOS,
	fib_29_m_axi_gmem_ARREGION,
	fib_29_m_axi_gmem_ARUSER,
	fib_29_m_axi_gmem_RREADY,
	fib_29_m_axi_gmem_RVALID,
	fib_29_m_axi_gmem_RID,
	fib_29_m_axi_gmem_RDATA,
	fib_29_m_axi_gmem_RRESP,
	fib_29_m_axi_gmem_RLAST,
	fib_29_m_axi_gmem_RUSER,
	fib_29_m_axi_gmem_AWREADY,
	fib_29_m_axi_gmem_AWVALID,
	fib_29_m_axi_gmem_AWID,
	fib_29_m_axi_gmem_AWADDR,
	fib_29_m_axi_gmem_AWLEN,
	fib_29_m_axi_gmem_AWSIZE,
	fib_29_m_axi_gmem_AWBURST,
	fib_29_m_axi_gmem_AWLOCK,
	fib_29_m_axi_gmem_AWCACHE,
	fib_29_m_axi_gmem_AWPROT,
	fib_29_m_axi_gmem_AWQOS,
	fib_29_m_axi_gmem_AWREGION,
	fib_29_m_axi_gmem_AWUSER,
	fib_29_m_axi_gmem_WREADY,
	fib_29_m_axi_gmem_WVALID,
	fib_29_m_axi_gmem_WDATA,
	fib_29_m_axi_gmem_WSTRB,
	fib_29_m_axi_gmem_WLAST,
	fib_29_m_axi_gmem_WUSER,
	fib_29_m_axi_gmem_BREADY,
	fib_29_m_axi_gmem_BVALID,
	fib_29_m_axi_gmem_BID,
	fib_29_m_axi_gmem_BRESP,
	fib_29_m_axi_gmem_BUSER,
	fib_29_s_axi_control_ARREADY,
	fib_29_s_axi_control_ARVALID,
	fib_29_s_axi_control_ARADDR,
	fib_29_s_axi_control_RREADY,
	fib_29_s_axi_control_RVALID,
	fib_29_s_axi_control_RDATA,
	fib_29_s_axi_control_RRESP,
	fib_29_s_axi_control_AWREADY,
	fib_29_s_axi_control_AWVALID,
	fib_29_s_axi_control_AWADDR,
	fib_29_s_axi_control_WREADY,
	fib_29_s_axi_control_WVALID,
	fib_29_s_axi_control_WDATA,
	fib_29_s_axi_control_WSTRB,
	fib_29_s_axi_control_BREADY,
	fib_29_s_axi_control_BVALID,
	fib_29_s_axi_control_BRESP,
	fib_30_m_axi_gmem_ARREADY,
	fib_30_m_axi_gmem_ARVALID,
	fib_30_m_axi_gmem_ARID,
	fib_30_m_axi_gmem_ARADDR,
	fib_30_m_axi_gmem_ARLEN,
	fib_30_m_axi_gmem_ARSIZE,
	fib_30_m_axi_gmem_ARBURST,
	fib_30_m_axi_gmem_ARLOCK,
	fib_30_m_axi_gmem_ARCACHE,
	fib_30_m_axi_gmem_ARPROT,
	fib_30_m_axi_gmem_ARQOS,
	fib_30_m_axi_gmem_ARREGION,
	fib_30_m_axi_gmem_ARUSER,
	fib_30_m_axi_gmem_RREADY,
	fib_30_m_axi_gmem_RVALID,
	fib_30_m_axi_gmem_RID,
	fib_30_m_axi_gmem_RDATA,
	fib_30_m_axi_gmem_RRESP,
	fib_30_m_axi_gmem_RLAST,
	fib_30_m_axi_gmem_RUSER,
	fib_30_m_axi_gmem_AWREADY,
	fib_30_m_axi_gmem_AWVALID,
	fib_30_m_axi_gmem_AWID,
	fib_30_m_axi_gmem_AWADDR,
	fib_30_m_axi_gmem_AWLEN,
	fib_30_m_axi_gmem_AWSIZE,
	fib_30_m_axi_gmem_AWBURST,
	fib_30_m_axi_gmem_AWLOCK,
	fib_30_m_axi_gmem_AWCACHE,
	fib_30_m_axi_gmem_AWPROT,
	fib_30_m_axi_gmem_AWQOS,
	fib_30_m_axi_gmem_AWREGION,
	fib_30_m_axi_gmem_AWUSER,
	fib_30_m_axi_gmem_WREADY,
	fib_30_m_axi_gmem_WVALID,
	fib_30_m_axi_gmem_WDATA,
	fib_30_m_axi_gmem_WSTRB,
	fib_30_m_axi_gmem_WLAST,
	fib_30_m_axi_gmem_WUSER,
	fib_30_m_axi_gmem_BREADY,
	fib_30_m_axi_gmem_BVALID,
	fib_30_m_axi_gmem_BID,
	fib_30_m_axi_gmem_BRESP,
	fib_30_m_axi_gmem_BUSER,
	fib_30_s_axi_control_ARREADY,
	fib_30_s_axi_control_ARVALID,
	fib_30_s_axi_control_ARADDR,
	fib_30_s_axi_control_RREADY,
	fib_30_s_axi_control_RVALID,
	fib_30_s_axi_control_RDATA,
	fib_30_s_axi_control_RRESP,
	fib_30_s_axi_control_AWREADY,
	fib_30_s_axi_control_AWVALID,
	fib_30_s_axi_control_AWADDR,
	fib_30_s_axi_control_WREADY,
	fib_30_s_axi_control_WVALID,
	fib_30_s_axi_control_WDATA,
	fib_30_s_axi_control_WSTRB,
	fib_30_s_axi_control_BREADY,
	fib_30_s_axi_control_BVALID,
	fib_30_s_axi_control_BRESP,
	fib_31_m_axi_gmem_ARREADY,
	fib_31_m_axi_gmem_ARVALID,
	fib_31_m_axi_gmem_ARID,
	fib_31_m_axi_gmem_ARADDR,
	fib_31_m_axi_gmem_ARLEN,
	fib_31_m_axi_gmem_ARSIZE,
	fib_31_m_axi_gmem_ARBURST,
	fib_31_m_axi_gmem_ARLOCK,
	fib_31_m_axi_gmem_ARCACHE,
	fib_31_m_axi_gmem_ARPROT,
	fib_31_m_axi_gmem_ARQOS,
	fib_31_m_axi_gmem_ARREGION,
	fib_31_m_axi_gmem_ARUSER,
	fib_31_m_axi_gmem_RREADY,
	fib_31_m_axi_gmem_RVALID,
	fib_31_m_axi_gmem_RID,
	fib_31_m_axi_gmem_RDATA,
	fib_31_m_axi_gmem_RRESP,
	fib_31_m_axi_gmem_RLAST,
	fib_31_m_axi_gmem_RUSER,
	fib_31_m_axi_gmem_AWREADY,
	fib_31_m_axi_gmem_AWVALID,
	fib_31_m_axi_gmem_AWID,
	fib_31_m_axi_gmem_AWADDR,
	fib_31_m_axi_gmem_AWLEN,
	fib_31_m_axi_gmem_AWSIZE,
	fib_31_m_axi_gmem_AWBURST,
	fib_31_m_axi_gmem_AWLOCK,
	fib_31_m_axi_gmem_AWCACHE,
	fib_31_m_axi_gmem_AWPROT,
	fib_31_m_axi_gmem_AWQOS,
	fib_31_m_axi_gmem_AWREGION,
	fib_31_m_axi_gmem_AWUSER,
	fib_31_m_axi_gmem_WREADY,
	fib_31_m_axi_gmem_WVALID,
	fib_31_m_axi_gmem_WDATA,
	fib_31_m_axi_gmem_WSTRB,
	fib_31_m_axi_gmem_WLAST,
	fib_31_m_axi_gmem_WUSER,
	fib_31_m_axi_gmem_BREADY,
	fib_31_m_axi_gmem_BVALID,
	fib_31_m_axi_gmem_BID,
	fib_31_m_axi_gmem_BRESP,
	fib_31_m_axi_gmem_BUSER,
	fib_31_s_axi_control_ARREADY,
	fib_31_s_axi_control_ARVALID,
	fib_31_s_axi_control_ARADDR,
	fib_31_s_axi_control_RREADY,
	fib_31_s_axi_control_RVALID,
	fib_31_s_axi_control_RDATA,
	fib_31_s_axi_control_RRESP,
	fib_31_s_axi_control_AWREADY,
	fib_31_s_axi_control_AWVALID,
	fib_31_s_axi_control_AWADDR,
	fib_31_s_axi_control_WREADY,
	fib_31_s_axi_control_WVALID,
	fib_31_s_axi_control_WDATA,
	fib_31_s_axi_control_WSTRB,
	fib_31_s_axi_control_BREADY,
	fib_31_s_axi_control_BVALID,
	fib_31_s_axi_control_BRESP,
	fib_32_m_axi_gmem_ARREADY,
	fib_32_m_axi_gmem_ARVALID,
	fib_32_m_axi_gmem_ARID,
	fib_32_m_axi_gmem_ARADDR,
	fib_32_m_axi_gmem_ARLEN,
	fib_32_m_axi_gmem_ARSIZE,
	fib_32_m_axi_gmem_ARBURST,
	fib_32_m_axi_gmem_ARLOCK,
	fib_32_m_axi_gmem_ARCACHE,
	fib_32_m_axi_gmem_ARPROT,
	fib_32_m_axi_gmem_ARQOS,
	fib_32_m_axi_gmem_ARREGION,
	fib_32_m_axi_gmem_ARUSER,
	fib_32_m_axi_gmem_RREADY,
	fib_32_m_axi_gmem_RVALID,
	fib_32_m_axi_gmem_RID,
	fib_32_m_axi_gmem_RDATA,
	fib_32_m_axi_gmem_RRESP,
	fib_32_m_axi_gmem_RLAST,
	fib_32_m_axi_gmem_RUSER,
	fib_32_m_axi_gmem_AWREADY,
	fib_32_m_axi_gmem_AWVALID,
	fib_32_m_axi_gmem_AWID,
	fib_32_m_axi_gmem_AWADDR,
	fib_32_m_axi_gmem_AWLEN,
	fib_32_m_axi_gmem_AWSIZE,
	fib_32_m_axi_gmem_AWBURST,
	fib_32_m_axi_gmem_AWLOCK,
	fib_32_m_axi_gmem_AWCACHE,
	fib_32_m_axi_gmem_AWPROT,
	fib_32_m_axi_gmem_AWQOS,
	fib_32_m_axi_gmem_AWREGION,
	fib_32_m_axi_gmem_AWUSER,
	fib_32_m_axi_gmem_WREADY,
	fib_32_m_axi_gmem_WVALID,
	fib_32_m_axi_gmem_WDATA,
	fib_32_m_axi_gmem_WSTRB,
	fib_32_m_axi_gmem_WLAST,
	fib_32_m_axi_gmem_WUSER,
	fib_32_m_axi_gmem_BREADY,
	fib_32_m_axi_gmem_BVALID,
	fib_32_m_axi_gmem_BID,
	fib_32_m_axi_gmem_BRESP,
	fib_32_m_axi_gmem_BUSER,
	fib_32_s_axi_control_ARREADY,
	fib_32_s_axi_control_ARVALID,
	fib_32_s_axi_control_ARADDR,
	fib_32_s_axi_control_RREADY,
	fib_32_s_axi_control_RVALID,
	fib_32_s_axi_control_RDATA,
	fib_32_s_axi_control_RRESP,
	fib_32_s_axi_control_AWREADY,
	fib_32_s_axi_control_AWVALID,
	fib_32_s_axi_control_AWADDR,
	fib_32_s_axi_control_WREADY,
	fib_32_s_axi_control_WVALID,
	fib_32_s_axi_control_WDATA,
	fib_32_s_axi_control_WSTRB,
	fib_32_s_axi_control_BREADY,
	fib_32_s_axi_control_BVALID,
	fib_32_s_axi_control_BRESP,
	fib_33_m_axi_gmem_ARREADY,
	fib_33_m_axi_gmem_ARVALID,
	fib_33_m_axi_gmem_ARID,
	fib_33_m_axi_gmem_ARADDR,
	fib_33_m_axi_gmem_ARLEN,
	fib_33_m_axi_gmem_ARSIZE,
	fib_33_m_axi_gmem_ARBURST,
	fib_33_m_axi_gmem_ARLOCK,
	fib_33_m_axi_gmem_ARCACHE,
	fib_33_m_axi_gmem_ARPROT,
	fib_33_m_axi_gmem_ARQOS,
	fib_33_m_axi_gmem_ARREGION,
	fib_33_m_axi_gmem_ARUSER,
	fib_33_m_axi_gmem_RREADY,
	fib_33_m_axi_gmem_RVALID,
	fib_33_m_axi_gmem_RID,
	fib_33_m_axi_gmem_RDATA,
	fib_33_m_axi_gmem_RRESP,
	fib_33_m_axi_gmem_RLAST,
	fib_33_m_axi_gmem_RUSER,
	fib_33_m_axi_gmem_AWREADY,
	fib_33_m_axi_gmem_AWVALID,
	fib_33_m_axi_gmem_AWID,
	fib_33_m_axi_gmem_AWADDR,
	fib_33_m_axi_gmem_AWLEN,
	fib_33_m_axi_gmem_AWSIZE,
	fib_33_m_axi_gmem_AWBURST,
	fib_33_m_axi_gmem_AWLOCK,
	fib_33_m_axi_gmem_AWCACHE,
	fib_33_m_axi_gmem_AWPROT,
	fib_33_m_axi_gmem_AWQOS,
	fib_33_m_axi_gmem_AWREGION,
	fib_33_m_axi_gmem_AWUSER,
	fib_33_m_axi_gmem_WREADY,
	fib_33_m_axi_gmem_WVALID,
	fib_33_m_axi_gmem_WDATA,
	fib_33_m_axi_gmem_WSTRB,
	fib_33_m_axi_gmem_WLAST,
	fib_33_m_axi_gmem_WUSER,
	fib_33_m_axi_gmem_BREADY,
	fib_33_m_axi_gmem_BVALID,
	fib_33_m_axi_gmem_BID,
	fib_33_m_axi_gmem_BRESP,
	fib_33_m_axi_gmem_BUSER,
	fib_33_s_axi_control_ARREADY,
	fib_33_s_axi_control_ARVALID,
	fib_33_s_axi_control_ARADDR,
	fib_33_s_axi_control_RREADY,
	fib_33_s_axi_control_RVALID,
	fib_33_s_axi_control_RDATA,
	fib_33_s_axi_control_RRESP,
	fib_33_s_axi_control_AWREADY,
	fib_33_s_axi_control_AWVALID,
	fib_33_s_axi_control_AWADDR,
	fib_33_s_axi_control_WREADY,
	fib_33_s_axi_control_WVALID,
	fib_33_s_axi_control_WDATA,
	fib_33_s_axi_control_WSTRB,
	fib_33_s_axi_control_BREADY,
	fib_33_s_axi_control_BVALID,
	fib_33_s_axi_control_BRESP,
	fib_34_m_axi_gmem_ARREADY,
	fib_34_m_axi_gmem_ARVALID,
	fib_34_m_axi_gmem_ARID,
	fib_34_m_axi_gmem_ARADDR,
	fib_34_m_axi_gmem_ARLEN,
	fib_34_m_axi_gmem_ARSIZE,
	fib_34_m_axi_gmem_ARBURST,
	fib_34_m_axi_gmem_ARLOCK,
	fib_34_m_axi_gmem_ARCACHE,
	fib_34_m_axi_gmem_ARPROT,
	fib_34_m_axi_gmem_ARQOS,
	fib_34_m_axi_gmem_ARREGION,
	fib_34_m_axi_gmem_ARUSER,
	fib_34_m_axi_gmem_RREADY,
	fib_34_m_axi_gmem_RVALID,
	fib_34_m_axi_gmem_RID,
	fib_34_m_axi_gmem_RDATA,
	fib_34_m_axi_gmem_RRESP,
	fib_34_m_axi_gmem_RLAST,
	fib_34_m_axi_gmem_RUSER,
	fib_34_m_axi_gmem_AWREADY,
	fib_34_m_axi_gmem_AWVALID,
	fib_34_m_axi_gmem_AWID,
	fib_34_m_axi_gmem_AWADDR,
	fib_34_m_axi_gmem_AWLEN,
	fib_34_m_axi_gmem_AWSIZE,
	fib_34_m_axi_gmem_AWBURST,
	fib_34_m_axi_gmem_AWLOCK,
	fib_34_m_axi_gmem_AWCACHE,
	fib_34_m_axi_gmem_AWPROT,
	fib_34_m_axi_gmem_AWQOS,
	fib_34_m_axi_gmem_AWREGION,
	fib_34_m_axi_gmem_AWUSER,
	fib_34_m_axi_gmem_WREADY,
	fib_34_m_axi_gmem_WVALID,
	fib_34_m_axi_gmem_WDATA,
	fib_34_m_axi_gmem_WSTRB,
	fib_34_m_axi_gmem_WLAST,
	fib_34_m_axi_gmem_WUSER,
	fib_34_m_axi_gmem_BREADY,
	fib_34_m_axi_gmem_BVALID,
	fib_34_m_axi_gmem_BID,
	fib_34_m_axi_gmem_BRESP,
	fib_34_m_axi_gmem_BUSER,
	fib_34_s_axi_control_ARREADY,
	fib_34_s_axi_control_ARVALID,
	fib_34_s_axi_control_ARADDR,
	fib_34_s_axi_control_RREADY,
	fib_34_s_axi_control_RVALID,
	fib_34_s_axi_control_RDATA,
	fib_34_s_axi_control_RRESP,
	fib_34_s_axi_control_AWREADY,
	fib_34_s_axi_control_AWVALID,
	fib_34_s_axi_control_AWADDR,
	fib_34_s_axi_control_WREADY,
	fib_34_s_axi_control_WVALID,
	fib_34_s_axi_control_WDATA,
	fib_34_s_axi_control_WSTRB,
	fib_34_s_axi_control_BREADY,
	fib_34_s_axi_control_BVALID,
	fib_34_s_axi_control_BRESP,
	fib_35_m_axi_gmem_ARREADY,
	fib_35_m_axi_gmem_ARVALID,
	fib_35_m_axi_gmem_ARID,
	fib_35_m_axi_gmem_ARADDR,
	fib_35_m_axi_gmem_ARLEN,
	fib_35_m_axi_gmem_ARSIZE,
	fib_35_m_axi_gmem_ARBURST,
	fib_35_m_axi_gmem_ARLOCK,
	fib_35_m_axi_gmem_ARCACHE,
	fib_35_m_axi_gmem_ARPROT,
	fib_35_m_axi_gmem_ARQOS,
	fib_35_m_axi_gmem_ARREGION,
	fib_35_m_axi_gmem_ARUSER,
	fib_35_m_axi_gmem_RREADY,
	fib_35_m_axi_gmem_RVALID,
	fib_35_m_axi_gmem_RID,
	fib_35_m_axi_gmem_RDATA,
	fib_35_m_axi_gmem_RRESP,
	fib_35_m_axi_gmem_RLAST,
	fib_35_m_axi_gmem_RUSER,
	fib_35_m_axi_gmem_AWREADY,
	fib_35_m_axi_gmem_AWVALID,
	fib_35_m_axi_gmem_AWID,
	fib_35_m_axi_gmem_AWADDR,
	fib_35_m_axi_gmem_AWLEN,
	fib_35_m_axi_gmem_AWSIZE,
	fib_35_m_axi_gmem_AWBURST,
	fib_35_m_axi_gmem_AWLOCK,
	fib_35_m_axi_gmem_AWCACHE,
	fib_35_m_axi_gmem_AWPROT,
	fib_35_m_axi_gmem_AWQOS,
	fib_35_m_axi_gmem_AWREGION,
	fib_35_m_axi_gmem_AWUSER,
	fib_35_m_axi_gmem_WREADY,
	fib_35_m_axi_gmem_WVALID,
	fib_35_m_axi_gmem_WDATA,
	fib_35_m_axi_gmem_WSTRB,
	fib_35_m_axi_gmem_WLAST,
	fib_35_m_axi_gmem_WUSER,
	fib_35_m_axi_gmem_BREADY,
	fib_35_m_axi_gmem_BVALID,
	fib_35_m_axi_gmem_BID,
	fib_35_m_axi_gmem_BRESP,
	fib_35_m_axi_gmem_BUSER,
	fib_35_s_axi_control_ARREADY,
	fib_35_s_axi_control_ARVALID,
	fib_35_s_axi_control_ARADDR,
	fib_35_s_axi_control_RREADY,
	fib_35_s_axi_control_RVALID,
	fib_35_s_axi_control_RDATA,
	fib_35_s_axi_control_RRESP,
	fib_35_s_axi_control_AWREADY,
	fib_35_s_axi_control_AWVALID,
	fib_35_s_axi_control_AWADDR,
	fib_35_s_axi_control_WREADY,
	fib_35_s_axi_control_WVALID,
	fib_35_s_axi_control_WDATA,
	fib_35_s_axi_control_WSTRB,
	fib_35_s_axi_control_BREADY,
	fib_35_s_axi_control_BVALID,
	fib_35_s_axi_control_BRESP,
	fib_36_m_axi_gmem_ARREADY,
	fib_36_m_axi_gmem_ARVALID,
	fib_36_m_axi_gmem_ARID,
	fib_36_m_axi_gmem_ARADDR,
	fib_36_m_axi_gmem_ARLEN,
	fib_36_m_axi_gmem_ARSIZE,
	fib_36_m_axi_gmem_ARBURST,
	fib_36_m_axi_gmem_ARLOCK,
	fib_36_m_axi_gmem_ARCACHE,
	fib_36_m_axi_gmem_ARPROT,
	fib_36_m_axi_gmem_ARQOS,
	fib_36_m_axi_gmem_ARREGION,
	fib_36_m_axi_gmem_ARUSER,
	fib_36_m_axi_gmem_RREADY,
	fib_36_m_axi_gmem_RVALID,
	fib_36_m_axi_gmem_RID,
	fib_36_m_axi_gmem_RDATA,
	fib_36_m_axi_gmem_RRESP,
	fib_36_m_axi_gmem_RLAST,
	fib_36_m_axi_gmem_RUSER,
	fib_36_m_axi_gmem_AWREADY,
	fib_36_m_axi_gmem_AWVALID,
	fib_36_m_axi_gmem_AWID,
	fib_36_m_axi_gmem_AWADDR,
	fib_36_m_axi_gmem_AWLEN,
	fib_36_m_axi_gmem_AWSIZE,
	fib_36_m_axi_gmem_AWBURST,
	fib_36_m_axi_gmem_AWLOCK,
	fib_36_m_axi_gmem_AWCACHE,
	fib_36_m_axi_gmem_AWPROT,
	fib_36_m_axi_gmem_AWQOS,
	fib_36_m_axi_gmem_AWREGION,
	fib_36_m_axi_gmem_AWUSER,
	fib_36_m_axi_gmem_WREADY,
	fib_36_m_axi_gmem_WVALID,
	fib_36_m_axi_gmem_WDATA,
	fib_36_m_axi_gmem_WSTRB,
	fib_36_m_axi_gmem_WLAST,
	fib_36_m_axi_gmem_WUSER,
	fib_36_m_axi_gmem_BREADY,
	fib_36_m_axi_gmem_BVALID,
	fib_36_m_axi_gmem_BID,
	fib_36_m_axi_gmem_BRESP,
	fib_36_m_axi_gmem_BUSER,
	fib_36_s_axi_control_ARREADY,
	fib_36_s_axi_control_ARVALID,
	fib_36_s_axi_control_ARADDR,
	fib_36_s_axi_control_RREADY,
	fib_36_s_axi_control_RVALID,
	fib_36_s_axi_control_RDATA,
	fib_36_s_axi_control_RRESP,
	fib_36_s_axi_control_AWREADY,
	fib_36_s_axi_control_AWVALID,
	fib_36_s_axi_control_AWADDR,
	fib_36_s_axi_control_WREADY,
	fib_36_s_axi_control_WVALID,
	fib_36_s_axi_control_WDATA,
	fib_36_s_axi_control_WSTRB,
	fib_36_s_axi_control_BREADY,
	fib_36_s_axi_control_BVALID,
	fib_36_s_axi_control_BRESP,
	fib_37_m_axi_gmem_ARREADY,
	fib_37_m_axi_gmem_ARVALID,
	fib_37_m_axi_gmem_ARID,
	fib_37_m_axi_gmem_ARADDR,
	fib_37_m_axi_gmem_ARLEN,
	fib_37_m_axi_gmem_ARSIZE,
	fib_37_m_axi_gmem_ARBURST,
	fib_37_m_axi_gmem_ARLOCK,
	fib_37_m_axi_gmem_ARCACHE,
	fib_37_m_axi_gmem_ARPROT,
	fib_37_m_axi_gmem_ARQOS,
	fib_37_m_axi_gmem_ARREGION,
	fib_37_m_axi_gmem_ARUSER,
	fib_37_m_axi_gmem_RREADY,
	fib_37_m_axi_gmem_RVALID,
	fib_37_m_axi_gmem_RID,
	fib_37_m_axi_gmem_RDATA,
	fib_37_m_axi_gmem_RRESP,
	fib_37_m_axi_gmem_RLAST,
	fib_37_m_axi_gmem_RUSER,
	fib_37_m_axi_gmem_AWREADY,
	fib_37_m_axi_gmem_AWVALID,
	fib_37_m_axi_gmem_AWID,
	fib_37_m_axi_gmem_AWADDR,
	fib_37_m_axi_gmem_AWLEN,
	fib_37_m_axi_gmem_AWSIZE,
	fib_37_m_axi_gmem_AWBURST,
	fib_37_m_axi_gmem_AWLOCK,
	fib_37_m_axi_gmem_AWCACHE,
	fib_37_m_axi_gmem_AWPROT,
	fib_37_m_axi_gmem_AWQOS,
	fib_37_m_axi_gmem_AWREGION,
	fib_37_m_axi_gmem_AWUSER,
	fib_37_m_axi_gmem_WREADY,
	fib_37_m_axi_gmem_WVALID,
	fib_37_m_axi_gmem_WDATA,
	fib_37_m_axi_gmem_WSTRB,
	fib_37_m_axi_gmem_WLAST,
	fib_37_m_axi_gmem_WUSER,
	fib_37_m_axi_gmem_BREADY,
	fib_37_m_axi_gmem_BVALID,
	fib_37_m_axi_gmem_BID,
	fib_37_m_axi_gmem_BRESP,
	fib_37_m_axi_gmem_BUSER,
	fib_37_s_axi_control_ARREADY,
	fib_37_s_axi_control_ARVALID,
	fib_37_s_axi_control_ARADDR,
	fib_37_s_axi_control_RREADY,
	fib_37_s_axi_control_RVALID,
	fib_37_s_axi_control_RDATA,
	fib_37_s_axi_control_RRESP,
	fib_37_s_axi_control_AWREADY,
	fib_37_s_axi_control_AWVALID,
	fib_37_s_axi_control_AWADDR,
	fib_37_s_axi_control_WREADY,
	fib_37_s_axi_control_WVALID,
	fib_37_s_axi_control_WDATA,
	fib_37_s_axi_control_WSTRB,
	fib_37_s_axi_control_BREADY,
	fib_37_s_axi_control_BVALID,
	fib_37_s_axi_control_BRESP,
	fib_38_m_axi_gmem_ARREADY,
	fib_38_m_axi_gmem_ARVALID,
	fib_38_m_axi_gmem_ARID,
	fib_38_m_axi_gmem_ARADDR,
	fib_38_m_axi_gmem_ARLEN,
	fib_38_m_axi_gmem_ARSIZE,
	fib_38_m_axi_gmem_ARBURST,
	fib_38_m_axi_gmem_ARLOCK,
	fib_38_m_axi_gmem_ARCACHE,
	fib_38_m_axi_gmem_ARPROT,
	fib_38_m_axi_gmem_ARQOS,
	fib_38_m_axi_gmem_ARREGION,
	fib_38_m_axi_gmem_ARUSER,
	fib_38_m_axi_gmem_RREADY,
	fib_38_m_axi_gmem_RVALID,
	fib_38_m_axi_gmem_RID,
	fib_38_m_axi_gmem_RDATA,
	fib_38_m_axi_gmem_RRESP,
	fib_38_m_axi_gmem_RLAST,
	fib_38_m_axi_gmem_RUSER,
	fib_38_m_axi_gmem_AWREADY,
	fib_38_m_axi_gmem_AWVALID,
	fib_38_m_axi_gmem_AWID,
	fib_38_m_axi_gmem_AWADDR,
	fib_38_m_axi_gmem_AWLEN,
	fib_38_m_axi_gmem_AWSIZE,
	fib_38_m_axi_gmem_AWBURST,
	fib_38_m_axi_gmem_AWLOCK,
	fib_38_m_axi_gmem_AWCACHE,
	fib_38_m_axi_gmem_AWPROT,
	fib_38_m_axi_gmem_AWQOS,
	fib_38_m_axi_gmem_AWREGION,
	fib_38_m_axi_gmem_AWUSER,
	fib_38_m_axi_gmem_WREADY,
	fib_38_m_axi_gmem_WVALID,
	fib_38_m_axi_gmem_WDATA,
	fib_38_m_axi_gmem_WSTRB,
	fib_38_m_axi_gmem_WLAST,
	fib_38_m_axi_gmem_WUSER,
	fib_38_m_axi_gmem_BREADY,
	fib_38_m_axi_gmem_BVALID,
	fib_38_m_axi_gmem_BID,
	fib_38_m_axi_gmem_BRESP,
	fib_38_m_axi_gmem_BUSER,
	fib_38_s_axi_control_ARREADY,
	fib_38_s_axi_control_ARVALID,
	fib_38_s_axi_control_ARADDR,
	fib_38_s_axi_control_RREADY,
	fib_38_s_axi_control_RVALID,
	fib_38_s_axi_control_RDATA,
	fib_38_s_axi_control_RRESP,
	fib_38_s_axi_control_AWREADY,
	fib_38_s_axi_control_AWVALID,
	fib_38_s_axi_control_AWADDR,
	fib_38_s_axi_control_WREADY,
	fib_38_s_axi_control_WVALID,
	fib_38_s_axi_control_WDATA,
	fib_38_s_axi_control_WSTRB,
	fib_38_s_axi_control_BREADY,
	fib_38_s_axi_control_BVALID,
	fib_38_s_axi_control_BRESP,
	fib_39_m_axi_gmem_ARREADY,
	fib_39_m_axi_gmem_ARVALID,
	fib_39_m_axi_gmem_ARID,
	fib_39_m_axi_gmem_ARADDR,
	fib_39_m_axi_gmem_ARLEN,
	fib_39_m_axi_gmem_ARSIZE,
	fib_39_m_axi_gmem_ARBURST,
	fib_39_m_axi_gmem_ARLOCK,
	fib_39_m_axi_gmem_ARCACHE,
	fib_39_m_axi_gmem_ARPROT,
	fib_39_m_axi_gmem_ARQOS,
	fib_39_m_axi_gmem_ARREGION,
	fib_39_m_axi_gmem_ARUSER,
	fib_39_m_axi_gmem_RREADY,
	fib_39_m_axi_gmem_RVALID,
	fib_39_m_axi_gmem_RID,
	fib_39_m_axi_gmem_RDATA,
	fib_39_m_axi_gmem_RRESP,
	fib_39_m_axi_gmem_RLAST,
	fib_39_m_axi_gmem_RUSER,
	fib_39_m_axi_gmem_AWREADY,
	fib_39_m_axi_gmem_AWVALID,
	fib_39_m_axi_gmem_AWID,
	fib_39_m_axi_gmem_AWADDR,
	fib_39_m_axi_gmem_AWLEN,
	fib_39_m_axi_gmem_AWSIZE,
	fib_39_m_axi_gmem_AWBURST,
	fib_39_m_axi_gmem_AWLOCK,
	fib_39_m_axi_gmem_AWCACHE,
	fib_39_m_axi_gmem_AWPROT,
	fib_39_m_axi_gmem_AWQOS,
	fib_39_m_axi_gmem_AWREGION,
	fib_39_m_axi_gmem_AWUSER,
	fib_39_m_axi_gmem_WREADY,
	fib_39_m_axi_gmem_WVALID,
	fib_39_m_axi_gmem_WDATA,
	fib_39_m_axi_gmem_WSTRB,
	fib_39_m_axi_gmem_WLAST,
	fib_39_m_axi_gmem_WUSER,
	fib_39_m_axi_gmem_BREADY,
	fib_39_m_axi_gmem_BVALID,
	fib_39_m_axi_gmem_BID,
	fib_39_m_axi_gmem_BRESP,
	fib_39_m_axi_gmem_BUSER,
	fib_39_s_axi_control_ARREADY,
	fib_39_s_axi_control_ARVALID,
	fib_39_s_axi_control_ARADDR,
	fib_39_s_axi_control_RREADY,
	fib_39_s_axi_control_RVALID,
	fib_39_s_axi_control_RDATA,
	fib_39_s_axi_control_RRESP,
	fib_39_s_axi_control_AWREADY,
	fib_39_s_axi_control_AWVALID,
	fib_39_s_axi_control_AWADDR,
	fib_39_s_axi_control_WREADY,
	fib_39_s_axi_control_WVALID,
	fib_39_s_axi_control_WDATA,
	fib_39_s_axi_control_WSTRB,
	fib_39_s_axi_control_BREADY,
	fib_39_s_axi_control_BVALID,
	fib_39_s_axi_control_BRESP,
	fib_40_m_axi_gmem_ARREADY,
	fib_40_m_axi_gmem_ARVALID,
	fib_40_m_axi_gmem_ARID,
	fib_40_m_axi_gmem_ARADDR,
	fib_40_m_axi_gmem_ARLEN,
	fib_40_m_axi_gmem_ARSIZE,
	fib_40_m_axi_gmem_ARBURST,
	fib_40_m_axi_gmem_ARLOCK,
	fib_40_m_axi_gmem_ARCACHE,
	fib_40_m_axi_gmem_ARPROT,
	fib_40_m_axi_gmem_ARQOS,
	fib_40_m_axi_gmem_ARREGION,
	fib_40_m_axi_gmem_ARUSER,
	fib_40_m_axi_gmem_RREADY,
	fib_40_m_axi_gmem_RVALID,
	fib_40_m_axi_gmem_RID,
	fib_40_m_axi_gmem_RDATA,
	fib_40_m_axi_gmem_RRESP,
	fib_40_m_axi_gmem_RLAST,
	fib_40_m_axi_gmem_RUSER,
	fib_40_m_axi_gmem_AWREADY,
	fib_40_m_axi_gmem_AWVALID,
	fib_40_m_axi_gmem_AWID,
	fib_40_m_axi_gmem_AWADDR,
	fib_40_m_axi_gmem_AWLEN,
	fib_40_m_axi_gmem_AWSIZE,
	fib_40_m_axi_gmem_AWBURST,
	fib_40_m_axi_gmem_AWLOCK,
	fib_40_m_axi_gmem_AWCACHE,
	fib_40_m_axi_gmem_AWPROT,
	fib_40_m_axi_gmem_AWQOS,
	fib_40_m_axi_gmem_AWREGION,
	fib_40_m_axi_gmem_AWUSER,
	fib_40_m_axi_gmem_WREADY,
	fib_40_m_axi_gmem_WVALID,
	fib_40_m_axi_gmem_WDATA,
	fib_40_m_axi_gmem_WSTRB,
	fib_40_m_axi_gmem_WLAST,
	fib_40_m_axi_gmem_WUSER,
	fib_40_m_axi_gmem_BREADY,
	fib_40_m_axi_gmem_BVALID,
	fib_40_m_axi_gmem_BID,
	fib_40_m_axi_gmem_BRESP,
	fib_40_m_axi_gmem_BUSER,
	fib_40_s_axi_control_ARREADY,
	fib_40_s_axi_control_ARVALID,
	fib_40_s_axi_control_ARADDR,
	fib_40_s_axi_control_RREADY,
	fib_40_s_axi_control_RVALID,
	fib_40_s_axi_control_RDATA,
	fib_40_s_axi_control_RRESP,
	fib_40_s_axi_control_AWREADY,
	fib_40_s_axi_control_AWVALID,
	fib_40_s_axi_control_AWADDR,
	fib_40_s_axi_control_WREADY,
	fib_40_s_axi_control_WVALID,
	fib_40_s_axi_control_WDATA,
	fib_40_s_axi_control_WSTRB,
	fib_40_s_axi_control_BREADY,
	fib_40_s_axi_control_BVALID,
	fib_40_s_axi_control_BRESP,
	fib_41_m_axi_gmem_ARREADY,
	fib_41_m_axi_gmem_ARVALID,
	fib_41_m_axi_gmem_ARID,
	fib_41_m_axi_gmem_ARADDR,
	fib_41_m_axi_gmem_ARLEN,
	fib_41_m_axi_gmem_ARSIZE,
	fib_41_m_axi_gmem_ARBURST,
	fib_41_m_axi_gmem_ARLOCK,
	fib_41_m_axi_gmem_ARCACHE,
	fib_41_m_axi_gmem_ARPROT,
	fib_41_m_axi_gmem_ARQOS,
	fib_41_m_axi_gmem_ARREGION,
	fib_41_m_axi_gmem_ARUSER,
	fib_41_m_axi_gmem_RREADY,
	fib_41_m_axi_gmem_RVALID,
	fib_41_m_axi_gmem_RID,
	fib_41_m_axi_gmem_RDATA,
	fib_41_m_axi_gmem_RRESP,
	fib_41_m_axi_gmem_RLAST,
	fib_41_m_axi_gmem_RUSER,
	fib_41_m_axi_gmem_AWREADY,
	fib_41_m_axi_gmem_AWVALID,
	fib_41_m_axi_gmem_AWID,
	fib_41_m_axi_gmem_AWADDR,
	fib_41_m_axi_gmem_AWLEN,
	fib_41_m_axi_gmem_AWSIZE,
	fib_41_m_axi_gmem_AWBURST,
	fib_41_m_axi_gmem_AWLOCK,
	fib_41_m_axi_gmem_AWCACHE,
	fib_41_m_axi_gmem_AWPROT,
	fib_41_m_axi_gmem_AWQOS,
	fib_41_m_axi_gmem_AWREGION,
	fib_41_m_axi_gmem_AWUSER,
	fib_41_m_axi_gmem_WREADY,
	fib_41_m_axi_gmem_WVALID,
	fib_41_m_axi_gmem_WDATA,
	fib_41_m_axi_gmem_WSTRB,
	fib_41_m_axi_gmem_WLAST,
	fib_41_m_axi_gmem_WUSER,
	fib_41_m_axi_gmem_BREADY,
	fib_41_m_axi_gmem_BVALID,
	fib_41_m_axi_gmem_BID,
	fib_41_m_axi_gmem_BRESP,
	fib_41_m_axi_gmem_BUSER,
	fib_41_s_axi_control_ARREADY,
	fib_41_s_axi_control_ARVALID,
	fib_41_s_axi_control_ARADDR,
	fib_41_s_axi_control_RREADY,
	fib_41_s_axi_control_RVALID,
	fib_41_s_axi_control_RDATA,
	fib_41_s_axi_control_RRESP,
	fib_41_s_axi_control_AWREADY,
	fib_41_s_axi_control_AWVALID,
	fib_41_s_axi_control_AWADDR,
	fib_41_s_axi_control_WREADY,
	fib_41_s_axi_control_WVALID,
	fib_41_s_axi_control_WDATA,
	fib_41_s_axi_control_WSTRB,
	fib_41_s_axi_control_BREADY,
	fib_41_s_axi_control_BVALID,
	fib_41_s_axi_control_BRESP,
	fib_42_m_axi_gmem_ARREADY,
	fib_42_m_axi_gmem_ARVALID,
	fib_42_m_axi_gmem_ARID,
	fib_42_m_axi_gmem_ARADDR,
	fib_42_m_axi_gmem_ARLEN,
	fib_42_m_axi_gmem_ARSIZE,
	fib_42_m_axi_gmem_ARBURST,
	fib_42_m_axi_gmem_ARLOCK,
	fib_42_m_axi_gmem_ARCACHE,
	fib_42_m_axi_gmem_ARPROT,
	fib_42_m_axi_gmem_ARQOS,
	fib_42_m_axi_gmem_ARREGION,
	fib_42_m_axi_gmem_ARUSER,
	fib_42_m_axi_gmem_RREADY,
	fib_42_m_axi_gmem_RVALID,
	fib_42_m_axi_gmem_RID,
	fib_42_m_axi_gmem_RDATA,
	fib_42_m_axi_gmem_RRESP,
	fib_42_m_axi_gmem_RLAST,
	fib_42_m_axi_gmem_RUSER,
	fib_42_m_axi_gmem_AWREADY,
	fib_42_m_axi_gmem_AWVALID,
	fib_42_m_axi_gmem_AWID,
	fib_42_m_axi_gmem_AWADDR,
	fib_42_m_axi_gmem_AWLEN,
	fib_42_m_axi_gmem_AWSIZE,
	fib_42_m_axi_gmem_AWBURST,
	fib_42_m_axi_gmem_AWLOCK,
	fib_42_m_axi_gmem_AWCACHE,
	fib_42_m_axi_gmem_AWPROT,
	fib_42_m_axi_gmem_AWQOS,
	fib_42_m_axi_gmem_AWREGION,
	fib_42_m_axi_gmem_AWUSER,
	fib_42_m_axi_gmem_WREADY,
	fib_42_m_axi_gmem_WVALID,
	fib_42_m_axi_gmem_WDATA,
	fib_42_m_axi_gmem_WSTRB,
	fib_42_m_axi_gmem_WLAST,
	fib_42_m_axi_gmem_WUSER,
	fib_42_m_axi_gmem_BREADY,
	fib_42_m_axi_gmem_BVALID,
	fib_42_m_axi_gmem_BID,
	fib_42_m_axi_gmem_BRESP,
	fib_42_m_axi_gmem_BUSER,
	fib_42_s_axi_control_ARREADY,
	fib_42_s_axi_control_ARVALID,
	fib_42_s_axi_control_ARADDR,
	fib_42_s_axi_control_RREADY,
	fib_42_s_axi_control_RVALID,
	fib_42_s_axi_control_RDATA,
	fib_42_s_axi_control_RRESP,
	fib_42_s_axi_control_AWREADY,
	fib_42_s_axi_control_AWVALID,
	fib_42_s_axi_control_AWADDR,
	fib_42_s_axi_control_WREADY,
	fib_42_s_axi_control_WVALID,
	fib_42_s_axi_control_WDATA,
	fib_42_s_axi_control_WSTRB,
	fib_42_s_axi_control_BREADY,
	fib_42_s_axi_control_BVALID,
	fib_42_s_axi_control_BRESP,
	fib_43_m_axi_gmem_ARREADY,
	fib_43_m_axi_gmem_ARVALID,
	fib_43_m_axi_gmem_ARID,
	fib_43_m_axi_gmem_ARADDR,
	fib_43_m_axi_gmem_ARLEN,
	fib_43_m_axi_gmem_ARSIZE,
	fib_43_m_axi_gmem_ARBURST,
	fib_43_m_axi_gmem_ARLOCK,
	fib_43_m_axi_gmem_ARCACHE,
	fib_43_m_axi_gmem_ARPROT,
	fib_43_m_axi_gmem_ARQOS,
	fib_43_m_axi_gmem_ARREGION,
	fib_43_m_axi_gmem_ARUSER,
	fib_43_m_axi_gmem_RREADY,
	fib_43_m_axi_gmem_RVALID,
	fib_43_m_axi_gmem_RID,
	fib_43_m_axi_gmem_RDATA,
	fib_43_m_axi_gmem_RRESP,
	fib_43_m_axi_gmem_RLAST,
	fib_43_m_axi_gmem_RUSER,
	fib_43_m_axi_gmem_AWREADY,
	fib_43_m_axi_gmem_AWVALID,
	fib_43_m_axi_gmem_AWID,
	fib_43_m_axi_gmem_AWADDR,
	fib_43_m_axi_gmem_AWLEN,
	fib_43_m_axi_gmem_AWSIZE,
	fib_43_m_axi_gmem_AWBURST,
	fib_43_m_axi_gmem_AWLOCK,
	fib_43_m_axi_gmem_AWCACHE,
	fib_43_m_axi_gmem_AWPROT,
	fib_43_m_axi_gmem_AWQOS,
	fib_43_m_axi_gmem_AWREGION,
	fib_43_m_axi_gmem_AWUSER,
	fib_43_m_axi_gmem_WREADY,
	fib_43_m_axi_gmem_WVALID,
	fib_43_m_axi_gmem_WDATA,
	fib_43_m_axi_gmem_WSTRB,
	fib_43_m_axi_gmem_WLAST,
	fib_43_m_axi_gmem_WUSER,
	fib_43_m_axi_gmem_BREADY,
	fib_43_m_axi_gmem_BVALID,
	fib_43_m_axi_gmem_BID,
	fib_43_m_axi_gmem_BRESP,
	fib_43_m_axi_gmem_BUSER,
	fib_43_s_axi_control_ARREADY,
	fib_43_s_axi_control_ARVALID,
	fib_43_s_axi_control_ARADDR,
	fib_43_s_axi_control_RREADY,
	fib_43_s_axi_control_RVALID,
	fib_43_s_axi_control_RDATA,
	fib_43_s_axi_control_RRESP,
	fib_43_s_axi_control_AWREADY,
	fib_43_s_axi_control_AWVALID,
	fib_43_s_axi_control_AWADDR,
	fib_43_s_axi_control_WREADY,
	fib_43_s_axi_control_WVALID,
	fib_43_s_axi_control_WDATA,
	fib_43_s_axi_control_WSTRB,
	fib_43_s_axi_control_BREADY,
	fib_43_s_axi_control_BVALID,
	fib_43_s_axi_control_BRESP,
	fib_44_m_axi_gmem_ARREADY,
	fib_44_m_axi_gmem_ARVALID,
	fib_44_m_axi_gmem_ARID,
	fib_44_m_axi_gmem_ARADDR,
	fib_44_m_axi_gmem_ARLEN,
	fib_44_m_axi_gmem_ARSIZE,
	fib_44_m_axi_gmem_ARBURST,
	fib_44_m_axi_gmem_ARLOCK,
	fib_44_m_axi_gmem_ARCACHE,
	fib_44_m_axi_gmem_ARPROT,
	fib_44_m_axi_gmem_ARQOS,
	fib_44_m_axi_gmem_ARREGION,
	fib_44_m_axi_gmem_ARUSER,
	fib_44_m_axi_gmem_RREADY,
	fib_44_m_axi_gmem_RVALID,
	fib_44_m_axi_gmem_RID,
	fib_44_m_axi_gmem_RDATA,
	fib_44_m_axi_gmem_RRESP,
	fib_44_m_axi_gmem_RLAST,
	fib_44_m_axi_gmem_RUSER,
	fib_44_m_axi_gmem_AWREADY,
	fib_44_m_axi_gmem_AWVALID,
	fib_44_m_axi_gmem_AWID,
	fib_44_m_axi_gmem_AWADDR,
	fib_44_m_axi_gmem_AWLEN,
	fib_44_m_axi_gmem_AWSIZE,
	fib_44_m_axi_gmem_AWBURST,
	fib_44_m_axi_gmem_AWLOCK,
	fib_44_m_axi_gmem_AWCACHE,
	fib_44_m_axi_gmem_AWPROT,
	fib_44_m_axi_gmem_AWQOS,
	fib_44_m_axi_gmem_AWREGION,
	fib_44_m_axi_gmem_AWUSER,
	fib_44_m_axi_gmem_WREADY,
	fib_44_m_axi_gmem_WVALID,
	fib_44_m_axi_gmem_WDATA,
	fib_44_m_axi_gmem_WSTRB,
	fib_44_m_axi_gmem_WLAST,
	fib_44_m_axi_gmem_WUSER,
	fib_44_m_axi_gmem_BREADY,
	fib_44_m_axi_gmem_BVALID,
	fib_44_m_axi_gmem_BID,
	fib_44_m_axi_gmem_BRESP,
	fib_44_m_axi_gmem_BUSER,
	fib_44_s_axi_control_ARREADY,
	fib_44_s_axi_control_ARVALID,
	fib_44_s_axi_control_ARADDR,
	fib_44_s_axi_control_RREADY,
	fib_44_s_axi_control_RVALID,
	fib_44_s_axi_control_RDATA,
	fib_44_s_axi_control_RRESP,
	fib_44_s_axi_control_AWREADY,
	fib_44_s_axi_control_AWVALID,
	fib_44_s_axi_control_AWADDR,
	fib_44_s_axi_control_WREADY,
	fib_44_s_axi_control_WVALID,
	fib_44_s_axi_control_WDATA,
	fib_44_s_axi_control_WSTRB,
	fib_44_s_axi_control_BREADY,
	fib_44_s_axi_control_BVALID,
	fib_44_s_axi_control_BRESP,
	fib_45_m_axi_gmem_ARREADY,
	fib_45_m_axi_gmem_ARVALID,
	fib_45_m_axi_gmem_ARID,
	fib_45_m_axi_gmem_ARADDR,
	fib_45_m_axi_gmem_ARLEN,
	fib_45_m_axi_gmem_ARSIZE,
	fib_45_m_axi_gmem_ARBURST,
	fib_45_m_axi_gmem_ARLOCK,
	fib_45_m_axi_gmem_ARCACHE,
	fib_45_m_axi_gmem_ARPROT,
	fib_45_m_axi_gmem_ARQOS,
	fib_45_m_axi_gmem_ARREGION,
	fib_45_m_axi_gmem_ARUSER,
	fib_45_m_axi_gmem_RREADY,
	fib_45_m_axi_gmem_RVALID,
	fib_45_m_axi_gmem_RID,
	fib_45_m_axi_gmem_RDATA,
	fib_45_m_axi_gmem_RRESP,
	fib_45_m_axi_gmem_RLAST,
	fib_45_m_axi_gmem_RUSER,
	fib_45_m_axi_gmem_AWREADY,
	fib_45_m_axi_gmem_AWVALID,
	fib_45_m_axi_gmem_AWID,
	fib_45_m_axi_gmem_AWADDR,
	fib_45_m_axi_gmem_AWLEN,
	fib_45_m_axi_gmem_AWSIZE,
	fib_45_m_axi_gmem_AWBURST,
	fib_45_m_axi_gmem_AWLOCK,
	fib_45_m_axi_gmem_AWCACHE,
	fib_45_m_axi_gmem_AWPROT,
	fib_45_m_axi_gmem_AWQOS,
	fib_45_m_axi_gmem_AWREGION,
	fib_45_m_axi_gmem_AWUSER,
	fib_45_m_axi_gmem_WREADY,
	fib_45_m_axi_gmem_WVALID,
	fib_45_m_axi_gmem_WDATA,
	fib_45_m_axi_gmem_WSTRB,
	fib_45_m_axi_gmem_WLAST,
	fib_45_m_axi_gmem_WUSER,
	fib_45_m_axi_gmem_BREADY,
	fib_45_m_axi_gmem_BVALID,
	fib_45_m_axi_gmem_BID,
	fib_45_m_axi_gmem_BRESP,
	fib_45_m_axi_gmem_BUSER,
	fib_45_s_axi_control_ARREADY,
	fib_45_s_axi_control_ARVALID,
	fib_45_s_axi_control_ARADDR,
	fib_45_s_axi_control_RREADY,
	fib_45_s_axi_control_RVALID,
	fib_45_s_axi_control_RDATA,
	fib_45_s_axi_control_RRESP,
	fib_45_s_axi_control_AWREADY,
	fib_45_s_axi_control_AWVALID,
	fib_45_s_axi_control_AWADDR,
	fib_45_s_axi_control_WREADY,
	fib_45_s_axi_control_WVALID,
	fib_45_s_axi_control_WDATA,
	fib_45_s_axi_control_WSTRB,
	fib_45_s_axi_control_BREADY,
	fib_45_s_axi_control_BVALID,
	fib_45_s_axi_control_BRESP,
	fib_46_m_axi_gmem_ARREADY,
	fib_46_m_axi_gmem_ARVALID,
	fib_46_m_axi_gmem_ARID,
	fib_46_m_axi_gmem_ARADDR,
	fib_46_m_axi_gmem_ARLEN,
	fib_46_m_axi_gmem_ARSIZE,
	fib_46_m_axi_gmem_ARBURST,
	fib_46_m_axi_gmem_ARLOCK,
	fib_46_m_axi_gmem_ARCACHE,
	fib_46_m_axi_gmem_ARPROT,
	fib_46_m_axi_gmem_ARQOS,
	fib_46_m_axi_gmem_ARREGION,
	fib_46_m_axi_gmem_ARUSER,
	fib_46_m_axi_gmem_RREADY,
	fib_46_m_axi_gmem_RVALID,
	fib_46_m_axi_gmem_RID,
	fib_46_m_axi_gmem_RDATA,
	fib_46_m_axi_gmem_RRESP,
	fib_46_m_axi_gmem_RLAST,
	fib_46_m_axi_gmem_RUSER,
	fib_46_m_axi_gmem_AWREADY,
	fib_46_m_axi_gmem_AWVALID,
	fib_46_m_axi_gmem_AWID,
	fib_46_m_axi_gmem_AWADDR,
	fib_46_m_axi_gmem_AWLEN,
	fib_46_m_axi_gmem_AWSIZE,
	fib_46_m_axi_gmem_AWBURST,
	fib_46_m_axi_gmem_AWLOCK,
	fib_46_m_axi_gmem_AWCACHE,
	fib_46_m_axi_gmem_AWPROT,
	fib_46_m_axi_gmem_AWQOS,
	fib_46_m_axi_gmem_AWREGION,
	fib_46_m_axi_gmem_AWUSER,
	fib_46_m_axi_gmem_WREADY,
	fib_46_m_axi_gmem_WVALID,
	fib_46_m_axi_gmem_WDATA,
	fib_46_m_axi_gmem_WSTRB,
	fib_46_m_axi_gmem_WLAST,
	fib_46_m_axi_gmem_WUSER,
	fib_46_m_axi_gmem_BREADY,
	fib_46_m_axi_gmem_BVALID,
	fib_46_m_axi_gmem_BID,
	fib_46_m_axi_gmem_BRESP,
	fib_46_m_axi_gmem_BUSER,
	fib_46_s_axi_control_ARREADY,
	fib_46_s_axi_control_ARVALID,
	fib_46_s_axi_control_ARADDR,
	fib_46_s_axi_control_RREADY,
	fib_46_s_axi_control_RVALID,
	fib_46_s_axi_control_RDATA,
	fib_46_s_axi_control_RRESP,
	fib_46_s_axi_control_AWREADY,
	fib_46_s_axi_control_AWVALID,
	fib_46_s_axi_control_AWADDR,
	fib_46_s_axi_control_WREADY,
	fib_46_s_axi_control_WVALID,
	fib_46_s_axi_control_WDATA,
	fib_46_s_axi_control_WSTRB,
	fib_46_s_axi_control_BREADY,
	fib_46_s_axi_control_BVALID,
	fib_46_s_axi_control_BRESP,
	fib_47_m_axi_gmem_ARREADY,
	fib_47_m_axi_gmem_ARVALID,
	fib_47_m_axi_gmem_ARID,
	fib_47_m_axi_gmem_ARADDR,
	fib_47_m_axi_gmem_ARLEN,
	fib_47_m_axi_gmem_ARSIZE,
	fib_47_m_axi_gmem_ARBURST,
	fib_47_m_axi_gmem_ARLOCK,
	fib_47_m_axi_gmem_ARCACHE,
	fib_47_m_axi_gmem_ARPROT,
	fib_47_m_axi_gmem_ARQOS,
	fib_47_m_axi_gmem_ARREGION,
	fib_47_m_axi_gmem_ARUSER,
	fib_47_m_axi_gmem_RREADY,
	fib_47_m_axi_gmem_RVALID,
	fib_47_m_axi_gmem_RID,
	fib_47_m_axi_gmem_RDATA,
	fib_47_m_axi_gmem_RRESP,
	fib_47_m_axi_gmem_RLAST,
	fib_47_m_axi_gmem_RUSER,
	fib_47_m_axi_gmem_AWREADY,
	fib_47_m_axi_gmem_AWVALID,
	fib_47_m_axi_gmem_AWID,
	fib_47_m_axi_gmem_AWADDR,
	fib_47_m_axi_gmem_AWLEN,
	fib_47_m_axi_gmem_AWSIZE,
	fib_47_m_axi_gmem_AWBURST,
	fib_47_m_axi_gmem_AWLOCK,
	fib_47_m_axi_gmem_AWCACHE,
	fib_47_m_axi_gmem_AWPROT,
	fib_47_m_axi_gmem_AWQOS,
	fib_47_m_axi_gmem_AWREGION,
	fib_47_m_axi_gmem_AWUSER,
	fib_47_m_axi_gmem_WREADY,
	fib_47_m_axi_gmem_WVALID,
	fib_47_m_axi_gmem_WDATA,
	fib_47_m_axi_gmem_WSTRB,
	fib_47_m_axi_gmem_WLAST,
	fib_47_m_axi_gmem_WUSER,
	fib_47_m_axi_gmem_BREADY,
	fib_47_m_axi_gmem_BVALID,
	fib_47_m_axi_gmem_BID,
	fib_47_m_axi_gmem_BRESP,
	fib_47_m_axi_gmem_BUSER,
	fib_47_s_axi_control_ARREADY,
	fib_47_s_axi_control_ARVALID,
	fib_47_s_axi_control_ARADDR,
	fib_47_s_axi_control_RREADY,
	fib_47_s_axi_control_RVALID,
	fib_47_s_axi_control_RDATA,
	fib_47_s_axi_control_RRESP,
	fib_47_s_axi_control_AWREADY,
	fib_47_s_axi_control_AWVALID,
	fib_47_s_axi_control_AWADDR,
	fib_47_s_axi_control_WREADY,
	fib_47_s_axi_control_WVALID,
	fib_47_s_axi_control_WDATA,
	fib_47_s_axi_control_WSTRB,
	fib_47_s_axi_control_BREADY,
	fib_47_s_axi_control_BVALID,
	fib_47_s_axi_control_BRESP,
	fib_48_m_axi_gmem_ARREADY,
	fib_48_m_axi_gmem_ARVALID,
	fib_48_m_axi_gmem_ARID,
	fib_48_m_axi_gmem_ARADDR,
	fib_48_m_axi_gmem_ARLEN,
	fib_48_m_axi_gmem_ARSIZE,
	fib_48_m_axi_gmem_ARBURST,
	fib_48_m_axi_gmem_ARLOCK,
	fib_48_m_axi_gmem_ARCACHE,
	fib_48_m_axi_gmem_ARPROT,
	fib_48_m_axi_gmem_ARQOS,
	fib_48_m_axi_gmem_ARREGION,
	fib_48_m_axi_gmem_ARUSER,
	fib_48_m_axi_gmem_RREADY,
	fib_48_m_axi_gmem_RVALID,
	fib_48_m_axi_gmem_RID,
	fib_48_m_axi_gmem_RDATA,
	fib_48_m_axi_gmem_RRESP,
	fib_48_m_axi_gmem_RLAST,
	fib_48_m_axi_gmem_RUSER,
	fib_48_m_axi_gmem_AWREADY,
	fib_48_m_axi_gmem_AWVALID,
	fib_48_m_axi_gmem_AWID,
	fib_48_m_axi_gmem_AWADDR,
	fib_48_m_axi_gmem_AWLEN,
	fib_48_m_axi_gmem_AWSIZE,
	fib_48_m_axi_gmem_AWBURST,
	fib_48_m_axi_gmem_AWLOCK,
	fib_48_m_axi_gmem_AWCACHE,
	fib_48_m_axi_gmem_AWPROT,
	fib_48_m_axi_gmem_AWQOS,
	fib_48_m_axi_gmem_AWREGION,
	fib_48_m_axi_gmem_AWUSER,
	fib_48_m_axi_gmem_WREADY,
	fib_48_m_axi_gmem_WVALID,
	fib_48_m_axi_gmem_WDATA,
	fib_48_m_axi_gmem_WSTRB,
	fib_48_m_axi_gmem_WLAST,
	fib_48_m_axi_gmem_WUSER,
	fib_48_m_axi_gmem_BREADY,
	fib_48_m_axi_gmem_BVALID,
	fib_48_m_axi_gmem_BID,
	fib_48_m_axi_gmem_BRESP,
	fib_48_m_axi_gmem_BUSER,
	fib_48_s_axi_control_ARREADY,
	fib_48_s_axi_control_ARVALID,
	fib_48_s_axi_control_ARADDR,
	fib_48_s_axi_control_RREADY,
	fib_48_s_axi_control_RVALID,
	fib_48_s_axi_control_RDATA,
	fib_48_s_axi_control_RRESP,
	fib_48_s_axi_control_AWREADY,
	fib_48_s_axi_control_AWVALID,
	fib_48_s_axi_control_AWADDR,
	fib_48_s_axi_control_WREADY,
	fib_48_s_axi_control_WVALID,
	fib_48_s_axi_control_WDATA,
	fib_48_s_axi_control_WSTRB,
	fib_48_s_axi_control_BREADY,
	fib_48_s_axi_control_BVALID,
	fib_48_s_axi_control_BRESP,
	fib_49_m_axi_gmem_ARREADY,
	fib_49_m_axi_gmem_ARVALID,
	fib_49_m_axi_gmem_ARID,
	fib_49_m_axi_gmem_ARADDR,
	fib_49_m_axi_gmem_ARLEN,
	fib_49_m_axi_gmem_ARSIZE,
	fib_49_m_axi_gmem_ARBURST,
	fib_49_m_axi_gmem_ARLOCK,
	fib_49_m_axi_gmem_ARCACHE,
	fib_49_m_axi_gmem_ARPROT,
	fib_49_m_axi_gmem_ARQOS,
	fib_49_m_axi_gmem_ARREGION,
	fib_49_m_axi_gmem_ARUSER,
	fib_49_m_axi_gmem_RREADY,
	fib_49_m_axi_gmem_RVALID,
	fib_49_m_axi_gmem_RID,
	fib_49_m_axi_gmem_RDATA,
	fib_49_m_axi_gmem_RRESP,
	fib_49_m_axi_gmem_RLAST,
	fib_49_m_axi_gmem_RUSER,
	fib_49_m_axi_gmem_AWREADY,
	fib_49_m_axi_gmem_AWVALID,
	fib_49_m_axi_gmem_AWID,
	fib_49_m_axi_gmem_AWADDR,
	fib_49_m_axi_gmem_AWLEN,
	fib_49_m_axi_gmem_AWSIZE,
	fib_49_m_axi_gmem_AWBURST,
	fib_49_m_axi_gmem_AWLOCK,
	fib_49_m_axi_gmem_AWCACHE,
	fib_49_m_axi_gmem_AWPROT,
	fib_49_m_axi_gmem_AWQOS,
	fib_49_m_axi_gmem_AWREGION,
	fib_49_m_axi_gmem_AWUSER,
	fib_49_m_axi_gmem_WREADY,
	fib_49_m_axi_gmem_WVALID,
	fib_49_m_axi_gmem_WDATA,
	fib_49_m_axi_gmem_WSTRB,
	fib_49_m_axi_gmem_WLAST,
	fib_49_m_axi_gmem_WUSER,
	fib_49_m_axi_gmem_BREADY,
	fib_49_m_axi_gmem_BVALID,
	fib_49_m_axi_gmem_BID,
	fib_49_m_axi_gmem_BRESP,
	fib_49_m_axi_gmem_BUSER,
	fib_49_s_axi_control_ARREADY,
	fib_49_s_axi_control_ARVALID,
	fib_49_s_axi_control_ARADDR,
	fib_49_s_axi_control_RREADY,
	fib_49_s_axi_control_RVALID,
	fib_49_s_axi_control_RDATA,
	fib_49_s_axi_control_RRESP,
	fib_49_s_axi_control_AWREADY,
	fib_49_s_axi_control_AWVALID,
	fib_49_s_axi_control_AWADDR,
	fib_49_s_axi_control_WREADY,
	fib_49_s_axi_control_WVALID,
	fib_49_s_axi_control_WDATA,
	fib_49_s_axi_control_WSTRB,
	fib_49_s_axi_control_BREADY,
	fib_49_s_axi_control_BVALID,
	fib_49_s_axi_control_BRESP,
	fib_50_m_axi_gmem_ARREADY,
	fib_50_m_axi_gmem_ARVALID,
	fib_50_m_axi_gmem_ARID,
	fib_50_m_axi_gmem_ARADDR,
	fib_50_m_axi_gmem_ARLEN,
	fib_50_m_axi_gmem_ARSIZE,
	fib_50_m_axi_gmem_ARBURST,
	fib_50_m_axi_gmem_ARLOCK,
	fib_50_m_axi_gmem_ARCACHE,
	fib_50_m_axi_gmem_ARPROT,
	fib_50_m_axi_gmem_ARQOS,
	fib_50_m_axi_gmem_ARREGION,
	fib_50_m_axi_gmem_ARUSER,
	fib_50_m_axi_gmem_RREADY,
	fib_50_m_axi_gmem_RVALID,
	fib_50_m_axi_gmem_RID,
	fib_50_m_axi_gmem_RDATA,
	fib_50_m_axi_gmem_RRESP,
	fib_50_m_axi_gmem_RLAST,
	fib_50_m_axi_gmem_RUSER,
	fib_50_m_axi_gmem_AWREADY,
	fib_50_m_axi_gmem_AWVALID,
	fib_50_m_axi_gmem_AWID,
	fib_50_m_axi_gmem_AWADDR,
	fib_50_m_axi_gmem_AWLEN,
	fib_50_m_axi_gmem_AWSIZE,
	fib_50_m_axi_gmem_AWBURST,
	fib_50_m_axi_gmem_AWLOCK,
	fib_50_m_axi_gmem_AWCACHE,
	fib_50_m_axi_gmem_AWPROT,
	fib_50_m_axi_gmem_AWQOS,
	fib_50_m_axi_gmem_AWREGION,
	fib_50_m_axi_gmem_AWUSER,
	fib_50_m_axi_gmem_WREADY,
	fib_50_m_axi_gmem_WVALID,
	fib_50_m_axi_gmem_WDATA,
	fib_50_m_axi_gmem_WSTRB,
	fib_50_m_axi_gmem_WLAST,
	fib_50_m_axi_gmem_WUSER,
	fib_50_m_axi_gmem_BREADY,
	fib_50_m_axi_gmem_BVALID,
	fib_50_m_axi_gmem_BID,
	fib_50_m_axi_gmem_BRESP,
	fib_50_m_axi_gmem_BUSER,
	fib_50_s_axi_control_ARREADY,
	fib_50_s_axi_control_ARVALID,
	fib_50_s_axi_control_ARADDR,
	fib_50_s_axi_control_RREADY,
	fib_50_s_axi_control_RVALID,
	fib_50_s_axi_control_RDATA,
	fib_50_s_axi_control_RRESP,
	fib_50_s_axi_control_AWREADY,
	fib_50_s_axi_control_AWVALID,
	fib_50_s_axi_control_AWADDR,
	fib_50_s_axi_control_WREADY,
	fib_50_s_axi_control_WVALID,
	fib_50_s_axi_control_WDATA,
	fib_50_s_axi_control_WSTRB,
	fib_50_s_axi_control_BREADY,
	fib_50_s_axi_control_BVALID,
	fib_50_s_axi_control_BRESP,
	fib_51_m_axi_gmem_ARREADY,
	fib_51_m_axi_gmem_ARVALID,
	fib_51_m_axi_gmem_ARID,
	fib_51_m_axi_gmem_ARADDR,
	fib_51_m_axi_gmem_ARLEN,
	fib_51_m_axi_gmem_ARSIZE,
	fib_51_m_axi_gmem_ARBURST,
	fib_51_m_axi_gmem_ARLOCK,
	fib_51_m_axi_gmem_ARCACHE,
	fib_51_m_axi_gmem_ARPROT,
	fib_51_m_axi_gmem_ARQOS,
	fib_51_m_axi_gmem_ARREGION,
	fib_51_m_axi_gmem_ARUSER,
	fib_51_m_axi_gmem_RREADY,
	fib_51_m_axi_gmem_RVALID,
	fib_51_m_axi_gmem_RID,
	fib_51_m_axi_gmem_RDATA,
	fib_51_m_axi_gmem_RRESP,
	fib_51_m_axi_gmem_RLAST,
	fib_51_m_axi_gmem_RUSER,
	fib_51_m_axi_gmem_AWREADY,
	fib_51_m_axi_gmem_AWVALID,
	fib_51_m_axi_gmem_AWID,
	fib_51_m_axi_gmem_AWADDR,
	fib_51_m_axi_gmem_AWLEN,
	fib_51_m_axi_gmem_AWSIZE,
	fib_51_m_axi_gmem_AWBURST,
	fib_51_m_axi_gmem_AWLOCK,
	fib_51_m_axi_gmem_AWCACHE,
	fib_51_m_axi_gmem_AWPROT,
	fib_51_m_axi_gmem_AWQOS,
	fib_51_m_axi_gmem_AWREGION,
	fib_51_m_axi_gmem_AWUSER,
	fib_51_m_axi_gmem_WREADY,
	fib_51_m_axi_gmem_WVALID,
	fib_51_m_axi_gmem_WDATA,
	fib_51_m_axi_gmem_WSTRB,
	fib_51_m_axi_gmem_WLAST,
	fib_51_m_axi_gmem_WUSER,
	fib_51_m_axi_gmem_BREADY,
	fib_51_m_axi_gmem_BVALID,
	fib_51_m_axi_gmem_BID,
	fib_51_m_axi_gmem_BRESP,
	fib_51_m_axi_gmem_BUSER,
	fib_51_s_axi_control_ARREADY,
	fib_51_s_axi_control_ARVALID,
	fib_51_s_axi_control_ARADDR,
	fib_51_s_axi_control_RREADY,
	fib_51_s_axi_control_RVALID,
	fib_51_s_axi_control_RDATA,
	fib_51_s_axi_control_RRESP,
	fib_51_s_axi_control_AWREADY,
	fib_51_s_axi_control_AWVALID,
	fib_51_s_axi_control_AWADDR,
	fib_51_s_axi_control_WREADY,
	fib_51_s_axi_control_WVALID,
	fib_51_s_axi_control_WDATA,
	fib_51_s_axi_control_WSTRB,
	fib_51_s_axi_control_BREADY,
	fib_51_s_axi_control_BVALID,
	fib_51_s_axi_control_BRESP,
	fib_52_m_axi_gmem_ARREADY,
	fib_52_m_axi_gmem_ARVALID,
	fib_52_m_axi_gmem_ARID,
	fib_52_m_axi_gmem_ARADDR,
	fib_52_m_axi_gmem_ARLEN,
	fib_52_m_axi_gmem_ARSIZE,
	fib_52_m_axi_gmem_ARBURST,
	fib_52_m_axi_gmem_ARLOCK,
	fib_52_m_axi_gmem_ARCACHE,
	fib_52_m_axi_gmem_ARPROT,
	fib_52_m_axi_gmem_ARQOS,
	fib_52_m_axi_gmem_ARREGION,
	fib_52_m_axi_gmem_ARUSER,
	fib_52_m_axi_gmem_RREADY,
	fib_52_m_axi_gmem_RVALID,
	fib_52_m_axi_gmem_RID,
	fib_52_m_axi_gmem_RDATA,
	fib_52_m_axi_gmem_RRESP,
	fib_52_m_axi_gmem_RLAST,
	fib_52_m_axi_gmem_RUSER,
	fib_52_m_axi_gmem_AWREADY,
	fib_52_m_axi_gmem_AWVALID,
	fib_52_m_axi_gmem_AWID,
	fib_52_m_axi_gmem_AWADDR,
	fib_52_m_axi_gmem_AWLEN,
	fib_52_m_axi_gmem_AWSIZE,
	fib_52_m_axi_gmem_AWBURST,
	fib_52_m_axi_gmem_AWLOCK,
	fib_52_m_axi_gmem_AWCACHE,
	fib_52_m_axi_gmem_AWPROT,
	fib_52_m_axi_gmem_AWQOS,
	fib_52_m_axi_gmem_AWREGION,
	fib_52_m_axi_gmem_AWUSER,
	fib_52_m_axi_gmem_WREADY,
	fib_52_m_axi_gmem_WVALID,
	fib_52_m_axi_gmem_WDATA,
	fib_52_m_axi_gmem_WSTRB,
	fib_52_m_axi_gmem_WLAST,
	fib_52_m_axi_gmem_WUSER,
	fib_52_m_axi_gmem_BREADY,
	fib_52_m_axi_gmem_BVALID,
	fib_52_m_axi_gmem_BID,
	fib_52_m_axi_gmem_BRESP,
	fib_52_m_axi_gmem_BUSER,
	fib_52_s_axi_control_ARREADY,
	fib_52_s_axi_control_ARVALID,
	fib_52_s_axi_control_ARADDR,
	fib_52_s_axi_control_RREADY,
	fib_52_s_axi_control_RVALID,
	fib_52_s_axi_control_RDATA,
	fib_52_s_axi_control_RRESP,
	fib_52_s_axi_control_AWREADY,
	fib_52_s_axi_control_AWVALID,
	fib_52_s_axi_control_AWADDR,
	fib_52_s_axi_control_WREADY,
	fib_52_s_axi_control_WVALID,
	fib_52_s_axi_control_WDATA,
	fib_52_s_axi_control_WSTRB,
	fib_52_s_axi_control_BREADY,
	fib_52_s_axi_control_BVALID,
	fib_52_s_axi_control_BRESP,
	fib_53_m_axi_gmem_ARREADY,
	fib_53_m_axi_gmem_ARVALID,
	fib_53_m_axi_gmem_ARID,
	fib_53_m_axi_gmem_ARADDR,
	fib_53_m_axi_gmem_ARLEN,
	fib_53_m_axi_gmem_ARSIZE,
	fib_53_m_axi_gmem_ARBURST,
	fib_53_m_axi_gmem_ARLOCK,
	fib_53_m_axi_gmem_ARCACHE,
	fib_53_m_axi_gmem_ARPROT,
	fib_53_m_axi_gmem_ARQOS,
	fib_53_m_axi_gmem_ARREGION,
	fib_53_m_axi_gmem_ARUSER,
	fib_53_m_axi_gmem_RREADY,
	fib_53_m_axi_gmem_RVALID,
	fib_53_m_axi_gmem_RID,
	fib_53_m_axi_gmem_RDATA,
	fib_53_m_axi_gmem_RRESP,
	fib_53_m_axi_gmem_RLAST,
	fib_53_m_axi_gmem_RUSER,
	fib_53_m_axi_gmem_AWREADY,
	fib_53_m_axi_gmem_AWVALID,
	fib_53_m_axi_gmem_AWID,
	fib_53_m_axi_gmem_AWADDR,
	fib_53_m_axi_gmem_AWLEN,
	fib_53_m_axi_gmem_AWSIZE,
	fib_53_m_axi_gmem_AWBURST,
	fib_53_m_axi_gmem_AWLOCK,
	fib_53_m_axi_gmem_AWCACHE,
	fib_53_m_axi_gmem_AWPROT,
	fib_53_m_axi_gmem_AWQOS,
	fib_53_m_axi_gmem_AWREGION,
	fib_53_m_axi_gmem_AWUSER,
	fib_53_m_axi_gmem_WREADY,
	fib_53_m_axi_gmem_WVALID,
	fib_53_m_axi_gmem_WDATA,
	fib_53_m_axi_gmem_WSTRB,
	fib_53_m_axi_gmem_WLAST,
	fib_53_m_axi_gmem_WUSER,
	fib_53_m_axi_gmem_BREADY,
	fib_53_m_axi_gmem_BVALID,
	fib_53_m_axi_gmem_BID,
	fib_53_m_axi_gmem_BRESP,
	fib_53_m_axi_gmem_BUSER,
	fib_53_s_axi_control_ARREADY,
	fib_53_s_axi_control_ARVALID,
	fib_53_s_axi_control_ARADDR,
	fib_53_s_axi_control_RREADY,
	fib_53_s_axi_control_RVALID,
	fib_53_s_axi_control_RDATA,
	fib_53_s_axi_control_RRESP,
	fib_53_s_axi_control_AWREADY,
	fib_53_s_axi_control_AWVALID,
	fib_53_s_axi_control_AWADDR,
	fib_53_s_axi_control_WREADY,
	fib_53_s_axi_control_WVALID,
	fib_53_s_axi_control_WDATA,
	fib_53_s_axi_control_WSTRB,
	fib_53_s_axi_control_BREADY,
	fib_53_s_axi_control_BVALID,
	fib_53_s_axi_control_BRESP,
	fib_54_m_axi_gmem_ARREADY,
	fib_54_m_axi_gmem_ARVALID,
	fib_54_m_axi_gmem_ARID,
	fib_54_m_axi_gmem_ARADDR,
	fib_54_m_axi_gmem_ARLEN,
	fib_54_m_axi_gmem_ARSIZE,
	fib_54_m_axi_gmem_ARBURST,
	fib_54_m_axi_gmem_ARLOCK,
	fib_54_m_axi_gmem_ARCACHE,
	fib_54_m_axi_gmem_ARPROT,
	fib_54_m_axi_gmem_ARQOS,
	fib_54_m_axi_gmem_ARREGION,
	fib_54_m_axi_gmem_ARUSER,
	fib_54_m_axi_gmem_RREADY,
	fib_54_m_axi_gmem_RVALID,
	fib_54_m_axi_gmem_RID,
	fib_54_m_axi_gmem_RDATA,
	fib_54_m_axi_gmem_RRESP,
	fib_54_m_axi_gmem_RLAST,
	fib_54_m_axi_gmem_RUSER,
	fib_54_m_axi_gmem_AWREADY,
	fib_54_m_axi_gmem_AWVALID,
	fib_54_m_axi_gmem_AWID,
	fib_54_m_axi_gmem_AWADDR,
	fib_54_m_axi_gmem_AWLEN,
	fib_54_m_axi_gmem_AWSIZE,
	fib_54_m_axi_gmem_AWBURST,
	fib_54_m_axi_gmem_AWLOCK,
	fib_54_m_axi_gmem_AWCACHE,
	fib_54_m_axi_gmem_AWPROT,
	fib_54_m_axi_gmem_AWQOS,
	fib_54_m_axi_gmem_AWREGION,
	fib_54_m_axi_gmem_AWUSER,
	fib_54_m_axi_gmem_WREADY,
	fib_54_m_axi_gmem_WVALID,
	fib_54_m_axi_gmem_WDATA,
	fib_54_m_axi_gmem_WSTRB,
	fib_54_m_axi_gmem_WLAST,
	fib_54_m_axi_gmem_WUSER,
	fib_54_m_axi_gmem_BREADY,
	fib_54_m_axi_gmem_BVALID,
	fib_54_m_axi_gmem_BID,
	fib_54_m_axi_gmem_BRESP,
	fib_54_m_axi_gmem_BUSER,
	fib_54_s_axi_control_ARREADY,
	fib_54_s_axi_control_ARVALID,
	fib_54_s_axi_control_ARADDR,
	fib_54_s_axi_control_RREADY,
	fib_54_s_axi_control_RVALID,
	fib_54_s_axi_control_RDATA,
	fib_54_s_axi_control_RRESP,
	fib_54_s_axi_control_AWREADY,
	fib_54_s_axi_control_AWVALID,
	fib_54_s_axi_control_AWADDR,
	fib_54_s_axi_control_WREADY,
	fib_54_s_axi_control_WVALID,
	fib_54_s_axi_control_WDATA,
	fib_54_s_axi_control_WSTRB,
	fib_54_s_axi_control_BREADY,
	fib_54_s_axi_control_BVALID,
	fib_54_s_axi_control_BRESP,
	fib_55_m_axi_gmem_ARREADY,
	fib_55_m_axi_gmem_ARVALID,
	fib_55_m_axi_gmem_ARID,
	fib_55_m_axi_gmem_ARADDR,
	fib_55_m_axi_gmem_ARLEN,
	fib_55_m_axi_gmem_ARSIZE,
	fib_55_m_axi_gmem_ARBURST,
	fib_55_m_axi_gmem_ARLOCK,
	fib_55_m_axi_gmem_ARCACHE,
	fib_55_m_axi_gmem_ARPROT,
	fib_55_m_axi_gmem_ARQOS,
	fib_55_m_axi_gmem_ARREGION,
	fib_55_m_axi_gmem_ARUSER,
	fib_55_m_axi_gmem_RREADY,
	fib_55_m_axi_gmem_RVALID,
	fib_55_m_axi_gmem_RID,
	fib_55_m_axi_gmem_RDATA,
	fib_55_m_axi_gmem_RRESP,
	fib_55_m_axi_gmem_RLAST,
	fib_55_m_axi_gmem_RUSER,
	fib_55_m_axi_gmem_AWREADY,
	fib_55_m_axi_gmem_AWVALID,
	fib_55_m_axi_gmem_AWID,
	fib_55_m_axi_gmem_AWADDR,
	fib_55_m_axi_gmem_AWLEN,
	fib_55_m_axi_gmem_AWSIZE,
	fib_55_m_axi_gmem_AWBURST,
	fib_55_m_axi_gmem_AWLOCK,
	fib_55_m_axi_gmem_AWCACHE,
	fib_55_m_axi_gmem_AWPROT,
	fib_55_m_axi_gmem_AWQOS,
	fib_55_m_axi_gmem_AWREGION,
	fib_55_m_axi_gmem_AWUSER,
	fib_55_m_axi_gmem_WREADY,
	fib_55_m_axi_gmem_WVALID,
	fib_55_m_axi_gmem_WDATA,
	fib_55_m_axi_gmem_WSTRB,
	fib_55_m_axi_gmem_WLAST,
	fib_55_m_axi_gmem_WUSER,
	fib_55_m_axi_gmem_BREADY,
	fib_55_m_axi_gmem_BVALID,
	fib_55_m_axi_gmem_BID,
	fib_55_m_axi_gmem_BRESP,
	fib_55_m_axi_gmem_BUSER,
	fib_55_s_axi_control_ARREADY,
	fib_55_s_axi_control_ARVALID,
	fib_55_s_axi_control_ARADDR,
	fib_55_s_axi_control_RREADY,
	fib_55_s_axi_control_RVALID,
	fib_55_s_axi_control_RDATA,
	fib_55_s_axi_control_RRESP,
	fib_55_s_axi_control_AWREADY,
	fib_55_s_axi_control_AWVALID,
	fib_55_s_axi_control_AWADDR,
	fib_55_s_axi_control_WREADY,
	fib_55_s_axi_control_WVALID,
	fib_55_s_axi_control_WDATA,
	fib_55_s_axi_control_WSTRB,
	fib_55_s_axi_control_BREADY,
	fib_55_s_axi_control_BVALID,
	fib_55_s_axi_control_BRESP,
	fib_56_m_axi_gmem_ARREADY,
	fib_56_m_axi_gmem_ARVALID,
	fib_56_m_axi_gmem_ARID,
	fib_56_m_axi_gmem_ARADDR,
	fib_56_m_axi_gmem_ARLEN,
	fib_56_m_axi_gmem_ARSIZE,
	fib_56_m_axi_gmem_ARBURST,
	fib_56_m_axi_gmem_ARLOCK,
	fib_56_m_axi_gmem_ARCACHE,
	fib_56_m_axi_gmem_ARPROT,
	fib_56_m_axi_gmem_ARQOS,
	fib_56_m_axi_gmem_ARREGION,
	fib_56_m_axi_gmem_ARUSER,
	fib_56_m_axi_gmem_RREADY,
	fib_56_m_axi_gmem_RVALID,
	fib_56_m_axi_gmem_RID,
	fib_56_m_axi_gmem_RDATA,
	fib_56_m_axi_gmem_RRESP,
	fib_56_m_axi_gmem_RLAST,
	fib_56_m_axi_gmem_RUSER,
	fib_56_m_axi_gmem_AWREADY,
	fib_56_m_axi_gmem_AWVALID,
	fib_56_m_axi_gmem_AWID,
	fib_56_m_axi_gmem_AWADDR,
	fib_56_m_axi_gmem_AWLEN,
	fib_56_m_axi_gmem_AWSIZE,
	fib_56_m_axi_gmem_AWBURST,
	fib_56_m_axi_gmem_AWLOCK,
	fib_56_m_axi_gmem_AWCACHE,
	fib_56_m_axi_gmem_AWPROT,
	fib_56_m_axi_gmem_AWQOS,
	fib_56_m_axi_gmem_AWREGION,
	fib_56_m_axi_gmem_AWUSER,
	fib_56_m_axi_gmem_WREADY,
	fib_56_m_axi_gmem_WVALID,
	fib_56_m_axi_gmem_WDATA,
	fib_56_m_axi_gmem_WSTRB,
	fib_56_m_axi_gmem_WLAST,
	fib_56_m_axi_gmem_WUSER,
	fib_56_m_axi_gmem_BREADY,
	fib_56_m_axi_gmem_BVALID,
	fib_56_m_axi_gmem_BID,
	fib_56_m_axi_gmem_BRESP,
	fib_56_m_axi_gmem_BUSER,
	fib_56_s_axi_control_ARREADY,
	fib_56_s_axi_control_ARVALID,
	fib_56_s_axi_control_ARADDR,
	fib_56_s_axi_control_RREADY,
	fib_56_s_axi_control_RVALID,
	fib_56_s_axi_control_RDATA,
	fib_56_s_axi_control_RRESP,
	fib_56_s_axi_control_AWREADY,
	fib_56_s_axi_control_AWVALID,
	fib_56_s_axi_control_AWADDR,
	fib_56_s_axi_control_WREADY,
	fib_56_s_axi_control_WVALID,
	fib_56_s_axi_control_WDATA,
	fib_56_s_axi_control_WSTRB,
	fib_56_s_axi_control_BREADY,
	fib_56_s_axi_control_BVALID,
	fib_56_s_axi_control_BRESP,
	fib_57_m_axi_gmem_ARREADY,
	fib_57_m_axi_gmem_ARVALID,
	fib_57_m_axi_gmem_ARID,
	fib_57_m_axi_gmem_ARADDR,
	fib_57_m_axi_gmem_ARLEN,
	fib_57_m_axi_gmem_ARSIZE,
	fib_57_m_axi_gmem_ARBURST,
	fib_57_m_axi_gmem_ARLOCK,
	fib_57_m_axi_gmem_ARCACHE,
	fib_57_m_axi_gmem_ARPROT,
	fib_57_m_axi_gmem_ARQOS,
	fib_57_m_axi_gmem_ARREGION,
	fib_57_m_axi_gmem_ARUSER,
	fib_57_m_axi_gmem_RREADY,
	fib_57_m_axi_gmem_RVALID,
	fib_57_m_axi_gmem_RID,
	fib_57_m_axi_gmem_RDATA,
	fib_57_m_axi_gmem_RRESP,
	fib_57_m_axi_gmem_RLAST,
	fib_57_m_axi_gmem_RUSER,
	fib_57_m_axi_gmem_AWREADY,
	fib_57_m_axi_gmem_AWVALID,
	fib_57_m_axi_gmem_AWID,
	fib_57_m_axi_gmem_AWADDR,
	fib_57_m_axi_gmem_AWLEN,
	fib_57_m_axi_gmem_AWSIZE,
	fib_57_m_axi_gmem_AWBURST,
	fib_57_m_axi_gmem_AWLOCK,
	fib_57_m_axi_gmem_AWCACHE,
	fib_57_m_axi_gmem_AWPROT,
	fib_57_m_axi_gmem_AWQOS,
	fib_57_m_axi_gmem_AWREGION,
	fib_57_m_axi_gmem_AWUSER,
	fib_57_m_axi_gmem_WREADY,
	fib_57_m_axi_gmem_WVALID,
	fib_57_m_axi_gmem_WDATA,
	fib_57_m_axi_gmem_WSTRB,
	fib_57_m_axi_gmem_WLAST,
	fib_57_m_axi_gmem_WUSER,
	fib_57_m_axi_gmem_BREADY,
	fib_57_m_axi_gmem_BVALID,
	fib_57_m_axi_gmem_BID,
	fib_57_m_axi_gmem_BRESP,
	fib_57_m_axi_gmem_BUSER,
	fib_57_s_axi_control_ARREADY,
	fib_57_s_axi_control_ARVALID,
	fib_57_s_axi_control_ARADDR,
	fib_57_s_axi_control_RREADY,
	fib_57_s_axi_control_RVALID,
	fib_57_s_axi_control_RDATA,
	fib_57_s_axi_control_RRESP,
	fib_57_s_axi_control_AWREADY,
	fib_57_s_axi_control_AWVALID,
	fib_57_s_axi_control_AWADDR,
	fib_57_s_axi_control_WREADY,
	fib_57_s_axi_control_WVALID,
	fib_57_s_axi_control_WDATA,
	fib_57_s_axi_control_WSTRB,
	fib_57_s_axi_control_BREADY,
	fib_57_s_axi_control_BVALID,
	fib_57_s_axi_control_BRESP,
	fib_58_m_axi_gmem_ARREADY,
	fib_58_m_axi_gmem_ARVALID,
	fib_58_m_axi_gmem_ARID,
	fib_58_m_axi_gmem_ARADDR,
	fib_58_m_axi_gmem_ARLEN,
	fib_58_m_axi_gmem_ARSIZE,
	fib_58_m_axi_gmem_ARBURST,
	fib_58_m_axi_gmem_ARLOCK,
	fib_58_m_axi_gmem_ARCACHE,
	fib_58_m_axi_gmem_ARPROT,
	fib_58_m_axi_gmem_ARQOS,
	fib_58_m_axi_gmem_ARREGION,
	fib_58_m_axi_gmem_ARUSER,
	fib_58_m_axi_gmem_RREADY,
	fib_58_m_axi_gmem_RVALID,
	fib_58_m_axi_gmem_RID,
	fib_58_m_axi_gmem_RDATA,
	fib_58_m_axi_gmem_RRESP,
	fib_58_m_axi_gmem_RLAST,
	fib_58_m_axi_gmem_RUSER,
	fib_58_m_axi_gmem_AWREADY,
	fib_58_m_axi_gmem_AWVALID,
	fib_58_m_axi_gmem_AWID,
	fib_58_m_axi_gmem_AWADDR,
	fib_58_m_axi_gmem_AWLEN,
	fib_58_m_axi_gmem_AWSIZE,
	fib_58_m_axi_gmem_AWBURST,
	fib_58_m_axi_gmem_AWLOCK,
	fib_58_m_axi_gmem_AWCACHE,
	fib_58_m_axi_gmem_AWPROT,
	fib_58_m_axi_gmem_AWQOS,
	fib_58_m_axi_gmem_AWREGION,
	fib_58_m_axi_gmem_AWUSER,
	fib_58_m_axi_gmem_WREADY,
	fib_58_m_axi_gmem_WVALID,
	fib_58_m_axi_gmem_WDATA,
	fib_58_m_axi_gmem_WSTRB,
	fib_58_m_axi_gmem_WLAST,
	fib_58_m_axi_gmem_WUSER,
	fib_58_m_axi_gmem_BREADY,
	fib_58_m_axi_gmem_BVALID,
	fib_58_m_axi_gmem_BID,
	fib_58_m_axi_gmem_BRESP,
	fib_58_m_axi_gmem_BUSER,
	fib_58_s_axi_control_ARREADY,
	fib_58_s_axi_control_ARVALID,
	fib_58_s_axi_control_ARADDR,
	fib_58_s_axi_control_RREADY,
	fib_58_s_axi_control_RVALID,
	fib_58_s_axi_control_RDATA,
	fib_58_s_axi_control_RRESP,
	fib_58_s_axi_control_AWREADY,
	fib_58_s_axi_control_AWVALID,
	fib_58_s_axi_control_AWADDR,
	fib_58_s_axi_control_WREADY,
	fib_58_s_axi_control_WVALID,
	fib_58_s_axi_control_WDATA,
	fib_58_s_axi_control_WSTRB,
	fib_58_s_axi_control_BREADY,
	fib_58_s_axi_control_BVALID,
	fib_58_s_axi_control_BRESP,
	fib_59_m_axi_gmem_ARREADY,
	fib_59_m_axi_gmem_ARVALID,
	fib_59_m_axi_gmem_ARID,
	fib_59_m_axi_gmem_ARADDR,
	fib_59_m_axi_gmem_ARLEN,
	fib_59_m_axi_gmem_ARSIZE,
	fib_59_m_axi_gmem_ARBURST,
	fib_59_m_axi_gmem_ARLOCK,
	fib_59_m_axi_gmem_ARCACHE,
	fib_59_m_axi_gmem_ARPROT,
	fib_59_m_axi_gmem_ARQOS,
	fib_59_m_axi_gmem_ARREGION,
	fib_59_m_axi_gmem_ARUSER,
	fib_59_m_axi_gmem_RREADY,
	fib_59_m_axi_gmem_RVALID,
	fib_59_m_axi_gmem_RID,
	fib_59_m_axi_gmem_RDATA,
	fib_59_m_axi_gmem_RRESP,
	fib_59_m_axi_gmem_RLAST,
	fib_59_m_axi_gmem_RUSER,
	fib_59_m_axi_gmem_AWREADY,
	fib_59_m_axi_gmem_AWVALID,
	fib_59_m_axi_gmem_AWID,
	fib_59_m_axi_gmem_AWADDR,
	fib_59_m_axi_gmem_AWLEN,
	fib_59_m_axi_gmem_AWSIZE,
	fib_59_m_axi_gmem_AWBURST,
	fib_59_m_axi_gmem_AWLOCK,
	fib_59_m_axi_gmem_AWCACHE,
	fib_59_m_axi_gmem_AWPROT,
	fib_59_m_axi_gmem_AWQOS,
	fib_59_m_axi_gmem_AWREGION,
	fib_59_m_axi_gmem_AWUSER,
	fib_59_m_axi_gmem_WREADY,
	fib_59_m_axi_gmem_WVALID,
	fib_59_m_axi_gmem_WDATA,
	fib_59_m_axi_gmem_WSTRB,
	fib_59_m_axi_gmem_WLAST,
	fib_59_m_axi_gmem_WUSER,
	fib_59_m_axi_gmem_BREADY,
	fib_59_m_axi_gmem_BVALID,
	fib_59_m_axi_gmem_BID,
	fib_59_m_axi_gmem_BRESP,
	fib_59_m_axi_gmem_BUSER,
	fib_59_s_axi_control_ARREADY,
	fib_59_s_axi_control_ARVALID,
	fib_59_s_axi_control_ARADDR,
	fib_59_s_axi_control_RREADY,
	fib_59_s_axi_control_RVALID,
	fib_59_s_axi_control_RDATA,
	fib_59_s_axi_control_RRESP,
	fib_59_s_axi_control_AWREADY,
	fib_59_s_axi_control_AWVALID,
	fib_59_s_axi_control_AWADDR,
	fib_59_s_axi_control_WREADY,
	fib_59_s_axi_control_WVALID,
	fib_59_s_axi_control_WDATA,
	fib_59_s_axi_control_WSTRB,
	fib_59_s_axi_control_BREADY,
	fib_59_s_axi_control_BVALID,
	fib_59_s_axi_control_BRESP,
	fib_60_m_axi_gmem_ARREADY,
	fib_60_m_axi_gmem_ARVALID,
	fib_60_m_axi_gmem_ARID,
	fib_60_m_axi_gmem_ARADDR,
	fib_60_m_axi_gmem_ARLEN,
	fib_60_m_axi_gmem_ARSIZE,
	fib_60_m_axi_gmem_ARBURST,
	fib_60_m_axi_gmem_ARLOCK,
	fib_60_m_axi_gmem_ARCACHE,
	fib_60_m_axi_gmem_ARPROT,
	fib_60_m_axi_gmem_ARQOS,
	fib_60_m_axi_gmem_ARREGION,
	fib_60_m_axi_gmem_ARUSER,
	fib_60_m_axi_gmem_RREADY,
	fib_60_m_axi_gmem_RVALID,
	fib_60_m_axi_gmem_RID,
	fib_60_m_axi_gmem_RDATA,
	fib_60_m_axi_gmem_RRESP,
	fib_60_m_axi_gmem_RLAST,
	fib_60_m_axi_gmem_RUSER,
	fib_60_m_axi_gmem_AWREADY,
	fib_60_m_axi_gmem_AWVALID,
	fib_60_m_axi_gmem_AWID,
	fib_60_m_axi_gmem_AWADDR,
	fib_60_m_axi_gmem_AWLEN,
	fib_60_m_axi_gmem_AWSIZE,
	fib_60_m_axi_gmem_AWBURST,
	fib_60_m_axi_gmem_AWLOCK,
	fib_60_m_axi_gmem_AWCACHE,
	fib_60_m_axi_gmem_AWPROT,
	fib_60_m_axi_gmem_AWQOS,
	fib_60_m_axi_gmem_AWREGION,
	fib_60_m_axi_gmem_AWUSER,
	fib_60_m_axi_gmem_WREADY,
	fib_60_m_axi_gmem_WVALID,
	fib_60_m_axi_gmem_WDATA,
	fib_60_m_axi_gmem_WSTRB,
	fib_60_m_axi_gmem_WLAST,
	fib_60_m_axi_gmem_WUSER,
	fib_60_m_axi_gmem_BREADY,
	fib_60_m_axi_gmem_BVALID,
	fib_60_m_axi_gmem_BID,
	fib_60_m_axi_gmem_BRESP,
	fib_60_m_axi_gmem_BUSER,
	fib_60_s_axi_control_ARREADY,
	fib_60_s_axi_control_ARVALID,
	fib_60_s_axi_control_ARADDR,
	fib_60_s_axi_control_RREADY,
	fib_60_s_axi_control_RVALID,
	fib_60_s_axi_control_RDATA,
	fib_60_s_axi_control_RRESP,
	fib_60_s_axi_control_AWREADY,
	fib_60_s_axi_control_AWVALID,
	fib_60_s_axi_control_AWADDR,
	fib_60_s_axi_control_WREADY,
	fib_60_s_axi_control_WVALID,
	fib_60_s_axi_control_WDATA,
	fib_60_s_axi_control_WSTRB,
	fib_60_s_axi_control_BREADY,
	fib_60_s_axi_control_BVALID,
	fib_60_s_axi_control_BRESP,
	fib_61_m_axi_gmem_ARREADY,
	fib_61_m_axi_gmem_ARVALID,
	fib_61_m_axi_gmem_ARID,
	fib_61_m_axi_gmem_ARADDR,
	fib_61_m_axi_gmem_ARLEN,
	fib_61_m_axi_gmem_ARSIZE,
	fib_61_m_axi_gmem_ARBURST,
	fib_61_m_axi_gmem_ARLOCK,
	fib_61_m_axi_gmem_ARCACHE,
	fib_61_m_axi_gmem_ARPROT,
	fib_61_m_axi_gmem_ARQOS,
	fib_61_m_axi_gmem_ARREGION,
	fib_61_m_axi_gmem_ARUSER,
	fib_61_m_axi_gmem_RREADY,
	fib_61_m_axi_gmem_RVALID,
	fib_61_m_axi_gmem_RID,
	fib_61_m_axi_gmem_RDATA,
	fib_61_m_axi_gmem_RRESP,
	fib_61_m_axi_gmem_RLAST,
	fib_61_m_axi_gmem_RUSER,
	fib_61_m_axi_gmem_AWREADY,
	fib_61_m_axi_gmem_AWVALID,
	fib_61_m_axi_gmem_AWID,
	fib_61_m_axi_gmem_AWADDR,
	fib_61_m_axi_gmem_AWLEN,
	fib_61_m_axi_gmem_AWSIZE,
	fib_61_m_axi_gmem_AWBURST,
	fib_61_m_axi_gmem_AWLOCK,
	fib_61_m_axi_gmem_AWCACHE,
	fib_61_m_axi_gmem_AWPROT,
	fib_61_m_axi_gmem_AWQOS,
	fib_61_m_axi_gmem_AWREGION,
	fib_61_m_axi_gmem_AWUSER,
	fib_61_m_axi_gmem_WREADY,
	fib_61_m_axi_gmem_WVALID,
	fib_61_m_axi_gmem_WDATA,
	fib_61_m_axi_gmem_WSTRB,
	fib_61_m_axi_gmem_WLAST,
	fib_61_m_axi_gmem_WUSER,
	fib_61_m_axi_gmem_BREADY,
	fib_61_m_axi_gmem_BVALID,
	fib_61_m_axi_gmem_BID,
	fib_61_m_axi_gmem_BRESP,
	fib_61_m_axi_gmem_BUSER,
	fib_61_s_axi_control_ARREADY,
	fib_61_s_axi_control_ARVALID,
	fib_61_s_axi_control_ARADDR,
	fib_61_s_axi_control_RREADY,
	fib_61_s_axi_control_RVALID,
	fib_61_s_axi_control_RDATA,
	fib_61_s_axi_control_RRESP,
	fib_61_s_axi_control_AWREADY,
	fib_61_s_axi_control_AWVALID,
	fib_61_s_axi_control_AWADDR,
	fib_61_s_axi_control_WREADY,
	fib_61_s_axi_control_WVALID,
	fib_61_s_axi_control_WDATA,
	fib_61_s_axi_control_WSTRB,
	fib_61_s_axi_control_BREADY,
	fib_61_s_axi_control_BVALID,
	fib_61_s_axi_control_BRESP,
	fib_62_m_axi_gmem_ARREADY,
	fib_62_m_axi_gmem_ARVALID,
	fib_62_m_axi_gmem_ARID,
	fib_62_m_axi_gmem_ARADDR,
	fib_62_m_axi_gmem_ARLEN,
	fib_62_m_axi_gmem_ARSIZE,
	fib_62_m_axi_gmem_ARBURST,
	fib_62_m_axi_gmem_ARLOCK,
	fib_62_m_axi_gmem_ARCACHE,
	fib_62_m_axi_gmem_ARPROT,
	fib_62_m_axi_gmem_ARQOS,
	fib_62_m_axi_gmem_ARREGION,
	fib_62_m_axi_gmem_ARUSER,
	fib_62_m_axi_gmem_RREADY,
	fib_62_m_axi_gmem_RVALID,
	fib_62_m_axi_gmem_RID,
	fib_62_m_axi_gmem_RDATA,
	fib_62_m_axi_gmem_RRESP,
	fib_62_m_axi_gmem_RLAST,
	fib_62_m_axi_gmem_RUSER,
	fib_62_m_axi_gmem_AWREADY,
	fib_62_m_axi_gmem_AWVALID,
	fib_62_m_axi_gmem_AWID,
	fib_62_m_axi_gmem_AWADDR,
	fib_62_m_axi_gmem_AWLEN,
	fib_62_m_axi_gmem_AWSIZE,
	fib_62_m_axi_gmem_AWBURST,
	fib_62_m_axi_gmem_AWLOCK,
	fib_62_m_axi_gmem_AWCACHE,
	fib_62_m_axi_gmem_AWPROT,
	fib_62_m_axi_gmem_AWQOS,
	fib_62_m_axi_gmem_AWREGION,
	fib_62_m_axi_gmem_AWUSER,
	fib_62_m_axi_gmem_WREADY,
	fib_62_m_axi_gmem_WVALID,
	fib_62_m_axi_gmem_WDATA,
	fib_62_m_axi_gmem_WSTRB,
	fib_62_m_axi_gmem_WLAST,
	fib_62_m_axi_gmem_WUSER,
	fib_62_m_axi_gmem_BREADY,
	fib_62_m_axi_gmem_BVALID,
	fib_62_m_axi_gmem_BID,
	fib_62_m_axi_gmem_BRESP,
	fib_62_m_axi_gmem_BUSER,
	fib_62_s_axi_control_ARREADY,
	fib_62_s_axi_control_ARVALID,
	fib_62_s_axi_control_ARADDR,
	fib_62_s_axi_control_RREADY,
	fib_62_s_axi_control_RVALID,
	fib_62_s_axi_control_RDATA,
	fib_62_s_axi_control_RRESP,
	fib_62_s_axi_control_AWREADY,
	fib_62_s_axi_control_AWVALID,
	fib_62_s_axi_control_AWADDR,
	fib_62_s_axi_control_WREADY,
	fib_62_s_axi_control_WVALID,
	fib_62_s_axi_control_WDATA,
	fib_62_s_axi_control_WSTRB,
	fib_62_s_axi_control_BREADY,
	fib_62_s_axi_control_BVALID,
	fib_62_s_axi_control_BRESP,
	fib_63_m_axi_gmem_ARREADY,
	fib_63_m_axi_gmem_ARVALID,
	fib_63_m_axi_gmem_ARID,
	fib_63_m_axi_gmem_ARADDR,
	fib_63_m_axi_gmem_ARLEN,
	fib_63_m_axi_gmem_ARSIZE,
	fib_63_m_axi_gmem_ARBURST,
	fib_63_m_axi_gmem_ARLOCK,
	fib_63_m_axi_gmem_ARCACHE,
	fib_63_m_axi_gmem_ARPROT,
	fib_63_m_axi_gmem_ARQOS,
	fib_63_m_axi_gmem_ARREGION,
	fib_63_m_axi_gmem_ARUSER,
	fib_63_m_axi_gmem_RREADY,
	fib_63_m_axi_gmem_RVALID,
	fib_63_m_axi_gmem_RID,
	fib_63_m_axi_gmem_RDATA,
	fib_63_m_axi_gmem_RRESP,
	fib_63_m_axi_gmem_RLAST,
	fib_63_m_axi_gmem_RUSER,
	fib_63_m_axi_gmem_AWREADY,
	fib_63_m_axi_gmem_AWVALID,
	fib_63_m_axi_gmem_AWID,
	fib_63_m_axi_gmem_AWADDR,
	fib_63_m_axi_gmem_AWLEN,
	fib_63_m_axi_gmem_AWSIZE,
	fib_63_m_axi_gmem_AWBURST,
	fib_63_m_axi_gmem_AWLOCK,
	fib_63_m_axi_gmem_AWCACHE,
	fib_63_m_axi_gmem_AWPROT,
	fib_63_m_axi_gmem_AWQOS,
	fib_63_m_axi_gmem_AWREGION,
	fib_63_m_axi_gmem_AWUSER,
	fib_63_m_axi_gmem_WREADY,
	fib_63_m_axi_gmem_WVALID,
	fib_63_m_axi_gmem_WDATA,
	fib_63_m_axi_gmem_WSTRB,
	fib_63_m_axi_gmem_WLAST,
	fib_63_m_axi_gmem_WUSER,
	fib_63_m_axi_gmem_BREADY,
	fib_63_m_axi_gmem_BVALID,
	fib_63_m_axi_gmem_BID,
	fib_63_m_axi_gmem_BRESP,
	fib_63_m_axi_gmem_BUSER,
	fib_63_s_axi_control_ARREADY,
	fib_63_s_axi_control_ARVALID,
	fib_63_s_axi_control_ARADDR,
	fib_63_s_axi_control_RREADY,
	fib_63_s_axi_control_RVALID,
	fib_63_s_axi_control_RDATA,
	fib_63_s_axi_control_RRESP,
	fib_63_s_axi_control_AWREADY,
	fib_63_s_axi_control_AWVALID,
	fib_63_s_axi_control_AWADDR,
	fib_63_s_axi_control_WREADY,
	fib_63_s_axi_control_WVALID,
	fib_63_s_axi_control_WDATA,
	fib_63_s_axi_control_WSTRB,
	fib_63_s_axi_control_BREADY,
	fib_63_s_axi_control_BVALID,
	fib_63_s_axi_control_BRESP,
	fib_schedulerAXI_0_ARREADY,
	fib_schedulerAXI_0_ARVALID,
	fib_schedulerAXI_0_ARID,
	fib_schedulerAXI_0_ARADDR,
	fib_schedulerAXI_0_ARLEN,
	fib_schedulerAXI_0_ARSIZE,
	fib_schedulerAXI_0_ARBURST,
	fib_schedulerAXI_0_ARLOCK,
	fib_schedulerAXI_0_ARCACHE,
	fib_schedulerAXI_0_ARPROT,
	fib_schedulerAXI_0_ARQOS,
	fib_schedulerAXI_0_ARREGION,
	fib_schedulerAXI_0_RREADY,
	fib_schedulerAXI_0_RVALID,
	fib_schedulerAXI_0_RID,
	fib_schedulerAXI_0_RDATA,
	fib_schedulerAXI_0_RRESP,
	fib_schedulerAXI_0_RLAST,
	fib_schedulerAXI_0_AWREADY,
	fib_schedulerAXI_0_AWVALID,
	fib_schedulerAXI_0_AWID,
	fib_schedulerAXI_0_AWADDR,
	fib_schedulerAXI_0_AWLEN,
	fib_schedulerAXI_0_AWSIZE,
	fib_schedulerAXI_0_AWBURST,
	fib_schedulerAXI_0_AWLOCK,
	fib_schedulerAXI_0_AWCACHE,
	fib_schedulerAXI_0_AWPROT,
	fib_schedulerAXI_0_AWQOS,
	fib_schedulerAXI_0_AWREGION,
	fib_schedulerAXI_0_WREADY,
	fib_schedulerAXI_0_WVALID,
	fib_schedulerAXI_0_WDATA,
	fib_schedulerAXI_0_WSTRB,
	fib_schedulerAXI_0_WLAST,
	fib_schedulerAXI_0_BREADY,
	fib_schedulerAXI_0_BVALID,
	fib_schedulerAXI_0_BID,
	fib_schedulerAXI_0_BRESP,
	sum_0_m_axi_gmem_ARREADY,
	sum_0_m_axi_gmem_ARVALID,
	sum_0_m_axi_gmem_ARID,
	sum_0_m_axi_gmem_ARADDR,
	sum_0_m_axi_gmem_ARLEN,
	sum_0_m_axi_gmem_ARSIZE,
	sum_0_m_axi_gmem_ARBURST,
	sum_0_m_axi_gmem_ARLOCK,
	sum_0_m_axi_gmem_ARCACHE,
	sum_0_m_axi_gmem_ARPROT,
	sum_0_m_axi_gmem_ARQOS,
	sum_0_m_axi_gmem_ARREGION,
	sum_0_m_axi_gmem_ARUSER,
	sum_0_m_axi_gmem_RREADY,
	sum_0_m_axi_gmem_RVALID,
	sum_0_m_axi_gmem_RID,
	sum_0_m_axi_gmem_RDATA,
	sum_0_m_axi_gmem_RRESP,
	sum_0_m_axi_gmem_RLAST,
	sum_0_m_axi_gmem_RUSER,
	sum_0_m_axi_gmem_AWREADY,
	sum_0_m_axi_gmem_AWVALID,
	sum_0_m_axi_gmem_AWID,
	sum_0_m_axi_gmem_AWADDR,
	sum_0_m_axi_gmem_AWLEN,
	sum_0_m_axi_gmem_AWSIZE,
	sum_0_m_axi_gmem_AWBURST,
	sum_0_m_axi_gmem_AWLOCK,
	sum_0_m_axi_gmem_AWCACHE,
	sum_0_m_axi_gmem_AWPROT,
	sum_0_m_axi_gmem_AWQOS,
	sum_0_m_axi_gmem_AWREGION,
	sum_0_m_axi_gmem_AWUSER,
	sum_0_m_axi_gmem_WREADY,
	sum_0_m_axi_gmem_WVALID,
	sum_0_m_axi_gmem_WDATA,
	sum_0_m_axi_gmem_WSTRB,
	sum_0_m_axi_gmem_WLAST,
	sum_0_m_axi_gmem_WUSER,
	sum_0_m_axi_gmem_BREADY,
	sum_0_m_axi_gmem_BVALID,
	sum_0_m_axi_gmem_BID,
	sum_0_m_axi_gmem_BRESP,
	sum_0_m_axi_gmem_BUSER,
	sum_0_s_axi_control_ARREADY,
	sum_0_s_axi_control_ARVALID,
	sum_0_s_axi_control_ARADDR,
	sum_0_s_axi_control_RREADY,
	sum_0_s_axi_control_RVALID,
	sum_0_s_axi_control_RDATA,
	sum_0_s_axi_control_RRESP,
	sum_0_s_axi_control_AWREADY,
	sum_0_s_axi_control_AWVALID,
	sum_0_s_axi_control_AWADDR,
	sum_0_s_axi_control_WREADY,
	sum_0_s_axi_control_WVALID,
	sum_0_s_axi_control_WDATA,
	sum_0_s_axi_control_WSTRB,
	sum_0_s_axi_control_BREADY,
	sum_0_s_axi_control_BVALID,
	sum_0_s_axi_control_BRESP,
	sum_1_m_axi_gmem_ARREADY,
	sum_1_m_axi_gmem_ARVALID,
	sum_1_m_axi_gmem_ARID,
	sum_1_m_axi_gmem_ARADDR,
	sum_1_m_axi_gmem_ARLEN,
	sum_1_m_axi_gmem_ARSIZE,
	sum_1_m_axi_gmem_ARBURST,
	sum_1_m_axi_gmem_ARLOCK,
	sum_1_m_axi_gmem_ARCACHE,
	sum_1_m_axi_gmem_ARPROT,
	sum_1_m_axi_gmem_ARQOS,
	sum_1_m_axi_gmem_ARREGION,
	sum_1_m_axi_gmem_ARUSER,
	sum_1_m_axi_gmem_RREADY,
	sum_1_m_axi_gmem_RVALID,
	sum_1_m_axi_gmem_RID,
	sum_1_m_axi_gmem_RDATA,
	sum_1_m_axi_gmem_RRESP,
	sum_1_m_axi_gmem_RLAST,
	sum_1_m_axi_gmem_RUSER,
	sum_1_m_axi_gmem_AWREADY,
	sum_1_m_axi_gmem_AWVALID,
	sum_1_m_axi_gmem_AWID,
	sum_1_m_axi_gmem_AWADDR,
	sum_1_m_axi_gmem_AWLEN,
	sum_1_m_axi_gmem_AWSIZE,
	sum_1_m_axi_gmem_AWBURST,
	sum_1_m_axi_gmem_AWLOCK,
	sum_1_m_axi_gmem_AWCACHE,
	sum_1_m_axi_gmem_AWPROT,
	sum_1_m_axi_gmem_AWQOS,
	sum_1_m_axi_gmem_AWREGION,
	sum_1_m_axi_gmem_AWUSER,
	sum_1_m_axi_gmem_WREADY,
	sum_1_m_axi_gmem_WVALID,
	sum_1_m_axi_gmem_WDATA,
	sum_1_m_axi_gmem_WSTRB,
	sum_1_m_axi_gmem_WLAST,
	sum_1_m_axi_gmem_WUSER,
	sum_1_m_axi_gmem_BREADY,
	sum_1_m_axi_gmem_BVALID,
	sum_1_m_axi_gmem_BID,
	sum_1_m_axi_gmem_BRESP,
	sum_1_m_axi_gmem_BUSER,
	sum_1_s_axi_control_ARREADY,
	sum_1_s_axi_control_ARVALID,
	sum_1_s_axi_control_ARADDR,
	sum_1_s_axi_control_RREADY,
	sum_1_s_axi_control_RVALID,
	sum_1_s_axi_control_RDATA,
	sum_1_s_axi_control_RRESP,
	sum_1_s_axi_control_AWREADY,
	sum_1_s_axi_control_AWVALID,
	sum_1_s_axi_control_AWADDR,
	sum_1_s_axi_control_WREADY,
	sum_1_s_axi_control_WVALID,
	sum_1_s_axi_control_WDATA,
	sum_1_s_axi_control_WSTRB,
	sum_1_s_axi_control_BREADY,
	sum_1_s_axi_control_BVALID,
	sum_1_s_axi_control_BRESP,
	sum_2_m_axi_gmem_ARREADY,
	sum_2_m_axi_gmem_ARVALID,
	sum_2_m_axi_gmem_ARID,
	sum_2_m_axi_gmem_ARADDR,
	sum_2_m_axi_gmem_ARLEN,
	sum_2_m_axi_gmem_ARSIZE,
	sum_2_m_axi_gmem_ARBURST,
	sum_2_m_axi_gmem_ARLOCK,
	sum_2_m_axi_gmem_ARCACHE,
	sum_2_m_axi_gmem_ARPROT,
	sum_2_m_axi_gmem_ARQOS,
	sum_2_m_axi_gmem_ARREGION,
	sum_2_m_axi_gmem_ARUSER,
	sum_2_m_axi_gmem_RREADY,
	sum_2_m_axi_gmem_RVALID,
	sum_2_m_axi_gmem_RID,
	sum_2_m_axi_gmem_RDATA,
	sum_2_m_axi_gmem_RRESP,
	sum_2_m_axi_gmem_RLAST,
	sum_2_m_axi_gmem_RUSER,
	sum_2_m_axi_gmem_AWREADY,
	sum_2_m_axi_gmem_AWVALID,
	sum_2_m_axi_gmem_AWID,
	sum_2_m_axi_gmem_AWADDR,
	sum_2_m_axi_gmem_AWLEN,
	sum_2_m_axi_gmem_AWSIZE,
	sum_2_m_axi_gmem_AWBURST,
	sum_2_m_axi_gmem_AWLOCK,
	sum_2_m_axi_gmem_AWCACHE,
	sum_2_m_axi_gmem_AWPROT,
	sum_2_m_axi_gmem_AWQOS,
	sum_2_m_axi_gmem_AWREGION,
	sum_2_m_axi_gmem_AWUSER,
	sum_2_m_axi_gmem_WREADY,
	sum_2_m_axi_gmem_WVALID,
	sum_2_m_axi_gmem_WDATA,
	sum_2_m_axi_gmem_WSTRB,
	sum_2_m_axi_gmem_WLAST,
	sum_2_m_axi_gmem_WUSER,
	sum_2_m_axi_gmem_BREADY,
	sum_2_m_axi_gmem_BVALID,
	sum_2_m_axi_gmem_BID,
	sum_2_m_axi_gmem_BRESP,
	sum_2_m_axi_gmem_BUSER,
	sum_2_s_axi_control_ARREADY,
	sum_2_s_axi_control_ARVALID,
	sum_2_s_axi_control_ARADDR,
	sum_2_s_axi_control_RREADY,
	sum_2_s_axi_control_RVALID,
	sum_2_s_axi_control_RDATA,
	sum_2_s_axi_control_RRESP,
	sum_2_s_axi_control_AWREADY,
	sum_2_s_axi_control_AWVALID,
	sum_2_s_axi_control_AWADDR,
	sum_2_s_axi_control_WREADY,
	sum_2_s_axi_control_WVALID,
	sum_2_s_axi_control_WDATA,
	sum_2_s_axi_control_WSTRB,
	sum_2_s_axi_control_BREADY,
	sum_2_s_axi_control_BVALID,
	sum_2_s_axi_control_BRESP,
	sum_3_m_axi_gmem_ARREADY,
	sum_3_m_axi_gmem_ARVALID,
	sum_3_m_axi_gmem_ARID,
	sum_3_m_axi_gmem_ARADDR,
	sum_3_m_axi_gmem_ARLEN,
	sum_3_m_axi_gmem_ARSIZE,
	sum_3_m_axi_gmem_ARBURST,
	sum_3_m_axi_gmem_ARLOCK,
	sum_3_m_axi_gmem_ARCACHE,
	sum_3_m_axi_gmem_ARPROT,
	sum_3_m_axi_gmem_ARQOS,
	sum_3_m_axi_gmem_ARREGION,
	sum_3_m_axi_gmem_ARUSER,
	sum_3_m_axi_gmem_RREADY,
	sum_3_m_axi_gmem_RVALID,
	sum_3_m_axi_gmem_RID,
	sum_3_m_axi_gmem_RDATA,
	sum_3_m_axi_gmem_RRESP,
	sum_3_m_axi_gmem_RLAST,
	sum_3_m_axi_gmem_RUSER,
	sum_3_m_axi_gmem_AWREADY,
	sum_3_m_axi_gmem_AWVALID,
	sum_3_m_axi_gmem_AWID,
	sum_3_m_axi_gmem_AWADDR,
	sum_3_m_axi_gmem_AWLEN,
	sum_3_m_axi_gmem_AWSIZE,
	sum_3_m_axi_gmem_AWBURST,
	sum_3_m_axi_gmem_AWLOCK,
	sum_3_m_axi_gmem_AWCACHE,
	sum_3_m_axi_gmem_AWPROT,
	sum_3_m_axi_gmem_AWQOS,
	sum_3_m_axi_gmem_AWREGION,
	sum_3_m_axi_gmem_AWUSER,
	sum_3_m_axi_gmem_WREADY,
	sum_3_m_axi_gmem_WVALID,
	sum_3_m_axi_gmem_WDATA,
	sum_3_m_axi_gmem_WSTRB,
	sum_3_m_axi_gmem_WLAST,
	sum_3_m_axi_gmem_WUSER,
	sum_3_m_axi_gmem_BREADY,
	sum_3_m_axi_gmem_BVALID,
	sum_3_m_axi_gmem_BID,
	sum_3_m_axi_gmem_BRESP,
	sum_3_m_axi_gmem_BUSER,
	sum_3_s_axi_control_ARREADY,
	sum_3_s_axi_control_ARVALID,
	sum_3_s_axi_control_ARADDR,
	sum_3_s_axi_control_RREADY,
	sum_3_s_axi_control_RVALID,
	sum_3_s_axi_control_RDATA,
	sum_3_s_axi_control_RRESP,
	sum_3_s_axi_control_AWREADY,
	sum_3_s_axi_control_AWVALID,
	sum_3_s_axi_control_AWADDR,
	sum_3_s_axi_control_WREADY,
	sum_3_s_axi_control_WVALID,
	sum_3_s_axi_control_WDATA,
	sum_3_s_axi_control_WSTRB,
	sum_3_s_axi_control_BREADY,
	sum_3_s_axi_control_BVALID,
	sum_3_s_axi_control_BRESP,
	sum_4_m_axi_gmem_ARREADY,
	sum_4_m_axi_gmem_ARVALID,
	sum_4_m_axi_gmem_ARID,
	sum_4_m_axi_gmem_ARADDR,
	sum_4_m_axi_gmem_ARLEN,
	sum_4_m_axi_gmem_ARSIZE,
	sum_4_m_axi_gmem_ARBURST,
	sum_4_m_axi_gmem_ARLOCK,
	sum_4_m_axi_gmem_ARCACHE,
	sum_4_m_axi_gmem_ARPROT,
	sum_4_m_axi_gmem_ARQOS,
	sum_4_m_axi_gmem_ARREGION,
	sum_4_m_axi_gmem_ARUSER,
	sum_4_m_axi_gmem_RREADY,
	sum_4_m_axi_gmem_RVALID,
	sum_4_m_axi_gmem_RID,
	sum_4_m_axi_gmem_RDATA,
	sum_4_m_axi_gmem_RRESP,
	sum_4_m_axi_gmem_RLAST,
	sum_4_m_axi_gmem_RUSER,
	sum_4_m_axi_gmem_AWREADY,
	sum_4_m_axi_gmem_AWVALID,
	sum_4_m_axi_gmem_AWID,
	sum_4_m_axi_gmem_AWADDR,
	sum_4_m_axi_gmem_AWLEN,
	sum_4_m_axi_gmem_AWSIZE,
	sum_4_m_axi_gmem_AWBURST,
	sum_4_m_axi_gmem_AWLOCK,
	sum_4_m_axi_gmem_AWCACHE,
	sum_4_m_axi_gmem_AWPROT,
	sum_4_m_axi_gmem_AWQOS,
	sum_4_m_axi_gmem_AWREGION,
	sum_4_m_axi_gmem_AWUSER,
	sum_4_m_axi_gmem_WREADY,
	sum_4_m_axi_gmem_WVALID,
	sum_4_m_axi_gmem_WDATA,
	sum_4_m_axi_gmem_WSTRB,
	sum_4_m_axi_gmem_WLAST,
	sum_4_m_axi_gmem_WUSER,
	sum_4_m_axi_gmem_BREADY,
	sum_4_m_axi_gmem_BVALID,
	sum_4_m_axi_gmem_BID,
	sum_4_m_axi_gmem_BRESP,
	sum_4_m_axi_gmem_BUSER,
	sum_4_s_axi_control_ARREADY,
	sum_4_s_axi_control_ARVALID,
	sum_4_s_axi_control_ARADDR,
	sum_4_s_axi_control_RREADY,
	sum_4_s_axi_control_RVALID,
	sum_4_s_axi_control_RDATA,
	sum_4_s_axi_control_RRESP,
	sum_4_s_axi_control_AWREADY,
	sum_4_s_axi_control_AWVALID,
	sum_4_s_axi_control_AWADDR,
	sum_4_s_axi_control_WREADY,
	sum_4_s_axi_control_WVALID,
	sum_4_s_axi_control_WDATA,
	sum_4_s_axi_control_WSTRB,
	sum_4_s_axi_control_BREADY,
	sum_4_s_axi_control_BVALID,
	sum_4_s_axi_control_BRESP,
	sum_5_m_axi_gmem_ARREADY,
	sum_5_m_axi_gmem_ARVALID,
	sum_5_m_axi_gmem_ARID,
	sum_5_m_axi_gmem_ARADDR,
	sum_5_m_axi_gmem_ARLEN,
	sum_5_m_axi_gmem_ARSIZE,
	sum_5_m_axi_gmem_ARBURST,
	sum_5_m_axi_gmem_ARLOCK,
	sum_5_m_axi_gmem_ARCACHE,
	sum_5_m_axi_gmem_ARPROT,
	sum_5_m_axi_gmem_ARQOS,
	sum_5_m_axi_gmem_ARREGION,
	sum_5_m_axi_gmem_ARUSER,
	sum_5_m_axi_gmem_RREADY,
	sum_5_m_axi_gmem_RVALID,
	sum_5_m_axi_gmem_RID,
	sum_5_m_axi_gmem_RDATA,
	sum_5_m_axi_gmem_RRESP,
	sum_5_m_axi_gmem_RLAST,
	sum_5_m_axi_gmem_RUSER,
	sum_5_m_axi_gmem_AWREADY,
	sum_5_m_axi_gmem_AWVALID,
	sum_5_m_axi_gmem_AWID,
	sum_5_m_axi_gmem_AWADDR,
	sum_5_m_axi_gmem_AWLEN,
	sum_5_m_axi_gmem_AWSIZE,
	sum_5_m_axi_gmem_AWBURST,
	sum_5_m_axi_gmem_AWLOCK,
	sum_5_m_axi_gmem_AWCACHE,
	sum_5_m_axi_gmem_AWPROT,
	sum_5_m_axi_gmem_AWQOS,
	sum_5_m_axi_gmem_AWREGION,
	sum_5_m_axi_gmem_AWUSER,
	sum_5_m_axi_gmem_WREADY,
	sum_5_m_axi_gmem_WVALID,
	sum_5_m_axi_gmem_WDATA,
	sum_5_m_axi_gmem_WSTRB,
	sum_5_m_axi_gmem_WLAST,
	sum_5_m_axi_gmem_WUSER,
	sum_5_m_axi_gmem_BREADY,
	sum_5_m_axi_gmem_BVALID,
	sum_5_m_axi_gmem_BID,
	sum_5_m_axi_gmem_BRESP,
	sum_5_m_axi_gmem_BUSER,
	sum_5_s_axi_control_ARREADY,
	sum_5_s_axi_control_ARVALID,
	sum_5_s_axi_control_ARADDR,
	sum_5_s_axi_control_RREADY,
	sum_5_s_axi_control_RVALID,
	sum_5_s_axi_control_RDATA,
	sum_5_s_axi_control_RRESP,
	sum_5_s_axi_control_AWREADY,
	sum_5_s_axi_control_AWVALID,
	sum_5_s_axi_control_AWADDR,
	sum_5_s_axi_control_WREADY,
	sum_5_s_axi_control_WVALID,
	sum_5_s_axi_control_WDATA,
	sum_5_s_axi_control_WSTRB,
	sum_5_s_axi_control_BREADY,
	sum_5_s_axi_control_BVALID,
	sum_5_s_axi_control_BRESP,
	sum_6_m_axi_gmem_ARREADY,
	sum_6_m_axi_gmem_ARVALID,
	sum_6_m_axi_gmem_ARID,
	sum_6_m_axi_gmem_ARADDR,
	sum_6_m_axi_gmem_ARLEN,
	sum_6_m_axi_gmem_ARSIZE,
	sum_6_m_axi_gmem_ARBURST,
	sum_6_m_axi_gmem_ARLOCK,
	sum_6_m_axi_gmem_ARCACHE,
	sum_6_m_axi_gmem_ARPROT,
	sum_6_m_axi_gmem_ARQOS,
	sum_6_m_axi_gmem_ARREGION,
	sum_6_m_axi_gmem_ARUSER,
	sum_6_m_axi_gmem_RREADY,
	sum_6_m_axi_gmem_RVALID,
	sum_6_m_axi_gmem_RID,
	sum_6_m_axi_gmem_RDATA,
	sum_6_m_axi_gmem_RRESP,
	sum_6_m_axi_gmem_RLAST,
	sum_6_m_axi_gmem_RUSER,
	sum_6_m_axi_gmem_AWREADY,
	sum_6_m_axi_gmem_AWVALID,
	sum_6_m_axi_gmem_AWID,
	sum_6_m_axi_gmem_AWADDR,
	sum_6_m_axi_gmem_AWLEN,
	sum_6_m_axi_gmem_AWSIZE,
	sum_6_m_axi_gmem_AWBURST,
	sum_6_m_axi_gmem_AWLOCK,
	sum_6_m_axi_gmem_AWCACHE,
	sum_6_m_axi_gmem_AWPROT,
	sum_6_m_axi_gmem_AWQOS,
	sum_6_m_axi_gmem_AWREGION,
	sum_6_m_axi_gmem_AWUSER,
	sum_6_m_axi_gmem_WREADY,
	sum_6_m_axi_gmem_WVALID,
	sum_6_m_axi_gmem_WDATA,
	sum_6_m_axi_gmem_WSTRB,
	sum_6_m_axi_gmem_WLAST,
	sum_6_m_axi_gmem_WUSER,
	sum_6_m_axi_gmem_BREADY,
	sum_6_m_axi_gmem_BVALID,
	sum_6_m_axi_gmem_BID,
	sum_6_m_axi_gmem_BRESP,
	sum_6_m_axi_gmem_BUSER,
	sum_6_s_axi_control_ARREADY,
	sum_6_s_axi_control_ARVALID,
	sum_6_s_axi_control_ARADDR,
	sum_6_s_axi_control_RREADY,
	sum_6_s_axi_control_RVALID,
	sum_6_s_axi_control_RDATA,
	sum_6_s_axi_control_RRESP,
	sum_6_s_axi_control_AWREADY,
	sum_6_s_axi_control_AWVALID,
	sum_6_s_axi_control_AWADDR,
	sum_6_s_axi_control_WREADY,
	sum_6_s_axi_control_WVALID,
	sum_6_s_axi_control_WDATA,
	sum_6_s_axi_control_WSTRB,
	sum_6_s_axi_control_BREADY,
	sum_6_s_axi_control_BVALID,
	sum_6_s_axi_control_BRESP,
	sum_7_m_axi_gmem_ARREADY,
	sum_7_m_axi_gmem_ARVALID,
	sum_7_m_axi_gmem_ARID,
	sum_7_m_axi_gmem_ARADDR,
	sum_7_m_axi_gmem_ARLEN,
	sum_7_m_axi_gmem_ARSIZE,
	sum_7_m_axi_gmem_ARBURST,
	sum_7_m_axi_gmem_ARLOCK,
	sum_7_m_axi_gmem_ARCACHE,
	sum_7_m_axi_gmem_ARPROT,
	sum_7_m_axi_gmem_ARQOS,
	sum_7_m_axi_gmem_ARREGION,
	sum_7_m_axi_gmem_ARUSER,
	sum_7_m_axi_gmem_RREADY,
	sum_7_m_axi_gmem_RVALID,
	sum_7_m_axi_gmem_RID,
	sum_7_m_axi_gmem_RDATA,
	sum_7_m_axi_gmem_RRESP,
	sum_7_m_axi_gmem_RLAST,
	sum_7_m_axi_gmem_RUSER,
	sum_7_m_axi_gmem_AWREADY,
	sum_7_m_axi_gmem_AWVALID,
	sum_7_m_axi_gmem_AWID,
	sum_7_m_axi_gmem_AWADDR,
	sum_7_m_axi_gmem_AWLEN,
	sum_7_m_axi_gmem_AWSIZE,
	sum_7_m_axi_gmem_AWBURST,
	sum_7_m_axi_gmem_AWLOCK,
	sum_7_m_axi_gmem_AWCACHE,
	sum_7_m_axi_gmem_AWPROT,
	sum_7_m_axi_gmem_AWQOS,
	sum_7_m_axi_gmem_AWREGION,
	sum_7_m_axi_gmem_AWUSER,
	sum_7_m_axi_gmem_WREADY,
	sum_7_m_axi_gmem_WVALID,
	sum_7_m_axi_gmem_WDATA,
	sum_7_m_axi_gmem_WSTRB,
	sum_7_m_axi_gmem_WLAST,
	sum_7_m_axi_gmem_WUSER,
	sum_7_m_axi_gmem_BREADY,
	sum_7_m_axi_gmem_BVALID,
	sum_7_m_axi_gmem_BID,
	sum_7_m_axi_gmem_BRESP,
	sum_7_m_axi_gmem_BUSER,
	sum_7_s_axi_control_ARREADY,
	sum_7_s_axi_control_ARVALID,
	sum_7_s_axi_control_ARADDR,
	sum_7_s_axi_control_RREADY,
	sum_7_s_axi_control_RVALID,
	sum_7_s_axi_control_RDATA,
	sum_7_s_axi_control_RRESP,
	sum_7_s_axi_control_AWREADY,
	sum_7_s_axi_control_AWVALID,
	sum_7_s_axi_control_AWADDR,
	sum_7_s_axi_control_WREADY,
	sum_7_s_axi_control_WVALID,
	sum_7_s_axi_control_WDATA,
	sum_7_s_axi_control_WSTRB,
	sum_7_s_axi_control_BREADY,
	sum_7_s_axi_control_BVALID,
	sum_7_s_axi_control_BRESP,
	sum_8_m_axi_gmem_ARREADY,
	sum_8_m_axi_gmem_ARVALID,
	sum_8_m_axi_gmem_ARID,
	sum_8_m_axi_gmem_ARADDR,
	sum_8_m_axi_gmem_ARLEN,
	sum_8_m_axi_gmem_ARSIZE,
	sum_8_m_axi_gmem_ARBURST,
	sum_8_m_axi_gmem_ARLOCK,
	sum_8_m_axi_gmem_ARCACHE,
	sum_8_m_axi_gmem_ARPROT,
	sum_8_m_axi_gmem_ARQOS,
	sum_8_m_axi_gmem_ARREGION,
	sum_8_m_axi_gmem_ARUSER,
	sum_8_m_axi_gmem_RREADY,
	sum_8_m_axi_gmem_RVALID,
	sum_8_m_axi_gmem_RID,
	sum_8_m_axi_gmem_RDATA,
	sum_8_m_axi_gmem_RRESP,
	sum_8_m_axi_gmem_RLAST,
	sum_8_m_axi_gmem_RUSER,
	sum_8_m_axi_gmem_AWREADY,
	sum_8_m_axi_gmem_AWVALID,
	sum_8_m_axi_gmem_AWID,
	sum_8_m_axi_gmem_AWADDR,
	sum_8_m_axi_gmem_AWLEN,
	sum_8_m_axi_gmem_AWSIZE,
	sum_8_m_axi_gmem_AWBURST,
	sum_8_m_axi_gmem_AWLOCK,
	sum_8_m_axi_gmem_AWCACHE,
	sum_8_m_axi_gmem_AWPROT,
	sum_8_m_axi_gmem_AWQOS,
	sum_8_m_axi_gmem_AWREGION,
	sum_8_m_axi_gmem_AWUSER,
	sum_8_m_axi_gmem_WREADY,
	sum_8_m_axi_gmem_WVALID,
	sum_8_m_axi_gmem_WDATA,
	sum_8_m_axi_gmem_WSTRB,
	sum_8_m_axi_gmem_WLAST,
	sum_8_m_axi_gmem_WUSER,
	sum_8_m_axi_gmem_BREADY,
	sum_8_m_axi_gmem_BVALID,
	sum_8_m_axi_gmem_BID,
	sum_8_m_axi_gmem_BRESP,
	sum_8_m_axi_gmem_BUSER,
	sum_8_s_axi_control_ARREADY,
	sum_8_s_axi_control_ARVALID,
	sum_8_s_axi_control_ARADDR,
	sum_8_s_axi_control_RREADY,
	sum_8_s_axi_control_RVALID,
	sum_8_s_axi_control_RDATA,
	sum_8_s_axi_control_RRESP,
	sum_8_s_axi_control_AWREADY,
	sum_8_s_axi_control_AWVALID,
	sum_8_s_axi_control_AWADDR,
	sum_8_s_axi_control_WREADY,
	sum_8_s_axi_control_WVALID,
	sum_8_s_axi_control_WDATA,
	sum_8_s_axi_control_WSTRB,
	sum_8_s_axi_control_BREADY,
	sum_8_s_axi_control_BVALID,
	sum_8_s_axi_control_BRESP,
	sum_9_m_axi_gmem_ARREADY,
	sum_9_m_axi_gmem_ARVALID,
	sum_9_m_axi_gmem_ARID,
	sum_9_m_axi_gmem_ARADDR,
	sum_9_m_axi_gmem_ARLEN,
	sum_9_m_axi_gmem_ARSIZE,
	sum_9_m_axi_gmem_ARBURST,
	sum_9_m_axi_gmem_ARLOCK,
	sum_9_m_axi_gmem_ARCACHE,
	sum_9_m_axi_gmem_ARPROT,
	sum_9_m_axi_gmem_ARQOS,
	sum_9_m_axi_gmem_ARREGION,
	sum_9_m_axi_gmem_ARUSER,
	sum_9_m_axi_gmem_RREADY,
	sum_9_m_axi_gmem_RVALID,
	sum_9_m_axi_gmem_RID,
	sum_9_m_axi_gmem_RDATA,
	sum_9_m_axi_gmem_RRESP,
	sum_9_m_axi_gmem_RLAST,
	sum_9_m_axi_gmem_RUSER,
	sum_9_m_axi_gmem_AWREADY,
	sum_9_m_axi_gmem_AWVALID,
	sum_9_m_axi_gmem_AWID,
	sum_9_m_axi_gmem_AWADDR,
	sum_9_m_axi_gmem_AWLEN,
	sum_9_m_axi_gmem_AWSIZE,
	sum_9_m_axi_gmem_AWBURST,
	sum_9_m_axi_gmem_AWLOCK,
	sum_9_m_axi_gmem_AWCACHE,
	sum_9_m_axi_gmem_AWPROT,
	sum_9_m_axi_gmem_AWQOS,
	sum_9_m_axi_gmem_AWREGION,
	sum_9_m_axi_gmem_AWUSER,
	sum_9_m_axi_gmem_WREADY,
	sum_9_m_axi_gmem_WVALID,
	sum_9_m_axi_gmem_WDATA,
	sum_9_m_axi_gmem_WSTRB,
	sum_9_m_axi_gmem_WLAST,
	sum_9_m_axi_gmem_WUSER,
	sum_9_m_axi_gmem_BREADY,
	sum_9_m_axi_gmem_BVALID,
	sum_9_m_axi_gmem_BID,
	sum_9_m_axi_gmem_BRESP,
	sum_9_m_axi_gmem_BUSER,
	sum_9_s_axi_control_ARREADY,
	sum_9_s_axi_control_ARVALID,
	sum_9_s_axi_control_ARADDR,
	sum_9_s_axi_control_RREADY,
	sum_9_s_axi_control_RVALID,
	sum_9_s_axi_control_RDATA,
	sum_9_s_axi_control_RRESP,
	sum_9_s_axi_control_AWREADY,
	sum_9_s_axi_control_AWVALID,
	sum_9_s_axi_control_AWADDR,
	sum_9_s_axi_control_WREADY,
	sum_9_s_axi_control_WVALID,
	sum_9_s_axi_control_WDATA,
	sum_9_s_axi_control_WSTRB,
	sum_9_s_axi_control_BREADY,
	sum_9_s_axi_control_BVALID,
	sum_9_s_axi_control_BRESP,
	sum_10_m_axi_gmem_ARREADY,
	sum_10_m_axi_gmem_ARVALID,
	sum_10_m_axi_gmem_ARID,
	sum_10_m_axi_gmem_ARADDR,
	sum_10_m_axi_gmem_ARLEN,
	sum_10_m_axi_gmem_ARSIZE,
	sum_10_m_axi_gmem_ARBURST,
	sum_10_m_axi_gmem_ARLOCK,
	sum_10_m_axi_gmem_ARCACHE,
	sum_10_m_axi_gmem_ARPROT,
	sum_10_m_axi_gmem_ARQOS,
	sum_10_m_axi_gmem_ARREGION,
	sum_10_m_axi_gmem_ARUSER,
	sum_10_m_axi_gmem_RREADY,
	sum_10_m_axi_gmem_RVALID,
	sum_10_m_axi_gmem_RID,
	sum_10_m_axi_gmem_RDATA,
	sum_10_m_axi_gmem_RRESP,
	sum_10_m_axi_gmem_RLAST,
	sum_10_m_axi_gmem_RUSER,
	sum_10_m_axi_gmem_AWREADY,
	sum_10_m_axi_gmem_AWVALID,
	sum_10_m_axi_gmem_AWID,
	sum_10_m_axi_gmem_AWADDR,
	sum_10_m_axi_gmem_AWLEN,
	sum_10_m_axi_gmem_AWSIZE,
	sum_10_m_axi_gmem_AWBURST,
	sum_10_m_axi_gmem_AWLOCK,
	sum_10_m_axi_gmem_AWCACHE,
	sum_10_m_axi_gmem_AWPROT,
	sum_10_m_axi_gmem_AWQOS,
	sum_10_m_axi_gmem_AWREGION,
	sum_10_m_axi_gmem_AWUSER,
	sum_10_m_axi_gmem_WREADY,
	sum_10_m_axi_gmem_WVALID,
	sum_10_m_axi_gmem_WDATA,
	sum_10_m_axi_gmem_WSTRB,
	sum_10_m_axi_gmem_WLAST,
	sum_10_m_axi_gmem_WUSER,
	sum_10_m_axi_gmem_BREADY,
	sum_10_m_axi_gmem_BVALID,
	sum_10_m_axi_gmem_BID,
	sum_10_m_axi_gmem_BRESP,
	sum_10_m_axi_gmem_BUSER,
	sum_10_s_axi_control_ARREADY,
	sum_10_s_axi_control_ARVALID,
	sum_10_s_axi_control_ARADDR,
	sum_10_s_axi_control_RREADY,
	sum_10_s_axi_control_RVALID,
	sum_10_s_axi_control_RDATA,
	sum_10_s_axi_control_RRESP,
	sum_10_s_axi_control_AWREADY,
	sum_10_s_axi_control_AWVALID,
	sum_10_s_axi_control_AWADDR,
	sum_10_s_axi_control_WREADY,
	sum_10_s_axi_control_WVALID,
	sum_10_s_axi_control_WDATA,
	sum_10_s_axi_control_WSTRB,
	sum_10_s_axi_control_BREADY,
	sum_10_s_axi_control_BVALID,
	sum_10_s_axi_control_BRESP,
	sum_11_m_axi_gmem_ARREADY,
	sum_11_m_axi_gmem_ARVALID,
	sum_11_m_axi_gmem_ARID,
	sum_11_m_axi_gmem_ARADDR,
	sum_11_m_axi_gmem_ARLEN,
	sum_11_m_axi_gmem_ARSIZE,
	sum_11_m_axi_gmem_ARBURST,
	sum_11_m_axi_gmem_ARLOCK,
	sum_11_m_axi_gmem_ARCACHE,
	sum_11_m_axi_gmem_ARPROT,
	sum_11_m_axi_gmem_ARQOS,
	sum_11_m_axi_gmem_ARREGION,
	sum_11_m_axi_gmem_ARUSER,
	sum_11_m_axi_gmem_RREADY,
	sum_11_m_axi_gmem_RVALID,
	sum_11_m_axi_gmem_RID,
	sum_11_m_axi_gmem_RDATA,
	sum_11_m_axi_gmem_RRESP,
	sum_11_m_axi_gmem_RLAST,
	sum_11_m_axi_gmem_RUSER,
	sum_11_m_axi_gmem_AWREADY,
	sum_11_m_axi_gmem_AWVALID,
	sum_11_m_axi_gmem_AWID,
	sum_11_m_axi_gmem_AWADDR,
	sum_11_m_axi_gmem_AWLEN,
	sum_11_m_axi_gmem_AWSIZE,
	sum_11_m_axi_gmem_AWBURST,
	sum_11_m_axi_gmem_AWLOCK,
	sum_11_m_axi_gmem_AWCACHE,
	sum_11_m_axi_gmem_AWPROT,
	sum_11_m_axi_gmem_AWQOS,
	sum_11_m_axi_gmem_AWREGION,
	sum_11_m_axi_gmem_AWUSER,
	sum_11_m_axi_gmem_WREADY,
	sum_11_m_axi_gmem_WVALID,
	sum_11_m_axi_gmem_WDATA,
	sum_11_m_axi_gmem_WSTRB,
	sum_11_m_axi_gmem_WLAST,
	sum_11_m_axi_gmem_WUSER,
	sum_11_m_axi_gmem_BREADY,
	sum_11_m_axi_gmem_BVALID,
	sum_11_m_axi_gmem_BID,
	sum_11_m_axi_gmem_BRESP,
	sum_11_m_axi_gmem_BUSER,
	sum_11_s_axi_control_ARREADY,
	sum_11_s_axi_control_ARVALID,
	sum_11_s_axi_control_ARADDR,
	sum_11_s_axi_control_RREADY,
	sum_11_s_axi_control_RVALID,
	sum_11_s_axi_control_RDATA,
	sum_11_s_axi_control_RRESP,
	sum_11_s_axi_control_AWREADY,
	sum_11_s_axi_control_AWVALID,
	sum_11_s_axi_control_AWADDR,
	sum_11_s_axi_control_WREADY,
	sum_11_s_axi_control_WVALID,
	sum_11_s_axi_control_WDATA,
	sum_11_s_axi_control_WSTRB,
	sum_11_s_axi_control_BREADY,
	sum_11_s_axi_control_BVALID,
	sum_11_s_axi_control_BRESP,
	sum_12_m_axi_gmem_ARREADY,
	sum_12_m_axi_gmem_ARVALID,
	sum_12_m_axi_gmem_ARID,
	sum_12_m_axi_gmem_ARADDR,
	sum_12_m_axi_gmem_ARLEN,
	sum_12_m_axi_gmem_ARSIZE,
	sum_12_m_axi_gmem_ARBURST,
	sum_12_m_axi_gmem_ARLOCK,
	sum_12_m_axi_gmem_ARCACHE,
	sum_12_m_axi_gmem_ARPROT,
	sum_12_m_axi_gmem_ARQOS,
	sum_12_m_axi_gmem_ARREGION,
	sum_12_m_axi_gmem_ARUSER,
	sum_12_m_axi_gmem_RREADY,
	sum_12_m_axi_gmem_RVALID,
	sum_12_m_axi_gmem_RID,
	sum_12_m_axi_gmem_RDATA,
	sum_12_m_axi_gmem_RRESP,
	sum_12_m_axi_gmem_RLAST,
	sum_12_m_axi_gmem_RUSER,
	sum_12_m_axi_gmem_AWREADY,
	sum_12_m_axi_gmem_AWVALID,
	sum_12_m_axi_gmem_AWID,
	sum_12_m_axi_gmem_AWADDR,
	sum_12_m_axi_gmem_AWLEN,
	sum_12_m_axi_gmem_AWSIZE,
	sum_12_m_axi_gmem_AWBURST,
	sum_12_m_axi_gmem_AWLOCK,
	sum_12_m_axi_gmem_AWCACHE,
	sum_12_m_axi_gmem_AWPROT,
	sum_12_m_axi_gmem_AWQOS,
	sum_12_m_axi_gmem_AWREGION,
	sum_12_m_axi_gmem_AWUSER,
	sum_12_m_axi_gmem_WREADY,
	sum_12_m_axi_gmem_WVALID,
	sum_12_m_axi_gmem_WDATA,
	sum_12_m_axi_gmem_WSTRB,
	sum_12_m_axi_gmem_WLAST,
	sum_12_m_axi_gmem_WUSER,
	sum_12_m_axi_gmem_BREADY,
	sum_12_m_axi_gmem_BVALID,
	sum_12_m_axi_gmem_BID,
	sum_12_m_axi_gmem_BRESP,
	sum_12_m_axi_gmem_BUSER,
	sum_12_s_axi_control_ARREADY,
	sum_12_s_axi_control_ARVALID,
	sum_12_s_axi_control_ARADDR,
	sum_12_s_axi_control_RREADY,
	sum_12_s_axi_control_RVALID,
	sum_12_s_axi_control_RDATA,
	sum_12_s_axi_control_RRESP,
	sum_12_s_axi_control_AWREADY,
	sum_12_s_axi_control_AWVALID,
	sum_12_s_axi_control_AWADDR,
	sum_12_s_axi_control_WREADY,
	sum_12_s_axi_control_WVALID,
	sum_12_s_axi_control_WDATA,
	sum_12_s_axi_control_WSTRB,
	sum_12_s_axi_control_BREADY,
	sum_12_s_axi_control_BVALID,
	sum_12_s_axi_control_BRESP,
	sum_13_m_axi_gmem_ARREADY,
	sum_13_m_axi_gmem_ARVALID,
	sum_13_m_axi_gmem_ARID,
	sum_13_m_axi_gmem_ARADDR,
	sum_13_m_axi_gmem_ARLEN,
	sum_13_m_axi_gmem_ARSIZE,
	sum_13_m_axi_gmem_ARBURST,
	sum_13_m_axi_gmem_ARLOCK,
	sum_13_m_axi_gmem_ARCACHE,
	sum_13_m_axi_gmem_ARPROT,
	sum_13_m_axi_gmem_ARQOS,
	sum_13_m_axi_gmem_ARREGION,
	sum_13_m_axi_gmem_ARUSER,
	sum_13_m_axi_gmem_RREADY,
	sum_13_m_axi_gmem_RVALID,
	sum_13_m_axi_gmem_RID,
	sum_13_m_axi_gmem_RDATA,
	sum_13_m_axi_gmem_RRESP,
	sum_13_m_axi_gmem_RLAST,
	sum_13_m_axi_gmem_RUSER,
	sum_13_m_axi_gmem_AWREADY,
	sum_13_m_axi_gmem_AWVALID,
	sum_13_m_axi_gmem_AWID,
	sum_13_m_axi_gmem_AWADDR,
	sum_13_m_axi_gmem_AWLEN,
	sum_13_m_axi_gmem_AWSIZE,
	sum_13_m_axi_gmem_AWBURST,
	sum_13_m_axi_gmem_AWLOCK,
	sum_13_m_axi_gmem_AWCACHE,
	sum_13_m_axi_gmem_AWPROT,
	sum_13_m_axi_gmem_AWQOS,
	sum_13_m_axi_gmem_AWREGION,
	sum_13_m_axi_gmem_AWUSER,
	sum_13_m_axi_gmem_WREADY,
	sum_13_m_axi_gmem_WVALID,
	sum_13_m_axi_gmem_WDATA,
	sum_13_m_axi_gmem_WSTRB,
	sum_13_m_axi_gmem_WLAST,
	sum_13_m_axi_gmem_WUSER,
	sum_13_m_axi_gmem_BREADY,
	sum_13_m_axi_gmem_BVALID,
	sum_13_m_axi_gmem_BID,
	sum_13_m_axi_gmem_BRESP,
	sum_13_m_axi_gmem_BUSER,
	sum_13_s_axi_control_ARREADY,
	sum_13_s_axi_control_ARVALID,
	sum_13_s_axi_control_ARADDR,
	sum_13_s_axi_control_RREADY,
	sum_13_s_axi_control_RVALID,
	sum_13_s_axi_control_RDATA,
	sum_13_s_axi_control_RRESP,
	sum_13_s_axi_control_AWREADY,
	sum_13_s_axi_control_AWVALID,
	sum_13_s_axi_control_AWADDR,
	sum_13_s_axi_control_WREADY,
	sum_13_s_axi_control_WVALID,
	sum_13_s_axi_control_WDATA,
	sum_13_s_axi_control_WSTRB,
	sum_13_s_axi_control_BREADY,
	sum_13_s_axi_control_BVALID,
	sum_13_s_axi_control_BRESP,
	sum_14_m_axi_gmem_ARREADY,
	sum_14_m_axi_gmem_ARVALID,
	sum_14_m_axi_gmem_ARID,
	sum_14_m_axi_gmem_ARADDR,
	sum_14_m_axi_gmem_ARLEN,
	sum_14_m_axi_gmem_ARSIZE,
	sum_14_m_axi_gmem_ARBURST,
	sum_14_m_axi_gmem_ARLOCK,
	sum_14_m_axi_gmem_ARCACHE,
	sum_14_m_axi_gmem_ARPROT,
	sum_14_m_axi_gmem_ARQOS,
	sum_14_m_axi_gmem_ARREGION,
	sum_14_m_axi_gmem_ARUSER,
	sum_14_m_axi_gmem_RREADY,
	sum_14_m_axi_gmem_RVALID,
	sum_14_m_axi_gmem_RID,
	sum_14_m_axi_gmem_RDATA,
	sum_14_m_axi_gmem_RRESP,
	sum_14_m_axi_gmem_RLAST,
	sum_14_m_axi_gmem_RUSER,
	sum_14_m_axi_gmem_AWREADY,
	sum_14_m_axi_gmem_AWVALID,
	sum_14_m_axi_gmem_AWID,
	sum_14_m_axi_gmem_AWADDR,
	sum_14_m_axi_gmem_AWLEN,
	sum_14_m_axi_gmem_AWSIZE,
	sum_14_m_axi_gmem_AWBURST,
	sum_14_m_axi_gmem_AWLOCK,
	sum_14_m_axi_gmem_AWCACHE,
	sum_14_m_axi_gmem_AWPROT,
	sum_14_m_axi_gmem_AWQOS,
	sum_14_m_axi_gmem_AWREGION,
	sum_14_m_axi_gmem_AWUSER,
	sum_14_m_axi_gmem_WREADY,
	sum_14_m_axi_gmem_WVALID,
	sum_14_m_axi_gmem_WDATA,
	sum_14_m_axi_gmem_WSTRB,
	sum_14_m_axi_gmem_WLAST,
	sum_14_m_axi_gmem_WUSER,
	sum_14_m_axi_gmem_BREADY,
	sum_14_m_axi_gmem_BVALID,
	sum_14_m_axi_gmem_BID,
	sum_14_m_axi_gmem_BRESP,
	sum_14_m_axi_gmem_BUSER,
	sum_14_s_axi_control_ARREADY,
	sum_14_s_axi_control_ARVALID,
	sum_14_s_axi_control_ARADDR,
	sum_14_s_axi_control_RREADY,
	sum_14_s_axi_control_RVALID,
	sum_14_s_axi_control_RDATA,
	sum_14_s_axi_control_RRESP,
	sum_14_s_axi_control_AWREADY,
	sum_14_s_axi_control_AWVALID,
	sum_14_s_axi_control_AWADDR,
	sum_14_s_axi_control_WREADY,
	sum_14_s_axi_control_WVALID,
	sum_14_s_axi_control_WDATA,
	sum_14_s_axi_control_WSTRB,
	sum_14_s_axi_control_BREADY,
	sum_14_s_axi_control_BVALID,
	sum_14_s_axi_control_BRESP,
	sum_15_m_axi_gmem_ARREADY,
	sum_15_m_axi_gmem_ARVALID,
	sum_15_m_axi_gmem_ARID,
	sum_15_m_axi_gmem_ARADDR,
	sum_15_m_axi_gmem_ARLEN,
	sum_15_m_axi_gmem_ARSIZE,
	sum_15_m_axi_gmem_ARBURST,
	sum_15_m_axi_gmem_ARLOCK,
	sum_15_m_axi_gmem_ARCACHE,
	sum_15_m_axi_gmem_ARPROT,
	sum_15_m_axi_gmem_ARQOS,
	sum_15_m_axi_gmem_ARREGION,
	sum_15_m_axi_gmem_ARUSER,
	sum_15_m_axi_gmem_RREADY,
	sum_15_m_axi_gmem_RVALID,
	sum_15_m_axi_gmem_RID,
	sum_15_m_axi_gmem_RDATA,
	sum_15_m_axi_gmem_RRESP,
	sum_15_m_axi_gmem_RLAST,
	sum_15_m_axi_gmem_RUSER,
	sum_15_m_axi_gmem_AWREADY,
	sum_15_m_axi_gmem_AWVALID,
	sum_15_m_axi_gmem_AWID,
	sum_15_m_axi_gmem_AWADDR,
	sum_15_m_axi_gmem_AWLEN,
	sum_15_m_axi_gmem_AWSIZE,
	sum_15_m_axi_gmem_AWBURST,
	sum_15_m_axi_gmem_AWLOCK,
	sum_15_m_axi_gmem_AWCACHE,
	sum_15_m_axi_gmem_AWPROT,
	sum_15_m_axi_gmem_AWQOS,
	sum_15_m_axi_gmem_AWREGION,
	sum_15_m_axi_gmem_AWUSER,
	sum_15_m_axi_gmem_WREADY,
	sum_15_m_axi_gmem_WVALID,
	sum_15_m_axi_gmem_WDATA,
	sum_15_m_axi_gmem_WSTRB,
	sum_15_m_axi_gmem_WLAST,
	sum_15_m_axi_gmem_WUSER,
	sum_15_m_axi_gmem_BREADY,
	sum_15_m_axi_gmem_BVALID,
	sum_15_m_axi_gmem_BID,
	sum_15_m_axi_gmem_BRESP,
	sum_15_m_axi_gmem_BUSER,
	sum_15_s_axi_control_ARREADY,
	sum_15_s_axi_control_ARVALID,
	sum_15_s_axi_control_ARADDR,
	sum_15_s_axi_control_RREADY,
	sum_15_s_axi_control_RVALID,
	sum_15_s_axi_control_RDATA,
	sum_15_s_axi_control_RRESP,
	sum_15_s_axi_control_AWREADY,
	sum_15_s_axi_control_AWVALID,
	sum_15_s_axi_control_AWADDR,
	sum_15_s_axi_control_WREADY,
	sum_15_s_axi_control_WVALID,
	sum_15_s_axi_control_WDATA,
	sum_15_s_axi_control_WSTRB,
	sum_15_s_axi_control_BREADY,
	sum_15_s_axi_control_BVALID,
	sum_15_s_axi_control_BRESP,
	sum_16_m_axi_gmem_ARREADY,
	sum_16_m_axi_gmem_ARVALID,
	sum_16_m_axi_gmem_ARID,
	sum_16_m_axi_gmem_ARADDR,
	sum_16_m_axi_gmem_ARLEN,
	sum_16_m_axi_gmem_ARSIZE,
	sum_16_m_axi_gmem_ARBURST,
	sum_16_m_axi_gmem_ARLOCK,
	sum_16_m_axi_gmem_ARCACHE,
	sum_16_m_axi_gmem_ARPROT,
	sum_16_m_axi_gmem_ARQOS,
	sum_16_m_axi_gmem_ARREGION,
	sum_16_m_axi_gmem_ARUSER,
	sum_16_m_axi_gmem_RREADY,
	sum_16_m_axi_gmem_RVALID,
	sum_16_m_axi_gmem_RID,
	sum_16_m_axi_gmem_RDATA,
	sum_16_m_axi_gmem_RRESP,
	sum_16_m_axi_gmem_RLAST,
	sum_16_m_axi_gmem_RUSER,
	sum_16_m_axi_gmem_AWREADY,
	sum_16_m_axi_gmem_AWVALID,
	sum_16_m_axi_gmem_AWID,
	sum_16_m_axi_gmem_AWADDR,
	sum_16_m_axi_gmem_AWLEN,
	sum_16_m_axi_gmem_AWSIZE,
	sum_16_m_axi_gmem_AWBURST,
	sum_16_m_axi_gmem_AWLOCK,
	sum_16_m_axi_gmem_AWCACHE,
	sum_16_m_axi_gmem_AWPROT,
	sum_16_m_axi_gmem_AWQOS,
	sum_16_m_axi_gmem_AWREGION,
	sum_16_m_axi_gmem_AWUSER,
	sum_16_m_axi_gmem_WREADY,
	sum_16_m_axi_gmem_WVALID,
	sum_16_m_axi_gmem_WDATA,
	sum_16_m_axi_gmem_WSTRB,
	sum_16_m_axi_gmem_WLAST,
	sum_16_m_axi_gmem_WUSER,
	sum_16_m_axi_gmem_BREADY,
	sum_16_m_axi_gmem_BVALID,
	sum_16_m_axi_gmem_BID,
	sum_16_m_axi_gmem_BRESP,
	sum_16_m_axi_gmem_BUSER,
	sum_16_s_axi_control_ARREADY,
	sum_16_s_axi_control_ARVALID,
	sum_16_s_axi_control_ARADDR,
	sum_16_s_axi_control_RREADY,
	sum_16_s_axi_control_RVALID,
	sum_16_s_axi_control_RDATA,
	sum_16_s_axi_control_RRESP,
	sum_16_s_axi_control_AWREADY,
	sum_16_s_axi_control_AWVALID,
	sum_16_s_axi_control_AWADDR,
	sum_16_s_axi_control_WREADY,
	sum_16_s_axi_control_WVALID,
	sum_16_s_axi_control_WDATA,
	sum_16_s_axi_control_WSTRB,
	sum_16_s_axi_control_BREADY,
	sum_16_s_axi_control_BVALID,
	sum_16_s_axi_control_BRESP,
	sum_17_m_axi_gmem_ARREADY,
	sum_17_m_axi_gmem_ARVALID,
	sum_17_m_axi_gmem_ARID,
	sum_17_m_axi_gmem_ARADDR,
	sum_17_m_axi_gmem_ARLEN,
	sum_17_m_axi_gmem_ARSIZE,
	sum_17_m_axi_gmem_ARBURST,
	sum_17_m_axi_gmem_ARLOCK,
	sum_17_m_axi_gmem_ARCACHE,
	sum_17_m_axi_gmem_ARPROT,
	sum_17_m_axi_gmem_ARQOS,
	sum_17_m_axi_gmem_ARREGION,
	sum_17_m_axi_gmem_ARUSER,
	sum_17_m_axi_gmem_RREADY,
	sum_17_m_axi_gmem_RVALID,
	sum_17_m_axi_gmem_RID,
	sum_17_m_axi_gmem_RDATA,
	sum_17_m_axi_gmem_RRESP,
	sum_17_m_axi_gmem_RLAST,
	sum_17_m_axi_gmem_RUSER,
	sum_17_m_axi_gmem_AWREADY,
	sum_17_m_axi_gmem_AWVALID,
	sum_17_m_axi_gmem_AWID,
	sum_17_m_axi_gmem_AWADDR,
	sum_17_m_axi_gmem_AWLEN,
	sum_17_m_axi_gmem_AWSIZE,
	sum_17_m_axi_gmem_AWBURST,
	sum_17_m_axi_gmem_AWLOCK,
	sum_17_m_axi_gmem_AWCACHE,
	sum_17_m_axi_gmem_AWPROT,
	sum_17_m_axi_gmem_AWQOS,
	sum_17_m_axi_gmem_AWREGION,
	sum_17_m_axi_gmem_AWUSER,
	sum_17_m_axi_gmem_WREADY,
	sum_17_m_axi_gmem_WVALID,
	sum_17_m_axi_gmem_WDATA,
	sum_17_m_axi_gmem_WSTRB,
	sum_17_m_axi_gmem_WLAST,
	sum_17_m_axi_gmem_WUSER,
	sum_17_m_axi_gmem_BREADY,
	sum_17_m_axi_gmem_BVALID,
	sum_17_m_axi_gmem_BID,
	sum_17_m_axi_gmem_BRESP,
	sum_17_m_axi_gmem_BUSER,
	sum_17_s_axi_control_ARREADY,
	sum_17_s_axi_control_ARVALID,
	sum_17_s_axi_control_ARADDR,
	sum_17_s_axi_control_RREADY,
	sum_17_s_axi_control_RVALID,
	sum_17_s_axi_control_RDATA,
	sum_17_s_axi_control_RRESP,
	sum_17_s_axi_control_AWREADY,
	sum_17_s_axi_control_AWVALID,
	sum_17_s_axi_control_AWADDR,
	sum_17_s_axi_control_WREADY,
	sum_17_s_axi_control_WVALID,
	sum_17_s_axi_control_WDATA,
	sum_17_s_axi_control_WSTRB,
	sum_17_s_axi_control_BREADY,
	sum_17_s_axi_control_BVALID,
	sum_17_s_axi_control_BRESP,
	sum_18_m_axi_gmem_ARREADY,
	sum_18_m_axi_gmem_ARVALID,
	sum_18_m_axi_gmem_ARID,
	sum_18_m_axi_gmem_ARADDR,
	sum_18_m_axi_gmem_ARLEN,
	sum_18_m_axi_gmem_ARSIZE,
	sum_18_m_axi_gmem_ARBURST,
	sum_18_m_axi_gmem_ARLOCK,
	sum_18_m_axi_gmem_ARCACHE,
	sum_18_m_axi_gmem_ARPROT,
	sum_18_m_axi_gmem_ARQOS,
	sum_18_m_axi_gmem_ARREGION,
	sum_18_m_axi_gmem_ARUSER,
	sum_18_m_axi_gmem_RREADY,
	sum_18_m_axi_gmem_RVALID,
	sum_18_m_axi_gmem_RID,
	sum_18_m_axi_gmem_RDATA,
	sum_18_m_axi_gmem_RRESP,
	sum_18_m_axi_gmem_RLAST,
	sum_18_m_axi_gmem_RUSER,
	sum_18_m_axi_gmem_AWREADY,
	sum_18_m_axi_gmem_AWVALID,
	sum_18_m_axi_gmem_AWID,
	sum_18_m_axi_gmem_AWADDR,
	sum_18_m_axi_gmem_AWLEN,
	sum_18_m_axi_gmem_AWSIZE,
	sum_18_m_axi_gmem_AWBURST,
	sum_18_m_axi_gmem_AWLOCK,
	sum_18_m_axi_gmem_AWCACHE,
	sum_18_m_axi_gmem_AWPROT,
	sum_18_m_axi_gmem_AWQOS,
	sum_18_m_axi_gmem_AWREGION,
	sum_18_m_axi_gmem_AWUSER,
	sum_18_m_axi_gmem_WREADY,
	sum_18_m_axi_gmem_WVALID,
	sum_18_m_axi_gmem_WDATA,
	sum_18_m_axi_gmem_WSTRB,
	sum_18_m_axi_gmem_WLAST,
	sum_18_m_axi_gmem_WUSER,
	sum_18_m_axi_gmem_BREADY,
	sum_18_m_axi_gmem_BVALID,
	sum_18_m_axi_gmem_BID,
	sum_18_m_axi_gmem_BRESP,
	sum_18_m_axi_gmem_BUSER,
	sum_18_s_axi_control_ARREADY,
	sum_18_s_axi_control_ARVALID,
	sum_18_s_axi_control_ARADDR,
	sum_18_s_axi_control_RREADY,
	sum_18_s_axi_control_RVALID,
	sum_18_s_axi_control_RDATA,
	sum_18_s_axi_control_RRESP,
	sum_18_s_axi_control_AWREADY,
	sum_18_s_axi_control_AWVALID,
	sum_18_s_axi_control_AWADDR,
	sum_18_s_axi_control_WREADY,
	sum_18_s_axi_control_WVALID,
	sum_18_s_axi_control_WDATA,
	sum_18_s_axi_control_WSTRB,
	sum_18_s_axi_control_BREADY,
	sum_18_s_axi_control_BVALID,
	sum_18_s_axi_control_BRESP,
	sum_19_m_axi_gmem_ARREADY,
	sum_19_m_axi_gmem_ARVALID,
	sum_19_m_axi_gmem_ARID,
	sum_19_m_axi_gmem_ARADDR,
	sum_19_m_axi_gmem_ARLEN,
	sum_19_m_axi_gmem_ARSIZE,
	sum_19_m_axi_gmem_ARBURST,
	sum_19_m_axi_gmem_ARLOCK,
	sum_19_m_axi_gmem_ARCACHE,
	sum_19_m_axi_gmem_ARPROT,
	sum_19_m_axi_gmem_ARQOS,
	sum_19_m_axi_gmem_ARREGION,
	sum_19_m_axi_gmem_ARUSER,
	sum_19_m_axi_gmem_RREADY,
	sum_19_m_axi_gmem_RVALID,
	sum_19_m_axi_gmem_RID,
	sum_19_m_axi_gmem_RDATA,
	sum_19_m_axi_gmem_RRESP,
	sum_19_m_axi_gmem_RLAST,
	sum_19_m_axi_gmem_RUSER,
	sum_19_m_axi_gmem_AWREADY,
	sum_19_m_axi_gmem_AWVALID,
	sum_19_m_axi_gmem_AWID,
	sum_19_m_axi_gmem_AWADDR,
	sum_19_m_axi_gmem_AWLEN,
	sum_19_m_axi_gmem_AWSIZE,
	sum_19_m_axi_gmem_AWBURST,
	sum_19_m_axi_gmem_AWLOCK,
	sum_19_m_axi_gmem_AWCACHE,
	sum_19_m_axi_gmem_AWPROT,
	sum_19_m_axi_gmem_AWQOS,
	sum_19_m_axi_gmem_AWREGION,
	sum_19_m_axi_gmem_AWUSER,
	sum_19_m_axi_gmem_WREADY,
	sum_19_m_axi_gmem_WVALID,
	sum_19_m_axi_gmem_WDATA,
	sum_19_m_axi_gmem_WSTRB,
	sum_19_m_axi_gmem_WLAST,
	sum_19_m_axi_gmem_WUSER,
	sum_19_m_axi_gmem_BREADY,
	sum_19_m_axi_gmem_BVALID,
	sum_19_m_axi_gmem_BID,
	sum_19_m_axi_gmem_BRESP,
	sum_19_m_axi_gmem_BUSER,
	sum_19_s_axi_control_ARREADY,
	sum_19_s_axi_control_ARVALID,
	sum_19_s_axi_control_ARADDR,
	sum_19_s_axi_control_RREADY,
	sum_19_s_axi_control_RVALID,
	sum_19_s_axi_control_RDATA,
	sum_19_s_axi_control_RRESP,
	sum_19_s_axi_control_AWREADY,
	sum_19_s_axi_control_AWVALID,
	sum_19_s_axi_control_AWADDR,
	sum_19_s_axi_control_WREADY,
	sum_19_s_axi_control_WVALID,
	sum_19_s_axi_control_WDATA,
	sum_19_s_axi_control_WSTRB,
	sum_19_s_axi_control_BREADY,
	sum_19_s_axi_control_BVALID,
	sum_19_s_axi_control_BRESP,
	sum_20_m_axi_gmem_ARREADY,
	sum_20_m_axi_gmem_ARVALID,
	sum_20_m_axi_gmem_ARID,
	sum_20_m_axi_gmem_ARADDR,
	sum_20_m_axi_gmem_ARLEN,
	sum_20_m_axi_gmem_ARSIZE,
	sum_20_m_axi_gmem_ARBURST,
	sum_20_m_axi_gmem_ARLOCK,
	sum_20_m_axi_gmem_ARCACHE,
	sum_20_m_axi_gmem_ARPROT,
	sum_20_m_axi_gmem_ARQOS,
	sum_20_m_axi_gmem_ARREGION,
	sum_20_m_axi_gmem_ARUSER,
	sum_20_m_axi_gmem_RREADY,
	sum_20_m_axi_gmem_RVALID,
	sum_20_m_axi_gmem_RID,
	sum_20_m_axi_gmem_RDATA,
	sum_20_m_axi_gmem_RRESP,
	sum_20_m_axi_gmem_RLAST,
	sum_20_m_axi_gmem_RUSER,
	sum_20_m_axi_gmem_AWREADY,
	sum_20_m_axi_gmem_AWVALID,
	sum_20_m_axi_gmem_AWID,
	sum_20_m_axi_gmem_AWADDR,
	sum_20_m_axi_gmem_AWLEN,
	sum_20_m_axi_gmem_AWSIZE,
	sum_20_m_axi_gmem_AWBURST,
	sum_20_m_axi_gmem_AWLOCK,
	sum_20_m_axi_gmem_AWCACHE,
	sum_20_m_axi_gmem_AWPROT,
	sum_20_m_axi_gmem_AWQOS,
	sum_20_m_axi_gmem_AWREGION,
	sum_20_m_axi_gmem_AWUSER,
	sum_20_m_axi_gmem_WREADY,
	sum_20_m_axi_gmem_WVALID,
	sum_20_m_axi_gmem_WDATA,
	sum_20_m_axi_gmem_WSTRB,
	sum_20_m_axi_gmem_WLAST,
	sum_20_m_axi_gmem_WUSER,
	sum_20_m_axi_gmem_BREADY,
	sum_20_m_axi_gmem_BVALID,
	sum_20_m_axi_gmem_BID,
	sum_20_m_axi_gmem_BRESP,
	sum_20_m_axi_gmem_BUSER,
	sum_20_s_axi_control_ARREADY,
	sum_20_s_axi_control_ARVALID,
	sum_20_s_axi_control_ARADDR,
	sum_20_s_axi_control_RREADY,
	sum_20_s_axi_control_RVALID,
	sum_20_s_axi_control_RDATA,
	sum_20_s_axi_control_RRESP,
	sum_20_s_axi_control_AWREADY,
	sum_20_s_axi_control_AWVALID,
	sum_20_s_axi_control_AWADDR,
	sum_20_s_axi_control_WREADY,
	sum_20_s_axi_control_WVALID,
	sum_20_s_axi_control_WDATA,
	sum_20_s_axi_control_WSTRB,
	sum_20_s_axi_control_BREADY,
	sum_20_s_axi_control_BVALID,
	sum_20_s_axi_control_BRESP,
	sum_21_m_axi_gmem_ARREADY,
	sum_21_m_axi_gmem_ARVALID,
	sum_21_m_axi_gmem_ARID,
	sum_21_m_axi_gmem_ARADDR,
	sum_21_m_axi_gmem_ARLEN,
	sum_21_m_axi_gmem_ARSIZE,
	sum_21_m_axi_gmem_ARBURST,
	sum_21_m_axi_gmem_ARLOCK,
	sum_21_m_axi_gmem_ARCACHE,
	sum_21_m_axi_gmem_ARPROT,
	sum_21_m_axi_gmem_ARQOS,
	sum_21_m_axi_gmem_ARREGION,
	sum_21_m_axi_gmem_ARUSER,
	sum_21_m_axi_gmem_RREADY,
	sum_21_m_axi_gmem_RVALID,
	sum_21_m_axi_gmem_RID,
	sum_21_m_axi_gmem_RDATA,
	sum_21_m_axi_gmem_RRESP,
	sum_21_m_axi_gmem_RLAST,
	sum_21_m_axi_gmem_RUSER,
	sum_21_m_axi_gmem_AWREADY,
	sum_21_m_axi_gmem_AWVALID,
	sum_21_m_axi_gmem_AWID,
	sum_21_m_axi_gmem_AWADDR,
	sum_21_m_axi_gmem_AWLEN,
	sum_21_m_axi_gmem_AWSIZE,
	sum_21_m_axi_gmem_AWBURST,
	sum_21_m_axi_gmem_AWLOCK,
	sum_21_m_axi_gmem_AWCACHE,
	sum_21_m_axi_gmem_AWPROT,
	sum_21_m_axi_gmem_AWQOS,
	sum_21_m_axi_gmem_AWREGION,
	sum_21_m_axi_gmem_AWUSER,
	sum_21_m_axi_gmem_WREADY,
	sum_21_m_axi_gmem_WVALID,
	sum_21_m_axi_gmem_WDATA,
	sum_21_m_axi_gmem_WSTRB,
	sum_21_m_axi_gmem_WLAST,
	sum_21_m_axi_gmem_WUSER,
	sum_21_m_axi_gmem_BREADY,
	sum_21_m_axi_gmem_BVALID,
	sum_21_m_axi_gmem_BID,
	sum_21_m_axi_gmem_BRESP,
	sum_21_m_axi_gmem_BUSER,
	sum_21_s_axi_control_ARREADY,
	sum_21_s_axi_control_ARVALID,
	sum_21_s_axi_control_ARADDR,
	sum_21_s_axi_control_RREADY,
	sum_21_s_axi_control_RVALID,
	sum_21_s_axi_control_RDATA,
	sum_21_s_axi_control_RRESP,
	sum_21_s_axi_control_AWREADY,
	sum_21_s_axi_control_AWVALID,
	sum_21_s_axi_control_AWADDR,
	sum_21_s_axi_control_WREADY,
	sum_21_s_axi_control_WVALID,
	sum_21_s_axi_control_WDATA,
	sum_21_s_axi_control_WSTRB,
	sum_21_s_axi_control_BREADY,
	sum_21_s_axi_control_BVALID,
	sum_21_s_axi_control_BRESP,
	sum_22_m_axi_gmem_ARREADY,
	sum_22_m_axi_gmem_ARVALID,
	sum_22_m_axi_gmem_ARID,
	sum_22_m_axi_gmem_ARADDR,
	sum_22_m_axi_gmem_ARLEN,
	sum_22_m_axi_gmem_ARSIZE,
	sum_22_m_axi_gmem_ARBURST,
	sum_22_m_axi_gmem_ARLOCK,
	sum_22_m_axi_gmem_ARCACHE,
	sum_22_m_axi_gmem_ARPROT,
	sum_22_m_axi_gmem_ARQOS,
	sum_22_m_axi_gmem_ARREGION,
	sum_22_m_axi_gmem_ARUSER,
	sum_22_m_axi_gmem_RREADY,
	sum_22_m_axi_gmem_RVALID,
	sum_22_m_axi_gmem_RID,
	sum_22_m_axi_gmem_RDATA,
	sum_22_m_axi_gmem_RRESP,
	sum_22_m_axi_gmem_RLAST,
	sum_22_m_axi_gmem_RUSER,
	sum_22_m_axi_gmem_AWREADY,
	sum_22_m_axi_gmem_AWVALID,
	sum_22_m_axi_gmem_AWID,
	sum_22_m_axi_gmem_AWADDR,
	sum_22_m_axi_gmem_AWLEN,
	sum_22_m_axi_gmem_AWSIZE,
	sum_22_m_axi_gmem_AWBURST,
	sum_22_m_axi_gmem_AWLOCK,
	sum_22_m_axi_gmem_AWCACHE,
	sum_22_m_axi_gmem_AWPROT,
	sum_22_m_axi_gmem_AWQOS,
	sum_22_m_axi_gmem_AWREGION,
	sum_22_m_axi_gmem_AWUSER,
	sum_22_m_axi_gmem_WREADY,
	sum_22_m_axi_gmem_WVALID,
	sum_22_m_axi_gmem_WDATA,
	sum_22_m_axi_gmem_WSTRB,
	sum_22_m_axi_gmem_WLAST,
	sum_22_m_axi_gmem_WUSER,
	sum_22_m_axi_gmem_BREADY,
	sum_22_m_axi_gmem_BVALID,
	sum_22_m_axi_gmem_BID,
	sum_22_m_axi_gmem_BRESP,
	sum_22_m_axi_gmem_BUSER,
	sum_22_s_axi_control_ARREADY,
	sum_22_s_axi_control_ARVALID,
	sum_22_s_axi_control_ARADDR,
	sum_22_s_axi_control_RREADY,
	sum_22_s_axi_control_RVALID,
	sum_22_s_axi_control_RDATA,
	sum_22_s_axi_control_RRESP,
	sum_22_s_axi_control_AWREADY,
	sum_22_s_axi_control_AWVALID,
	sum_22_s_axi_control_AWADDR,
	sum_22_s_axi_control_WREADY,
	sum_22_s_axi_control_WVALID,
	sum_22_s_axi_control_WDATA,
	sum_22_s_axi_control_WSTRB,
	sum_22_s_axi_control_BREADY,
	sum_22_s_axi_control_BVALID,
	sum_22_s_axi_control_BRESP,
	sum_23_m_axi_gmem_ARREADY,
	sum_23_m_axi_gmem_ARVALID,
	sum_23_m_axi_gmem_ARID,
	sum_23_m_axi_gmem_ARADDR,
	sum_23_m_axi_gmem_ARLEN,
	sum_23_m_axi_gmem_ARSIZE,
	sum_23_m_axi_gmem_ARBURST,
	sum_23_m_axi_gmem_ARLOCK,
	sum_23_m_axi_gmem_ARCACHE,
	sum_23_m_axi_gmem_ARPROT,
	sum_23_m_axi_gmem_ARQOS,
	sum_23_m_axi_gmem_ARREGION,
	sum_23_m_axi_gmem_ARUSER,
	sum_23_m_axi_gmem_RREADY,
	sum_23_m_axi_gmem_RVALID,
	sum_23_m_axi_gmem_RID,
	sum_23_m_axi_gmem_RDATA,
	sum_23_m_axi_gmem_RRESP,
	sum_23_m_axi_gmem_RLAST,
	sum_23_m_axi_gmem_RUSER,
	sum_23_m_axi_gmem_AWREADY,
	sum_23_m_axi_gmem_AWVALID,
	sum_23_m_axi_gmem_AWID,
	sum_23_m_axi_gmem_AWADDR,
	sum_23_m_axi_gmem_AWLEN,
	sum_23_m_axi_gmem_AWSIZE,
	sum_23_m_axi_gmem_AWBURST,
	sum_23_m_axi_gmem_AWLOCK,
	sum_23_m_axi_gmem_AWCACHE,
	sum_23_m_axi_gmem_AWPROT,
	sum_23_m_axi_gmem_AWQOS,
	sum_23_m_axi_gmem_AWREGION,
	sum_23_m_axi_gmem_AWUSER,
	sum_23_m_axi_gmem_WREADY,
	sum_23_m_axi_gmem_WVALID,
	sum_23_m_axi_gmem_WDATA,
	sum_23_m_axi_gmem_WSTRB,
	sum_23_m_axi_gmem_WLAST,
	sum_23_m_axi_gmem_WUSER,
	sum_23_m_axi_gmem_BREADY,
	sum_23_m_axi_gmem_BVALID,
	sum_23_m_axi_gmem_BID,
	sum_23_m_axi_gmem_BRESP,
	sum_23_m_axi_gmem_BUSER,
	sum_23_s_axi_control_ARREADY,
	sum_23_s_axi_control_ARVALID,
	sum_23_s_axi_control_ARADDR,
	sum_23_s_axi_control_RREADY,
	sum_23_s_axi_control_RVALID,
	sum_23_s_axi_control_RDATA,
	sum_23_s_axi_control_RRESP,
	sum_23_s_axi_control_AWREADY,
	sum_23_s_axi_control_AWVALID,
	sum_23_s_axi_control_AWADDR,
	sum_23_s_axi_control_WREADY,
	sum_23_s_axi_control_WVALID,
	sum_23_s_axi_control_WDATA,
	sum_23_s_axi_control_WSTRB,
	sum_23_s_axi_control_BREADY,
	sum_23_s_axi_control_BVALID,
	sum_23_s_axi_control_BRESP,
	sum_24_m_axi_gmem_ARREADY,
	sum_24_m_axi_gmem_ARVALID,
	sum_24_m_axi_gmem_ARID,
	sum_24_m_axi_gmem_ARADDR,
	sum_24_m_axi_gmem_ARLEN,
	sum_24_m_axi_gmem_ARSIZE,
	sum_24_m_axi_gmem_ARBURST,
	sum_24_m_axi_gmem_ARLOCK,
	sum_24_m_axi_gmem_ARCACHE,
	sum_24_m_axi_gmem_ARPROT,
	sum_24_m_axi_gmem_ARQOS,
	sum_24_m_axi_gmem_ARREGION,
	sum_24_m_axi_gmem_ARUSER,
	sum_24_m_axi_gmem_RREADY,
	sum_24_m_axi_gmem_RVALID,
	sum_24_m_axi_gmem_RID,
	sum_24_m_axi_gmem_RDATA,
	sum_24_m_axi_gmem_RRESP,
	sum_24_m_axi_gmem_RLAST,
	sum_24_m_axi_gmem_RUSER,
	sum_24_m_axi_gmem_AWREADY,
	sum_24_m_axi_gmem_AWVALID,
	sum_24_m_axi_gmem_AWID,
	sum_24_m_axi_gmem_AWADDR,
	sum_24_m_axi_gmem_AWLEN,
	sum_24_m_axi_gmem_AWSIZE,
	sum_24_m_axi_gmem_AWBURST,
	sum_24_m_axi_gmem_AWLOCK,
	sum_24_m_axi_gmem_AWCACHE,
	sum_24_m_axi_gmem_AWPROT,
	sum_24_m_axi_gmem_AWQOS,
	sum_24_m_axi_gmem_AWREGION,
	sum_24_m_axi_gmem_AWUSER,
	sum_24_m_axi_gmem_WREADY,
	sum_24_m_axi_gmem_WVALID,
	sum_24_m_axi_gmem_WDATA,
	sum_24_m_axi_gmem_WSTRB,
	sum_24_m_axi_gmem_WLAST,
	sum_24_m_axi_gmem_WUSER,
	sum_24_m_axi_gmem_BREADY,
	sum_24_m_axi_gmem_BVALID,
	sum_24_m_axi_gmem_BID,
	sum_24_m_axi_gmem_BRESP,
	sum_24_m_axi_gmem_BUSER,
	sum_24_s_axi_control_ARREADY,
	sum_24_s_axi_control_ARVALID,
	sum_24_s_axi_control_ARADDR,
	sum_24_s_axi_control_RREADY,
	sum_24_s_axi_control_RVALID,
	sum_24_s_axi_control_RDATA,
	sum_24_s_axi_control_RRESP,
	sum_24_s_axi_control_AWREADY,
	sum_24_s_axi_control_AWVALID,
	sum_24_s_axi_control_AWADDR,
	sum_24_s_axi_control_WREADY,
	sum_24_s_axi_control_WVALID,
	sum_24_s_axi_control_WDATA,
	sum_24_s_axi_control_WSTRB,
	sum_24_s_axi_control_BREADY,
	sum_24_s_axi_control_BVALID,
	sum_24_s_axi_control_BRESP,
	sum_25_m_axi_gmem_ARREADY,
	sum_25_m_axi_gmem_ARVALID,
	sum_25_m_axi_gmem_ARID,
	sum_25_m_axi_gmem_ARADDR,
	sum_25_m_axi_gmem_ARLEN,
	sum_25_m_axi_gmem_ARSIZE,
	sum_25_m_axi_gmem_ARBURST,
	sum_25_m_axi_gmem_ARLOCK,
	sum_25_m_axi_gmem_ARCACHE,
	sum_25_m_axi_gmem_ARPROT,
	sum_25_m_axi_gmem_ARQOS,
	sum_25_m_axi_gmem_ARREGION,
	sum_25_m_axi_gmem_ARUSER,
	sum_25_m_axi_gmem_RREADY,
	sum_25_m_axi_gmem_RVALID,
	sum_25_m_axi_gmem_RID,
	sum_25_m_axi_gmem_RDATA,
	sum_25_m_axi_gmem_RRESP,
	sum_25_m_axi_gmem_RLAST,
	sum_25_m_axi_gmem_RUSER,
	sum_25_m_axi_gmem_AWREADY,
	sum_25_m_axi_gmem_AWVALID,
	sum_25_m_axi_gmem_AWID,
	sum_25_m_axi_gmem_AWADDR,
	sum_25_m_axi_gmem_AWLEN,
	sum_25_m_axi_gmem_AWSIZE,
	sum_25_m_axi_gmem_AWBURST,
	sum_25_m_axi_gmem_AWLOCK,
	sum_25_m_axi_gmem_AWCACHE,
	sum_25_m_axi_gmem_AWPROT,
	sum_25_m_axi_gmem_AWQOS,
	sum_25_m_axi_gmem_AWREGION,
	sum_25_m_axi_gmem_AWUSER,
	sum_25_m_axi_gmem_WREADY,
	sum_25_m_axi_gmem_WVALID,
	sum_25_m_axi_gmem_WDATA,
	sum_25_m_axi_gmem_WSTRB,
	sum_25_m_axi_gmem_WLAST,
	sum_25_m_axi_gmem_WUSER,
	sum_25_m_axi_gmem_BREADY,
	sum_25_m_axi_gmem_BVALID,
	sum_25_m_axi_gmem_BID,
	sum_25_m_axi_gmem_BRESP,
	sum_25_m_axi_gmem_BUSER,
	sum_25_s_axi_control_ARREADY,
	sum_25_s_axi_control_ARVALID,
	sum_25_s_axi_control_ARADDR,
	sum_25_s_axi_control_RREADY,
	sum_25_s_axi_control_RVALID,
	sum_25_s_axi_control_RDATA,
	sum_25_s_axi_control_RRESP,
	sum_25_s_axi_control_AWREADY,
	sum_25_s_axi_control_AWVALID,
	sum_25_s_axi_control_AWADDR,
	sum_25_s_axi_control_WREADY,
	sum_25_s_axi_control_WVALID,
	sum_25_s_axi_control_WDATA,
	sum_25_s_axi_control_WSTRB,
	sum_25_s_axi_control_BREADY,
	sum_25_s_axi_control_BVALID,
	sum_25_s_axi_control_BRESP,
	sum_26_m_axi_gmem_ARREADY,
	sum_26_m_axi_gmem_ARVALID,
	sum_26_m_axi_gmem_ARID,
	sum_26_m_axi_gmem_ARADDR,
	sum_26_m_axi_gmem_ARLEN,
	sum_26_m_axi_gmem_ARSIZE,
	sum_26_m_axi_gmem_ARBURST,
	sum_26_m_axi_gmem_ARLOCK,
	sum_26_m_axi_gmem_ARCACHE,
	sum_26_m_axi_gmem_ARPROT,
	sum_26_m_axi_gmem_ARQOS,
	sum_26_m_axi_gmem_ARREGION,
	sum_26_m_axi_gmem_ARUSER,
	sum_26_m_axi_gmem_RREADY,
	sum_26_m_axi_gmem_RVALID,
	sum_26_m_axi_gmem_RID,
	sum_26_m_axi_gmem_RDATA,
	sum_26_m_axi_gmem_RRESP,
	sum_26_m_axi_gmem_RLAST,
	sum_26_m_axi_gmem_RUSER,
	sum_26_m_axi_gmem_AWREADY,
	sum_26_m_axi_gmem_AWVALID,
	sum_26_m_axi_gmem_AWID,
	sum_26_m_axi_gmem_AWADDR,
	sum_26_m_axi_gmem_AWLEN,
	sum_26_m_axi_gmem_AWSIZE,
	sum_26_m_axi_gmem_AWBURST,
	sum_26_m_axi_gmem_AWLOCK,
	sum_26_m_axi_gmem_AWCACHE,
	sum_26_m_axi_gmem_AWPROT,
	sum_26_m_axi_gmem_AWQOS,
	sum_26_m_axi_gmem_AWREGION,
	sum_26_m_axi_gmem_AWUSER,
	sum_26_m_axi_gmem_WREADY,
	sum_26_m_axi_gmem_WVALID,
	sum_26_m_axi_gmem_WDATA,
	sum_26_m_axi_gmem_WSTRB,
	sum_26_m_axi_gmem_WLAST,
	sum_26_m_axi_gmem_WUSER,
	sum_26_m_axi_gmem_BREADY,
	sum_26_m_axi_gmem_BVALID,
	sum_26_m_axi_gmem_BID,
	sum_26_m_axi_gmem_BRESP,
	sum_26_m_axi_gmem_BUSER,
	sum_26_s_axi_control_ARREADY,
	sum_26_s_axi_control_ARVALID,
	sum_26_s_axi_control_ARADDR,
	sum_26_s_axi_control_RREADY,
	sum_26_s_axi_control_RVALID,
	sum_26_s_axi_control_RDATA,
	sum_26_s_axi_control_RRESP,
	sum_26_s_axi_control_AWREADY,
	sum_26_s_axi_control_AWVALID,
	sum_26_s_axi_control_AWADDR,
	sum_26_s_axi_control_WREADY,
	sum_26_s_axi_control_WVALID,
	sum_26_s_axi_control_WDATA,
	sum_26_s_axi_control_WSTRB,
	sum_26_s_axi_control_BREADY,
	sum_26_s_axi_control_BVALID,
	sum_26_s_axi_control_BRESP,
	sum_27_m_axi_gmem_ARREADY,
	sum_27_m_axi_gmem_ARVALID,
	sum_27_m_axi_gmem_ARID,
	sum_27_m_axi_gmem_ARADDR,
	sum_27_m_axi_gmem_ARLEN,
	sum_27_m_axi_gmem_ARSIZE,
	sum_27_m_axi_gmem_ARBURST,
	sum_27_m_axi_gmem_ARLOCK,
	sum_27_m_axi_gmem_ARCACHE,
	sum_27_m_axi_gmem_ARPROT,
	sum_27_m_axi_gmem_ARQOS,
	sum_27_m_axi_gmem_ARREGION,
	sum_27_m_axi_gmem_ARUSER,
	sum_27_m_axi_gmem_RREADY,
	sum_27_m_axi_gmem_RVALID,
	sum_27_m_axi_gmem_RID,
	sum_27_m_axi_gmem_RDATA,
	sum_27_m_axi_gmem_RRESP,
	sum_27_m_axi_gmem_RLAST,
	sum_27_m_axi_gmem_RUSER,
	sum_27_m_axi_gmem_AWREADY,
	sum_27_m_axi_gmem_AWVALID,
	sum_27_m_axi_gmem_AWID,
	sum_27_m_axi_gmem_AWADDR,
	sum_27_m_axi_gmem_AWLEN,
	sum_27_m_axi_gmem_AWSIZE,
	sum_27_m_axi_gmem_AWBURST,
	sum_27_m_axi_gmem_AWLOCK,
	sum_27_m_axi_gmem_AWCACHE,
	sum_27_m_axi_gmem_AWPROT,
	sum_27_m_axi_gmem_AWQOS,
	sum_27_m_axi_gmem_AWREGION,
	sum_27_m_axi_gmem_AWUSER,
	sum_27_m_axi_gmem_WREADY,
	sum_27_m_axi_gmem_WVALID,
	sum_27_m_axi_gmem_WDATA,
	sum_27_m_axi_gmem_WSTRB,
	sum_27_m_axi_gmem_WLAST,
	sum_27_m_axi_gmem_WUSER,
	sum_27_m_axi_gmem_BREADY,
	sum_27_m_axi_gmem_BVALID,
	sum_27_m_axi_gmem_BID,
	sum_27_m_axi_gmem_BRESP,
	sum_27_m_axi_gmem_BUSER,
	sum_27_s_axi_control_ARREADY,
	sum_27_s_axi_control_ARVALID,
	sum_27_s_axi_control_ARADDR,
	sum_27_s_axi_control_RREADY,
	sum_27_s_axi_control_RVALID,
	sum_27_s_axi_control_RDATA,
	sum_27_s_axi_control_RRESP,
	sum_27_s_axi_control_AWREADY,
	sum_27_s_axi_control_AWVALID,
	sum_27_s_axi_control_AWADDR,
	sum_27_s_axi_control_WREADY,
	sum_27_s_axi_control_WVALID,
	sum_27_s_axi_control_WDATA,
	sum_27_s_axi_control_WSTRB,
	sum_27_s_axi_control_BREADY,
	sum_27_s_axi_control_BVALID,
	sum_27_s_axi_control_BRESP,
	sum_28_m_axi_gmem_ARREADY,
	sum_28_m_axi_gmem_ARVALID,
	sum_28_m_axi_gmem_ARID,
	sum_28_m_axi_gmem_ARADDR,
	sum_28_m_axi_gmem_ARLEN,
	sum_28_m_axi_gmem_ARSIZE,
	sum_28_m_axi_gmem_ARBURST,
	sum_28_m_axi_gmem_ARLOCK,
	sum_28_m_axi_gmem_ARCACHE,
	sum_28_m_axi_gmem_ARPROT,
	sum_28_m_axi_gmem_ARQOS,
	sum_28_m_axi_gmem_ARREGION,
	sum_28_m_axi_gmem_ARUSER,
	sum_28_m_axi_gmem_RREADY,
	sum_28_m_axi_gmem_RVALID,
	sum_28_m_axi_gmem_RID,
	sum_28_m_axi_gmem_RDATA,
	sum_28_m_axi_gmem_RRESP,
	sum_28_m_axi_gmem_RLAST,
	sum_28_m_axi_gmem_RUSER,
	sum_28_m_axi_gmem_AWREADY,
	sum_28_m_axi_gmem_AWVALID,
	sum_28_m_axi_gmem_AWID,
	sum_28_m_axi_gmem_AWADDR,
	sum_28_m_axi_gmem_AWLEN,
	sum_28_m_axi_gmem_AWSIZE,
	sum_28_m_axi_gmem_AWBURST,
	sum_28_m_axi_gmem_AWLOCK,
	sum_28_m_axi_gmem_AWCACHE,
	sum_28_m_axi_gmem_AWPROT,
	sum_28_m_axi_gmem_AWQOS,
	sum_28_m_axi_gmem_AWREGION,
	sum_28_m_axi_gmem_AWUSER,
	sum_28_m_axi_gmem_WREADY,
	sum_28_m_axi_gmem_WVALID,
	sum_28_m_axi_gmem_WDATA,
	sum_28_m_axi_gmem_WSTRB,
	sum_28_m_axi_gmem_WLAST,
	sum_28_m_axi_gmem_WUSER,
	sum_28_m_axi_gmem_BREADY,
	sum_28_m_axi_gmem_BVALID,
	sum_28_m_axi_gmem_BID,
	sum_28_m_axi_gmem_BRESP,
	sum_28_m_axi_gmem_BUSER,
	sum_28_s_axi_control_ARREADY,
	sum_28_s_axi_control_ARVALID,
	sum_28_s_axi_control_ARADDR,
	sum_28_s_axi_control_RREADY,
	sum_28_s_axi_control_RVALID,
	sum_28_s_axi_control_RDATA,
	sum_28_s_axi_control_RRESP,
	sum_28_s_axi_control_AWREADY,
	sum_28_s_axi_control_AWVALID,
	sum_28_s_axi_control_AWADDR,
	sum_28_s_axi_control_WREADY,
	sum_28_s_axi_control_WVALID,
	sum_28_s_axi_control_WDATA,
	sum_28_s_axi_control_WSTRB,
	sum_28_s_axi_control_BREADY,
	sum_28_s_axi_control_BVALID,
	sum_28_s_axi_control_BRESP,
	sum_29_m_axi_gmem_ARREADY,
	sum_29_m_axi_gmem_ARVALID,
	sum_29_m_axi_gmem_ARID,
	sum_29_m_axi_gmem_ARADDR,
	sum_29_m_axi_gmem_ARLEN,
	sum_29_m_axi_gmem_ARSIZE,
	sum_29_m_axi_gmem_ARBURST,
	sum_29_m_axi_gmem_ARLOCK,
	sum_29_m_axi_gmem_ARCACHE,
	sum_29_m_axi_gmem_ARPROT,
	sum_29_m_axi_gmem_ARQOS,
	sum_29_m_axi_gmem_ARREGION,
	sum_29_m_axi_gmem_ARUSER,
	sum_29_m_axi_gmem_RREADY,
	sum_29_m_axi_gmem_RVALID,
	sum_29_m_axi_gmem_RID,
	sum_29_m_axi_gmem_RDATA,
	sum_29_m_axi_gmem_RRESP,
	sum_29_m_axi_gmem_RLAST,
	sum_29_m_axi_gmem_RUSER,
	sum_29_m_axi_gmem_AWREADY,
	sum_29_m_axi_gmem_AWVALID,
	sum_29_m_axi_gmem_AWID,
	sum_29_m_axi_gmem_AWADDR,
	sum_29_m_axi_gmem_AWLEN,
	sum_29_m_axi_gmem_AWSIZE,
	sum_29_m_axi_gmem_AWBURST,
	sum_29_m_axi_gmem_AWLOCK,
	sum_29_m_axi_gmem_AWCACHE,
	sum_29_m_axi_gmem_AWPROT,
	sum_29_m_axi_gmem_AWQOS,
	sum_29_m_axi_gmem_AWREGION,
	sum_29_m_axi_gmem_AWUSER,
	sum_29_m_axi_gmem_WREADY,
	sum_29_m_axi_gmem_WVALID,
	sum_29_m_axi_gmem_WDATA,
	sum_29_m_axi_gmem_WSTRB,
	sum_29_m_axi_gmem_WLAST,
	sum_29_m_axi_gmem_WUSER,
	sum_29_m_axi_gmem_BREADY,
	sum_29_m_axi_gmem_BVALID,
	sum_29_m_axi_gmem_BID,
	sum_29_m_axi_gmem_BRESP,
	sum_29_m_axi_gmem_BUSER,
	sum_29_s_axi_control_ARREADY,
	sum_29_s_axi_control_ARVALID,
	sum_29_s_axi_control_ARADDR,
	sum_29_s_axi_control_RREADY,
	sum_29_s_axi_control_RVALID,
	sum_29_s_axi_control_RDATA,
	sum_29_s_axi_control_RRESP,
	sum_29_s_axi_control_AWREADY,
	sum_29_s_axi_control_AWVALID,
	sum_29_s_axi_control_AWADDR,
	sum_29_s_axi_control_WREADY,
	sum_29_s_axi_control_WVALID,
	sum_29_s_axi_control_WDATA,
	sum_29_s_axi_control_WSTRB,
	sum_29_s_axi_control_BREADY,
	sum_29_s_axi_control_BVALID,
	sum_29_s_axi_control_BRESP,
	sum_30_m_axi_gmem_ARREADY,
	sum_30_m_axi_gmem_ARVALID,
	sum_30_m_axi_gmem_ARID,
	sum_30_m_axi_gmem_ARADDR,
	sum_30_m_axi_gmem_ARLEN,
	sum_30_m_axi_gmem_ARSIZE,
	sum_30_m_axi_gmem_ARBURST,
	sum_30_m_axi_gmem_ARLOCK,
	sum_30_m_axi_gmem_ARCACHE,
	sum_30_m_axi_gmem_ARPROT,
	sum_30_m_axi_gmem_ARQOS,
	sum_30_m_axi_gmem_ARREGION,
	sum_30_m_axi_gmem_ARUSER,
	sum_30_m_axi_gmem_RREADY,
	sum_30_m_axi_gmem_RVALID,
	sum_30_m_axi_gmem_RID,
	sum_30_m_axi_gmem_RDATA,
	sum_30_m_axi_gmem_RRESP,
	sum_30_m_axi_gmem_RLAST,
	sum_30_m_axi_gmem_RUSER,
	sum_30_m_axi_gmem_AWREADY,
	sum_30_m_axi_gmem_AWVALID,
	sum_30_m_axi_gmem_AWID,
	sum_30_m_axi_gmem_AWADDR,
	sum_30_m_axi_gmem_AWLEN,
	sum_30_m_axi_gmem_AWSIZE,
	sum_30_m_axi_gmem_AWBURST,
	sum_30_m_axi_gmem_AWLOCK,
	sum_30_m_axi_gmem_AWCACHE,
	sum_30_m_axi_gmem_AWPROT,
	sum_30_m_axi_gmem_AWQOS,
	sum_30_m_axi_gmem_AWREGION,
	sum_30_m_axi_gmem_AWUSER,
	sum_30_m_axi_gmem_WREADY,
	sum_30_m_axi_gmem_WVALID,
	sum_30_m_axi_gmem_WDATA,
	sum_30_m_axi_gmem_WSTRB,
	sum_30_m_axi_gmem_WLAST,
	sum_30_m_axi_gmem_WUSER,
	sum_30_m_axi_gmem_BREADY,
	sum_30_m_axi_gmem_BVALID,
	sum_30_m_axi_gmem_BID,
	sum_30_m_axi_gmem_BRESP,
	sum_30_m_axi_gmem_BUSER,
	sum_30_s_axi_control_ARREADY,
	sum_30_s_axi_control_ARVALID,
	sum_30_s_axi_control_ARADDR,
	sum_30_s_axi_control_RREADY,
	sum_30_s_axi_control_RVALID,
	sum_30_s_axi_control_RDATA,
	sum_30_s_axi_control_RRESP,
	sum_30_s_axi_control_AWREADY,
	sum_30_s_axi_control_AWVALID,
	sum_30_s_axi_control_AWADDR,
	sum_30_s_axi_control_WREADY,
	sum_30_s_axi_control_WVALID,
	sum_30_s_axi_control_WDATA,
	sum_30_s_axi_control_WSTRB,
	sum_30_s_axi_control_BREADY,
	sum_30_s_axi_control_BVALID,
	sum_30_s_axi_control_BRESP,
	sum_31_m_axi_gmem_ARREADY,
	sum_31_m_axi_gmem_ARVALID,
	sum_31_m_axi_gmem_ARID,
	sum_31_m_axi_gmem_ARADDR,
	sum_31_m_axi_gmem_ARLEN,
	sum_31_m_axi_gmem_ARSIZE,
	sum_31_m_axi_gmem_ARBURST,
	sum_31_m_axi_gmem_ARLOCK,
	sum_31_m_axi_gmem_ARCACHE,
	sum_31_m_axi_gmem_ARPROT,
	sum_31_m_axi_gmem_ARQOS,
	sum_31_m_axi_gmem_ARREGION,
	sum_31_m_axi_gmem_ARUSER,
	sum_31_m_axi_gmem_RREADY,
	sum_31_m_axi_gmem_RVALID,
	sum_31_m_axi_gmem_RID,
	sum_31_m_axi_gmem_RDATA,
	sum_31_m_axi_gmem_RRESP,
	sum_31_m_axi_gmem_RLAST,
	sum_31_m_axi_gmem_RUSER,
	sum_31_m_axi_gmem_AWREADY,
	sum_31_m_axi_gmem_AWVALID,
	sum_31_m_axi_gmem_AWID,
	sum_31_m_axi_gmem_AWADDR,
	sum_31_m_axi_gmem_AWLEN,
	sum_31_m_axi_gmem_AWSIZE,
	sum_31_m_axi_gmem_AWBURST,
	sum_31_m_axi_gmem_AWLOCK,
	sum_31_m_axi_gmem_AWCACHE,
	sum_31_m_axi_gmem_AWPROT,
	sum_31_m_axi_gmem_AWQOS,
	sum_31_m_axi_gmem_AWREGION,
	sum_31_m_axi_gmem_AWUSER,
	sum_31_m_axi_gmem_WREADY,
	sum_31_m_axi_gmem_WVALID,
	sum_31_m_axi_gmem_WDATA,
	sum_31_m_axi_gmem_WSTRB,
	sum_31_m_axi_gmem_WLAST,
	sum_31_m_axi_gmem_WUSER,
	sum_31_m_axi_gmem_BREADY,
	sum_31_m_axi_gmem_BVALID,
	sum_31_m_axi_gmem_BID,
	sum_31_m_axi_gmem_BRESP,
	sum_31_m_axi_gmem_BUSER,
	sum_31_s_axi_control_ARREADY,
	sum_31_s_axi_control_ARVALID,
	sum_31_s_axi_control_ARADDR,
	sum_31_s_axi_control_RREADY,
	sum_31_s_axi_control_RVALID,
	sum_31_s_axi_control_RDATA,
	sum_31_s_axi_control_RRESP,
	sum_31_s_axi_control_AWREADY,
	sum_31_s_axi_control_AWVALID,
	sum_31_s_axi_control_AWADDR,
	sum_31_s_axi_control_WREADY,
	sum_31_s_axi_control_WVALID,
	sum_31_s_axi_control_WDATA,
	sum_31_s_axi_control_WSTRB,
	sum_31_s_axi_control_BREADY,
	sum_31_s_axi_control_BVALID,
	sum_31_s_axi_control_BRESP,
	sum_32_m_axi_gmem_ARREADY,
	sum_32_m_axi_gmem_ARVALID,
	sum_32_m_axi_gmem_ARID,
	sum_32_m_axi_gmem_ARADDR,
	sum_32_m_axi_gmem_ARLEN,
	sum_32_m_axi_gmem_ARSIZE,
	sum_32_m_axi_gmem_ARBURST,
	sum_32_m_axi_gmem_ARLOCK,
	sum_32_m_axi_gmem_ARCACHE,
	sum_32_m_axi_gmem_ARPROT,
	sum_32_m_axi_gmem_ARQOS,
	sum_32_m_axi_gmem_ARREGION,
	sum_32_m_axi_gmem_ARUSER,
	sum_32_m_axi_gmem_RREADY,
	sum_32_m_axi_gmem_RVALID,
	sum_32_m_axi_gmem_RID,
	sum_32_m_axi_gmem_RDATA,
	sum_32_m_axi_gmem_RRESP,
	sum_32_m_axi_gmem_RLAST,
	sum_32_m_axi_gmem_RUSER,
	sum_32_m_axi_gmem_AWREADY,
	sum_32_m_axi_gmem_AWVALID,
	sum_32_m_axi_gmem_AWID,
	sum_32_m_axi_gmem_AWADDR,
	sum_32_m_axi_gmem_AWLEN,
	sum_32_m_axi_gmem_AWSIZE,
	sum_32_m_axi_gmem_AWBURST,
	sum_32_m_axi_gmem_AWLOCK,
	sum_32_m_axi_gmem_AWCACHE,
	sum_32_m_axi_gmem_AWPROT,
	sum_32_m_axi_gmem_AWQOS,
	sum_32_m_axi_gmem_AWREGION,
	sum_32_m_axi_gmem_AWUSER,
	sum_32_m_axi_gmem_WREADY,
	sum_32_m_axi_gmem_WVALID,
	sum_32_m_axi_gmem_WDATA,
	sum_32_m_axi_gmem_WSTRB,
	sum_32_m_axi_gmem_WLAST,
	sum_32_m_axi_gmem_WUSER,
	sum_32_m_axi_gmem_BREADY,
	sum_32_m_axi_gmem_BVALID,
	sum_32_m_axi_gmem_BID,
	sum_32_m_axi_gmem_BRESP,
	sum_32_m_axi_gmem_BUSER,
	sum_32_s_axi_control_ARREADY,
	sum_32_s_axi_control_ARVALID,
	sum_32_s_axi_control_ARADDR,
	sum_32_s_axi_control_RREADY,
	sum_32_s_axi_control_RVALID,
	sum_32_s_axi_control_RDATA,
	sum_32_s_axi_control_RRESP,
	sum_32_s_axi_control_AWREADY,
	sum_32_s_axi_control_AWVALID,
	sum_32_s_axi_control_AWADDR,
	sum_32_s_axi_control_WREADY,
	sum_32_s_axi_control_WVALID,
	sum_32_s_axi_control_WDATA,
	sum_32_s_axi_control_WSTRB,
	sum_32_s_axi_control_BREADY,
	sum_32_s_axi_control_BVALID,
	sum_32_s_axi_control_BRESP,
	sum_33_m_axi_gmem_ARREADY,
	sum_33_m_axi_gmem_ARVALID,
	sum_33_m_axi_gmem_ARID,
	sum_33_m_axi_gmem_ARADDR,
	sum_33_m_axi_gmem_ARLEN,
	sum_33_m_axi_gmem_ARSIZE,
	sum_33_m_axi_gmem_ARBURST,
	sum_33_m_axi_gmem_ARLOCK,
	sum_33_m_axi_gmem_ARCACHE,
	sum_33_m_axi_gmem_ARPROT,
	sum_33_m_axi_gmem_ARQOS,
	sum_33_m_axi_gmem_ARREGION,
	sum_33_m_axi_gmem_ARUSER,
	sum_33_m_axi_gmem_RREADY,
	sum_33_m_axi_gmem_RVALID,
	sum_33_m_axi_gmem_RID,
	sum_33_m_axi_gmem_RDATA,
	sum_33_m_axi_gmem_RRESP,
	sum_33_m_axi_gmem_RLAST,
	sum_33_m_axi_gmem_RUSER,
	sum_33_m_axi_gmem_AWREADY,
	sum_33_m_axi_gmem_AWVALID,
	sum_33_m_axi_gmem_AWID,
	sum_33_m_axi_gmem_AWADDR,
	sum_33_m_axi_gmem_AWLEN,
	sum_33_m_axi_gmem_AWSIZE,
	sum_33_m_axi_gmem_AWBURST,
	sum_33_m_axi_gmem_AWLOCK,
	sum_33_m_axi_gmem_AWCACHE,
	sum_33_m_axi_gmem_AWPROT,
	sum_33_m_axi_gmem_AWQOS,
	sum_33_m_axi_gmem_AWREGION,
	sum_33_m_axi_gmem_AWUSER,
	sum_33_m_axi_gmem_WREADY,
	sum_33_m_axi_gmem_WVALID,
	sum_33_m_axi_gmem_WDATA,
	sum_33_m_axi_gmem_WSTRB,
	sum_33_m_axi_gmem_WLAST,
	sum_33_m_axi_gmem_WUSER,
	sum_33_m_axi_gmem_BREADY,
	sum_33_m_axi_gmem_BVALID,
	sum_33_m_axi_gmem_BID,
	sum_33_m_axi_gmem_BRESP,
	sum_33_m_axi_gmem_BUSER,
	sum_33_s_axi_control_ARREADY,
	sum_33_s_axi_control_ARVALID,
	sum_33_s_axi_control_ARADDR,
	sum_33_s_axi_control_RREADY,
	sum_33_s_axi_control_RVALID,
	sum_33_s_axi_control_RDATA,
	sum_33_s_axi_control_RRESP,
	sum_33_s_axi_control_AWREADY,
	sum_33_s_axi_control_AWVALID,
	sum_33_s_axi_control_AWADDR,
	sum_33_s_axi_control_WREADY,
	sum_33_s_axi_control_WVALID,
	sum_33_s_axi_control_WDATA,
	sum_33_s_axi_control_WSTRB,
	sum_33_s_axi_control_BREADY,
	sum_33_s_axi_control_BVALID,
	sum_33_s_axi_control_BRESP,
	sum_34_m_axi_gmem_ARREADY,
	sum_34_m_axi_gmem_ARVALID,
	sum_34_m_axi_gmem_ARID,
	sum_34_m_axi_gmem_ARADDR,
	sum_34_m_axi_gmem_ARLEN,
	sum_34_m_axi_gmem_ARSIZE,
	sum_34_m_axi_gmem_ARBURST,
	sum_34_m_axi_gmem_ARLOCK,
	sum_34_m_axi_gmem_ARCACHE,
	sum_34_m_axi_gmem_ARPROT,
	sum_34_m_axi_gmem_ARQOS,
	sum_34_m_axi_gmem_ARREGION,
	sum_34_m_axi_gmem_ARUSER,
	sum_34_m_axi_gmem_RREADY,
	sum_34_m_axi_gmem_RVALID,
	sum_34_m_axi_gmem_RID,
	sum_34_m_axi_gmem_RDATA,
	sum_34_m_axi_gmem_RRESP,
	sum_34_m_axi_gmem_RLAST,
	sum_34_m_axi_gmem_RUSER,
	sum_34_m_axi_gmem_AWREADY,
	sum_34_m_axi_gmem_AWVALID,
	sum_34_m_axi_gmem_AWID,
	sum_34_m_axi_gmem_AWADDR,
	sum_34_m_axi_gmem_AWLEN,
	sum_34_m_axi_gmem_AWSIZE,
	sum_34_m_axi_gmem_AWBURST,
	sum_34_m_axi_gmem_AWLOCK,
	sum_34_m_axi_gmem_AWCACHE,
	sum_34_m_axi_gmem_AWPROT,
	sum_34_m_axi_gmem_AWQOS,
	sum_34_m_axi_gmem_AWREGION,
	sum_34_m_axi_gmem_AWUSER,
	sum_34_m_axi_gmem_WREADY,
	sum_34_m_axi_gmem_WVALID,
	sum_34_m_axi_gmem_WDATA,
	sum_34_m_axi_gmem_WSTRB,
	sum_34_m_axi_gmem_WLAST,
	sum_34_m_axi_gmem_WUSER,
	sum_34_m_axi_gmem_BREADY,
	sum_34_m_axi_gmem_BVALID,
	sum_34_m_axi_gmem_BID,
	sum_34_m_axi_gmem_BRESP,
	sum_34_m_axi_gmem_BUSER,
	sum_34_s_axi_control_ARREADY,
	sum_34_s_axi_control_ARVALID,
	sum_34_s_axi_control_ARADDR,
	sum_34_s_axi_control_RREADY,
	sum_34_s_axi_control_RVALID,
	sum_34_s_axi_control_RDATA,
	sum_34_s_axi_control_RRESP,
	sum_34_s_axi_control_AWREADY,
	sum_34_s_axi_control_AWVALID,
	sum_34_s_axi_control_AWADDR,
	sum_34_s_axi_control_WREADY,
	sum_34_s_axi_control_WVALID,
	sum_34_s_axi_control_WDATA,
	sum_34_s_axi_control_WSTRB,
	sum_34_s_axi_control_BREADY,
	sum_34_s_axi_control_BVALID,
	sum_34_s_axi_control_BRESP,
	sum_35_m_axi_gmem_ARREADY,
	sum_35_m_axi_gmem_ARVALID,
	sum_35_m_axi_gmem_ARID,
	sum_35_m_axi_gmem_ARADDR,
	sum_35_m_axi_gmem_ARLEN,
	sum_35_m_axi_gmem_ARSIZE,
	sum_35_m_axi_gmem_ARBURST,
	sum_35_m_axi_gmem_ARLOCK,
	sum_35_m_axi_gmem_ARCACHE,
	sum_35_m_axi_gmem_ARPROT,
	sum_35_m_axi_gmem_ARQOS,
	sum_35_m_axi_gmem_ARREGION,
	sum_35_m_axi_gmem_ARUSER,
	sum_35_m_axi_gmem_RREADY,
	sum_35_m_axi_gmem_RVALID,
	sum_35_m_axi_gmem_RID,
	sum_35_m_axi_gmem_RDATA,
	sum_35_m_axi_gmem_RRESP,
	sum_35_m_axi_gmem_RLAST,
	sum_35_m_axi_gmem_RUSER,
	sum_35_m_axi_gmem_AWREADY,
	sum_35_m_axi_gmem_AWVALID,
	sum_35_m_axi_gmem_AWID,
	sum_35_m_axi_gmem_AWADDR,
	sum_35_m_axi_gmem_AWLEN,
	sum_35_m_axi_gmem_AWSIZE,
	sum_35_m_axi_gmem_AWBURST,
	sum_35_m_axi_gmem_AWLOCK,
	sum_35_m_axi_gmem_AWCACHE,
	sum_35_m_axi_gmem_AWPROT,
	sum_35_m_axi_gmem_AWQOS,
	sum_35_m_axi_gmem_AWREGION,
	sum_35_m_axi_gmem_AWUSER,
	sum_35_m_axi_gmem_WREADY,
	sum_35_m_axi_gmem_WVALID,
	sum_35_m_axi_gmem_WDATA,
	sum_35_m_axi_gmem_WSTRB,
	sum_35_m_axi_gmem_WLAST,
	sum_35_m_axi_gmem_WUSER,
	sum_35_m_axi_gmem_BREADY,
	sum_35_m_axi_gmem_BVALID,
	sum_35_m_axi_gmem_BID,
	sum_35_m_axi_gmem_BRESP,
	sum_35_m_axi_gmem_BUSER,
	sum_35_s_axi_control_ARREADY,
	sum_35_s_axi_control_ARVALID,
	sum_35_s_axi_control_ARADDR,
	sum_35_s_axi_control_RREADY,
	sum_35_s_axi_control_RVALID,
	sum_35_s_axi_control_RDATA,
	sum_35_s_axi_control_RRESP,
	sum_35_s_axi_control_AWREADY,
	sum_35_s_axi_control_AWVALID,
	sum_35_s_axi_control_AWADDR,
	sum_35_s_axi_control_WREADY,
	sum_35_s_axi_control_WVALID,
	sum_35_s_axi_control_WDATA,
	sum_35_s_axi_control_WSTRB,
	sum_35_s_axi_control_BREADY,
	sum_35_s_axi_control_BVALID,
	sum_35_s_axi_control_BRESP,
	sum_36_m_axi_gmem_ARREADY,
	sum_36_m_axi_gmem_ARVALID,
	sum_36_m_axi_gmem_ARID,
	sum_36_m_axi_gmem_ARADDR,
	sum_36_m_axi_gmem_ARLEN,
	sum_36_m_axi_gmem_ARSIZE,
	sum_36_m_axi_gmem_ARBURST,
	sum_36_m_axi_gmem_ARLOCK,
	sum_36_m_axi_gmem_ARCACHE,
	sum_36_m_axi_gmem_ARPROT,
	sum_36_m_axi_gmem_ARQOS,
	sum_36_m_axi_gmem_ARREGION,
	sum_36_m_axi_gmem_ARUSER,
	sum_36_m_axi_gmem_RREADY,
	sum_36_m_axi_gmem_RVALID,
	sum_36_m_axi_gmem_RID,
	sum_36_m_axi_gmem_RDATA,
	sum_36_m_axi_gmem_RRESP,
	sum_36_m_axi_gmem_RLAST,
	sum_36_m_axi_gmem_RUSER,
	sum_36_m_axi_gmem_AWREADY,
	sum_36_m_axi_gmem_AWVALID,
	sum_36_m_axi_gmem_AWID,
	sum_36_m_axi_gmem_AWADDR,
	sum_36_m_axi_gmem_AWLEN,
	sum_36_m_axi_gmem_AWSIZE,
	sum_36_m_axi_gmem_AWBURST,
	sum_36_m_axi_gmem_AWLOCK,
	sum_36_m_axi_gmem_AWCACHE,
	sum_36_m_axi_gmem_AWPROT,
	sum_36_m_axi_gmem_AWQOS,
	sum_36_m_axi_gmem_AWREGION,
	sum_36_m_axi_gmem_AWUSER,
	sum_36_m_axi_gmem_WREADY,
	sum_36_m_axi_gmem_WVALID,
	sum_36_m_axi_gmem_WDATA,
	sum_36_m_axi_gmem_WSTRB,
	sum_36_m_axi_gmem_WLAST,
	sum_36_m_axi_gmem_WUSER,
	sum_36_m_axi_gmem_BREADY,
	sum_36_m_axi_gmem_BVALID,
	sum_36_m_axi_gmem_BID,
	sum_36_m_axi_gmem_BRESP,
	sum_36_m_axi_gmem_BUSER,
	sum_36_s_axi_control_ARREADY,
	sum_36_s_axi_control_ARVALID,
	sum_36_s_axi_control_ARADDR,
	sum_36_s_axi_control_RREADY,
	sum_36_s_axi_control_RVALID,
	sum_36_s_axi_control_RDATA,
	sum_36_s_axi_control_RRESP,
	sum_36_s_axi_control_AWREADY,
	sum_36_s_axi_control_AWVALID,
	sum_36_s_axi_control_AWADDR,
	sum_36_s_axi_control_WREADY,
	sum_36_s_axi_control_WVALID,
	sum_36_s_axi_control_WDATA,
	sum_36_s_axi_control_WSTRB,
	sum_36_s_axi_control_BREADY,
	sum_36_s_axi_control_BVALID,
	sum_36_s_axi_control_BRESP,
	sum_37_m_axi_gmem_ARREADY,
	sum_37_m_axi_gmem_ARVALID,
	sum_37_m_axi_gmem_ARID,
	sum_37_m_axi_gmem_ARADDR,
	sum_37_m_axi_gmem_ARLEN,
	sum_37_m_axi_gmem_ARSIZE,
	sum_37_m_axi_gmem_ARBURST,
	sum_37_m_axi_gmem_ARLOCK,
	sum_37_m_axi_gmem_ARCACHE,
	sum_37_m_axi_gmem_ARPROT,
	sum_37_m_axi_gmem_ARQOS,
	sum_37_m_axi_gmem_ARREGION,
	sum_37_m_axi_gmem_ARUSER,
	sum_37_m_axi_gmem_RREADY,
	sum_37_m_axi_gmem_RVALID,
	sum_37_m_axi_gmem_RID,
	sum_37_m_axi_gmem_RDATA,
	sum_37_m_axi_gmem_RRESP,
	sum_37_m_axi_gmem_RLAST,
	sum_37_m_axi_gmem_RUSER,
	sum_37_m_axi_gmem_AWREADY,
	sum_37_m_axi_gmem_AWVALID,
	sum_37_m_axi_gmem_AWID,
	sum_37_m_axi_gmem_AWADDR,
	sum_37_m_axi_gmem_AWLEN,
	sum_37_m_axi_gmem_AWSIZE,
	sum_37_m_axi_gmem_AWBURST,
	sum_37_m_axi_gmem_AWLOCK,
	sum_37_m_axi_gmem_AWCACHE,
	sum_37_m_axi_gmem_AWPROT,
	sum_37_m_axi_gmem_AWQOS,
	sum_37_m_axi_gmem_AWREGION,
	sum_37_m_axi_gmem_AWUSER,
	sum_37_m_axi_gmem_WREADY,
	sum_37_m_axi_gmem_WVALID,
	sum_37_m_axi_gmem_WDATA,
	sum_37_m_axi_gmem_WSTRB,
	sum_37_m_axi_gmem_WLAST,
	sum_37_m_axi_gmem_WUSER,
	sum_37_m_axi_gmem_BREADY,
	sum_37_m_axi_gmem_BVALID,
	sum_37_m_axi_gmem_BID,
	sum_37_m_axi_gmem_BRESP,
	sum_37_m_axi_gmem_BUSER,
	sum_37_s_axi_control_ARREADY,
	sum_37_s_axi_control_ARVALID,
	sum_37_s_axi_control_ARADDR,
	sum_37_s_axi_control_RREADY,
	sum_37_s_axi_control_RVALID,
	sum_37_s_axi_control_RDATA,
	sum_37_s_axi_control_RRESP,
	sum_37_s_axi_control_AWREADY,
	sum_37_s_axi_control_AWVALID,
	sum_37_s_axi_control_AWADDR,
	sum_37_s_axi_control_WREADY,
	sum_37_s_axi_control_WVALID,
	sum_37_s_axi_control_WDATA,
	sum_37_s_axi_control_WSTRB,
	sum_37_s_axi_control_BREADY,
	sum_37_s_axi_control_BVALID,
	sum_37_s_axi_control_BRESP,
	sum_38_m_axi_gmem_ARREADY,
	sum_38_m_axi_gmem_ARVALID,
	sum_38_m_axi_gmem_ARID,
	sum_38_m_axi_gmem_ARADDR,
	sum_38_m_axi_gmem_ARLEN,
	sum_38_m_axi_gmem_ARSIZE,
	sum_38_m_axi_gmem_ARBURST,
	sum_38_m_axi_gmem_ARLOCK,
	sum_38_m_axi_gmem_ARCACHE,
	sum_38_m_axi_gmem_ARPROT,
	sum_38_m_axi_gmem_ARQOS,
	sum_38_m_axi_gmem_ARREGION,
	sum_38_m_axi_gmem_ARUSER,
	sum_38_m_axi_gmem_RREADY,
	sum_38_m_axi_gmem_RVALID,
	sum_38_m_axi_gmem_RID,
	sum_38_m_axi_gmem_RDATA,
	sum_38_m_axi_gmem_RRESP,
	sum_38_m_axi_gmem_RLAST,
	sum_38_m_axi_gmem_RUSER,
	sum_38_m_axi_gmem_AWREADY,
	sum_38_m_axi_gmem_AWVALID,
	sum_38_m_axi_gmem_AWID,
	sum_38_m_axi_gmem_AWADDR,
	sum_38_m_axi_gmem_AWLEN,
	sum_38_m_axi_gmem_AWSIZE,
	sum_38_m_axi_gmem_AWBURST,
	sum_38_m_axi_gmem_AWLOCK,
	sum_38_m_axi_gmem_AWCACHE,
	sum_38_m_axi_gmem_AWPROT,
	sum_38_m_axi_gmem_AWQOS,
	sum_38_m_axi_gmem_AWREGION,
	sum_38_m_axi_gmem_AWUSER,
	sum_38_m_axi_gmem_WREADY,
	sum_38_m_axi_gmem_WVALID,
	sum_38_m_axi_gmem_WDATA,
	sum_38_m_axi_gmem_WSTRB,
	sum_38_m_axi_gmem_WLAST,
	sum_38_m_axi_gmem_WUSER,
	sum_38_m_axi_gmem_BREADY,
	sum_38_m_axi_gmem_BVALID,
	sum_38_m_axi_gmem_BID,
	sum_38_m_axi_gmem_BRESP,
	sum_38_m_axi_gmem_BUSER,
	sum_38_s_axi_control_ARREADY,
	sum_38_s_axi_control_ARVALID,
	sum_38_s_axi_control_ARADDR,
	sum_38_s_axi_control_RREADY,
	sum_38_s_axi_control_RVALID,
	sum_38_s_axi_control_RDATA,
	sum_38_s_axi_control_RRESP,
	sum_38_s_axi_control_AWREADY,
	sum_38_s_axi_control_AWVALID,
	sum_38_s_axi_control_AWADDR,
	sum_38_s_axi_control_WREADY,
	sum_38_s_axi_control_WVALID,
	sum_38_s_axi_control_WDATA,
	sum_38_s_axi_control_WSTRB,
	sum_38_s_axi_control_BREADY,
	sum_38_s_axi_control_BVALID,
	sum_38_s_axi_control_BRESP,
	sum_39_m_axi_gmem_ARREADY,
	sum_39_m_axi_gmem_ARVALID,
	sum_39_m_axi_gmem_ARID,
	sum_39_m_axi_gmem_ARADDR,
	sum_39_m_axi_gmem_ARLEN,
	sum_39_m_axi_gmem_ARSIZE,
	sum_39_m_axi_gmem_ARBURST,
	sum_39_m_axi_gmem_ARLOCK,
	sum_39_m_axi_gmem_ARCACHE,
	sum_39_m_axi_gmem_ARPROT,
	sum_39_m_axi_gmem_ARQOS,
	sum_39_m_axi_gmem_ARREGION,
	sum_39_m_axi_gmem_ARUSER,
	sum_39_m_axi_gmem_RREADY,
	sum_39_m_axi_gmem_RVALID,
	sum_39_m_axi_gmem_RID,
	sum_39_m_axi_gmem_RDATA,
	sum_39_m_axi_gmem_RRESP,
	sum_39_m_axi_gmem_RLAST,
	sum_39_m_axi_gmem_RUSER,
	sum_39_m_axi_gmem_AWREADY,
	sum_39_m_axi_gmem_AWVALID,
	sum_39_m_axi_gmem_AWID,
	sum_39_m_axi_gmem_AWADDR,
	sum_39_m_axi_gmem_AWLEN,
	sum_39_m_axi_gmem_AWSIZE,
	sum_39_m_axi_gmem_AWBURST,
	sum_39_m_axi_gmem_AWLOCK,
	sum_39_m_axi_gmem_AWCACHE,
	sum_39_m_axi_gmem_AWPROT,
	sum_39_m_axi_gmem_AWQOS,
	sum_39_m_axi_gmem_AWREGION,
	sum_39_m_axi_gmem_AWUSER,
	sum_39_m_axi_gmem_WREADY,
	sum_39_m_axi_gmem_WVALID,
	sum_39_m_axi_gmem_WDATA,
	sum_39_m_axi_gmem_WSTRB,
	sum_39_m_axi_gmem_WLAST,
	sum_39_m_axi_gmem_WUSER,
	sum_39_m_axi_gmem_BREADY,
	sum_39_m_axi_gmem_BVALID,
	sum_39_m_axi_gmem_BID,
	sum_39_m_axi_gmem_BRESP,
	sum_39_m_axi_gmem_BUSER,
	sum_39_s_axi_control_ARREADY,
	sum_39_s_axi_control_ARVALID,
	sum_39_s_axi_control_ARADDR,
	sum_39_s_axi_control_RREADY,
	sum_39_s_axi_control_RVALID,
	sum_39_s_axi_control_RDATA,
	sum_39_s_axi_control_RRESP,
	sum_39_s_axi_control_AWREADY,
	sum_39_s_axi_control_AWVALID,
	sum_39_s_axi_control_AWADDR,
	sum_39_s_axi_control_WREADY,
	sum_39_s_axi_control_WVALID,
	sum_39_s_axi_control_WDATA,
	sum_39_s_axi_control_WSTRB,
	sum_39_s_axi_control_BREADY,
	sum_39_s_axi_control_BVALID,
	sum_39_s_axi_control_BRESP,
	sum_40_m_axi_gmem_ARREADY,
	sum_40_m_axi_gmem_ARVALID,
	sum_40_m_axi_gmem_ARID,
	sum_40_m_axi_gmem_ARADDR,
	sum_40_m_axi_gmem_ARLEN,
	sum_40_m_axi_gmem_ARSIZE,
	sum_40_m_axi_gmem_ARBURST,
	sum_40_m_axi_gmem_ARLOCK,
	sum_40_m_axi_gmem_ARCACHE,
	sum_40_m_axi_gmem_ARPROT,
	sum_40_m_axi_gmem_ARQOS,
	sum_40_m_axi_gmem_ARREGION,
	sum_40_m_axi_gmem_ARUSER,
	sum_40_m_axi_gmem_RREADY,
	sum_40_m_axi_gmem_RVALID,
	sum_40_m_axi_gmem_RID,
	sum_40_m_axi_gmem_RDATA,
	sum_40_m_axi_gmem_RRESP,
	sum_40_m_axi_gmem_RLAST,
	sum_40_m_axi_gmem_RUSER,
	sum_40_m_axi_gmem_AWREADY,
	sum_40_m_axi_gmem_AWVALID,
	sum_40_m_axi_gmem_AWID,
	sum_40_m_axi_gmem_AWADDR,
	sum_40_m_axi_gmem_AWLEN,
	sum_40_m_axi_gmem_AWSIZE,
	sum_40_m_axi_gmem_AWBURST,
	sum_40_m_axi_gmem_AWLOCK,
	sum_40_m_axi_gmem_AWCACHE,
	sum_40_m_axi_gmem_AWPROT,
	sum_40_m_axi_gmem_AWQOS,
	sum_40_m_axi_gmem_AWREGION,
	sum_40_m_axi_gmem_AWUSER,
	sum_40_m_axi_gmem_WREADY,
	sum_40_m_axi_gmem_WVALID,
	sum_40_m_axi_gmem_WDATA,
	sum_40_m_axi_gmem_WSTRB,
	sum_40_m_axi_gmem_WLAST,
	sum_40_m_axi_gmem_WUSER,
	sum_40_m_axi_gmem_BREADY,
	sum_40_m_axi_gmem_BVALID,
	sum_40_m_axi_gmem_BID,
	sum_40_m_axi_gmem_BRESP,
	sum_40_m_axi_gmem_BUSER,
	sum_40_s_axi_control_ARREADY,
	sum_40_s_axi_control_ARVALID,
	sum_40_s_axi_control_ARADDR,
	sum_40_s_axi_control_RREADY,
	sum_40_s_axi_control_RVALID,
	sum_40_s_axi_control_RDATA,
	sum_40_s_axi_control_RRESP,
	sum_40_s_axi_control_AWREADY,
	sum_40_s_axi_control_AWVALID,
	sum_40_s_axi_control_AWADDR,
	sum_40_s_axi_control_WREADY,
	sum_40_s_axi_control_WVALID,
	sum_40_s_axi_control_WDATA,
	sum_40_s_axi_control_WSTRB,
	sum_40_s_axi_control_BREADY,
	sum_40_s_axi_control_BVALID,
	sum_40_s_axi_control_BRESP,
	sum_41_m_axi_gmem_ARREADY,
	sum_41_m_axi_gmem_ARVALID,
	sum_41_m_axi_gmem_ARID,
	sum_41_m_axi_gmem_ARADDR,
	sum_41_m_axi_gmem_ARLEN,
	sum_41_m_axi_gmem_ARSIZE,
	sum_41_m_axi_gmem_ARBURST,
	sum_41_m_axi_gmem_ARLOCK,
	sum_41_m_axi_gmem_ARCACHE,
	sum_41_m_axi_gmem_ARPROT,
	sum_41_m_axi_gmem_ARQOS,
	sum_41_m_axi_gmem_ARREGION,
	sum_41_m_axi_gmem_ARUSER,
	sum_41_m_axi_gmem_RREADY,
	sum_41_m_axi_gmem_RVALID,
	sum_41_m_axi_gmem_RID,
	sum_41_m_axi_gmem_RDATA,
	sum_41_m_axi_gmem_RRESP,
	sum_41_m_axi_gmem_RLAST,
	sum_41_m_axi_gmem_RUSER,
	sum_41_m_axi_gmem_AWREADY,
	sum_41_m_axi_gmem_AWVALID,
	sum_41_m_axi_gmem_AWID,
	sum_41_m_axi_gmem_AWADDR,
	sum_41_m_axi_gmem_AWLEN,
	sum_41_m_axi_gmem_AWSIZE,
	sum_41_m_axi_gmem_AWBURST,
	sum_41_m_axi_gmem_AWLOCK,
	sum_41_m_axi_gmem_AWCACHE,
	sum_41_m_axi_gmem_AWPROT,
	sum_41_m_axi_gmem_AWQOS,
	sum_41_m_axi_gmem_AWREGION,
	sum_41_m_axi_gmem_AWUSER,
	sum_41_m_axi_gmem_WREADY,
	sum_41_m_axi_gmem_WVALID,
	sum_41_m_axi_gmem_WDATA,
	sum_41_m_axi_gmem_WSTRB,
	sum_41_m_axi_gmem_WLAST,
	sum_41_m_axi_gmem_WUSER,
	sum_41_m_axi_gmem_BREADY,
	sum_41_m_axi_gmem_BVALID,
	sum_41_m_axi_gmem_BID,
	sum_41_m_axi_gmem_BRESP,
	sum_41_m_axi_gmem_BUSER,
	sum_41_s_axi_control_ARREADY,
	sum_41_s_axi_control_ARVALID,
	sum_41_s_axi_control_ARADDR,
	sum_41_s_axi_control_RREADY,
	sum_41_s_axi_control_RVALID,
	sum_41_s_axi_control_RDATA,
	sum_41_s_axi_control_RRESP,
	sum_41_s_axi_control_AWREADY,
	sum_41_s_axi_control_AWVALID,
	sum_41_s_axi_control_AWADDR,
	sum_41_s_axi_control_WREADY,
	sum_41_s_axi_control_WVALID,
	sum_41_s_axi_control_WDATA,
	sum_41_s_axi_control_WSTRB,
	sum_41_s_axi_control_BREADY,
	sum_41_s_axi_control_BVALID,
	sum_41_s_axi_control_BRESP,
	sum_42_m_axi_gmem_ARREADY,
	sum_42_m_axi_gmem_ARVALID,
	sum_42_m_axi_gmem_ARID,
	sum_42_m_axi_gmem_ARADDR,
	sum_42_m_axi_gmem_ARLEN,
	sum_42_m_axi_gmem_ARSIZE,
	sum_42_m_axi_gmem_ARBURST,
	sum_42_m_axi_gmem_ARLOCK,
	sum_42_m_axi_gmem_ARCACHE,
	sum_42_m_axi_gmem_ARPROT,
	sum_42_m_axi_gmem_ARQOS,
	sum_42_m_axi_gmem_ARREGION,
	sum_42_m_axi_gmem_ARUSER,
	sum_42_m_axi_gmem_RREADY,
	sum_42_m_axi_gmem_RVALID,
	sum_42_m_axi_gmem_RID,
	sum_42_m_axi_gmem_RDATA,
	sum_42_m_axi_gmem_RRESP,
	sum_42_m_axi_gmem_RLAST,
	sum_42_m_axi_gmem_RUSER,
	sum_42_m_axi_gmem_AWREADY,
	sum_42_m_axi_gmem_AWVALID,
	sum_42_m_axi_gmem_AWID,
	sum_42_m_axi_gmem_AWADDR,
	sum_42_m_axi_gmem_AWLEN,
	sum_42_m_axi_gmem_AWSIZE,
	sum_42_m_axi_gmem_AWBURST,
	sum_42_m_axi_gmem_AWLOCK,
	sum_42_m_axi_gmem_AWCACHE,
	sum_42_m_axi_gmem_AWPROT,
	sum_42_m_axi_gmem_AWQOS,
	sum_42_m_axi_gmem_AWREGION,
	sum_42_m_axi_gmem_AWUSER,
	sum_42_m_axi_gmem_WREADY,
	sum_42_m_axi_gmem_WVALID,
	sum_42_m_axi_gmem_WDATA,
	sum_42_m_axi_gmem_WSTRB,
	sum_42_m_axi_gmem_WLAST,
	sum_42_m_axi_gmem_WUSER,
	sum_42_m_axi_gmem_BREADY,
	sum_42_m_axi_gmem_BVALID,
	sum_42_m_axi_gmem_BID,
	sum_42_m_axi_gmem_BRESP,
	sum_42_m_axi_gmem_BUSER,
	sum_42_s_axi_control_ARREADY,
	sum_42_s_axi_control_ARVALID,
	sum_42_s_axi_control_ARADDR,
	sum_42_s_axi_control_RREADY,
	sum_42_s_axi_control_RVALID,
	sum_42_s_axi_control_RDATA,
	sum_42_s_axi_control_RRESP,
	sum_42_s_axi_control_AWREADY,
	sum_42_s_axi_control_AWVALID,
	sum_42_s_axi_control_AWADDR,
	sum_42_s_axi_control_WREADY,
	sum_42_s_axi_control_WVALID,
	sum_42_s_axi_control_WDATA,
	sum_42_s_axi_control_WSTRB,
	sum_42_s_axi_control_BREADY,
	sum_42_s_axi_control_BVALID,
	sum_42_s_axi_control_BRESP,
	sum_43_m_axi_gmem_ARREADY,
	sum_43_m_axi_gmem_ARVALID,
	sum_43_m_axi_gmem_ARID,
	sum_43_m_axi_gmem_ARADDR,
	sum_43_m_axi_gmem_ARLEN,
	sum_43_m_axi_gmem_ARSIZE,
	sum_43_m_axi_gmem_ARBURST,
	sum_43_m_axi_gmem_ARLOCK,
	sum_43_m_axi_gmem_ARCACHE,
	sum_43_m_axi_gmem_ARPROT,
	sum_43_m_axi_gmem_ARQOS,
	sum_43_m_axi_gmem_ARREGION,
	sum_43_m_axi_gmem_ARUSER,
	sum_43_m_axi_gmem_RREADY,
	sum_43_m_axi_gmem_RVALID,
	sum_43_m_axi_gmem_RID,
	sum_43_m_axi_gmem_RDATA,
	sum_43_m_axi_gmem_RRESP,
	sum_43_m_axi_gmem_RLAST,
	sum_43_m_axi_gmem_RUSER,
	sum_43_m_axi_gmem_AWREADY,
	sum_43_m_axi_gmem_AWVALID,
	sum_43_m_axi_gmem_AWID,
	sum_43_m_axi_gmem_AWADDR,
	sum_43_m_axi_gmem_AWLEN,
	sum_43_m_axi_gmem_AWSIZE,
	sum_43_m_axi_gmem_AWBURST,
	sum_43_m_axi_gmem_AWLOCK,
	sum_43_m_axi_gmem_AWCACHE,
	sum_43_m_axi_gmem_AWPROT,
	sum_43_m_axi_gmem_AWQOS,
	sum_43_m_axi_gmem_AWREGION,
	sum_43_m_axi_gmem_AWUSER,
	sum_43_m_axi_gmem_WREADY,
	sum_43_m_axi_gmem_WVALID,
	sum_43_m_axi_gmem_WDATA,
	sum_43_m_axi_gmem_WSTRB,
	sum_43_m_axi_gmem_WLAST,
	sum_43_m_axi_gmem_WUSER,
	sum_43_m_axi_gmem_BREADY,
	sum_43_m_axi_gmem_BVALID,
	sum_43_m_axi_gmem_BID,
	sum_43_m_axi_gmem_BRESP,
	sum_43_m_axi_gmem_BUSER,
	sum_43_s_axi_control_ARREADY,
	sum_43_s_axi_control_ARVALID,
	sum_43_s_axi_control_ARADDR,
	sum_43_s_axi_control_RREADY,
	sum_43_s_axi_control_RVALID,
	sum_43_s_axi_control_RDATA,
	sum_43_s_axi_control_RRESP,
	sum_43_s_axi_control_AWREADY,
	sum_43_s_axi_control_AWVALID,
	sum_43_s_axi_control_AWADDR,
	sum_43_s_axi_control_WREADY,
	sum_43_s_axi_control_WVALID,
	sum_43_s_axi_control_WDATA,
	sum_43_s_axi_control_WSTRB,
	sum_43_s_axi_control_BREADY,
	sum_43_s_axi_control_BVALID,
	sum_43_s_axi_control_BRESP,
	sum_44_m_axi_gmem_ARREADY,
	sum_44_m_axi_gmem_ARVALID,
	sum_44_m_axi_gmem_ARID,
	sum_44_m_axi_gmem_ARADDR,
	sum_44_m_axi_gmem_ARLEN,
	sum_44_m_axi_gmem_ARSIZE,
	sum_44_m_axi_gmem_ARBURST,
	sum_44_m_axi_gmem_ARLOCK,
	sum_44_m_axi_gmem_ARCACHE,
	sum_44_m_axi_gmem_ARPROT,
	sum_44_m_axi_gmem_ARQOS,
	sum_44_m_axi_gmem_ARREGION,
	sum_44_m_axi_gmem_ARUSER,
	sum_44_m_axi_gmem_RREADY,
	sum_44_m_axi_gmem_RVALID,
	sum_44_m_axi_gmem_RID,
	sum_44_m_axi_gmem_RDATA,
	sum_44_m_axi_gmem_RRESP,
	sum_44_m_axi_gmem_RLAST,
	sum_44_m_axi_gmem_RUSER,
	sum_44_m_axi_gmem_AWREADY,
	sum_44_m_axi_gmem_AWVALID,
	sum_44_m_axi_gmem_AWID,
	sum_44_m_axi_gmem_AWADDR,
	sum_44_m_axi_gmem_AWLEN,
	sum_44_m_axi_gmem_AWSIZE,
	sum_44_m_axi_gmem_AWBURST,
	sum_44_m_axi_gmem_AWLOCK,
	sum_44_m_axi_gmem_AWCACHE,
	sum_44_m_axi_gmem_AWPROT,
	sum_44_m_axi_gmem_AWQOS,
	sum_44_m_axi_gmem_AWREGION,
	sum_44_m_axi_gmem_AWUSER,
	sum_44_m_axi_gmem_WREADY,
	sum_44_m_axi_gmem_WVALID,
	sum_44_m_axi_gmem_WDATA,
	sum_44_m_axi_gmem_WSTRB,
	sum_44_m_axi_gmem_WLAST,
	sum_44_m_axi_gmem_WUSER,
	sum_44_m_axi_gmem_BREADY,
	sum_44_m_axi_gmem_BVALID,
	sum_44_m_axi_gmem_BID,
	sum_44_m_axi_gmem_BRESP,
	sum_44_m_axi_gmem_BUSER,
	sum_44_s_axi_control_ARREADY,
	sum_44_s_axi_control_ARVALID,
	sum_44_s_axi_control_ARADDR,
	sum_44_s_axi_control_RREADY,
	sum_44_s_axi_control_RVALID,
	sum_44_s_axi_control_RDATA,
	sum_44_s_axi_control_RRESP,
	sum_44_s_axi_control_AWREADY,
	sum_44_s_axi_control_AWVALID,
	sum_44_s_axi_control_AWADDR,
	sum_44_s_axi_control_WREADY,
	sum_44_s_axi_control_WVALID,
	sum_44_s_axi_control_WDATA,
	sum_44_s_axi_control_WSTRB,
	sum_44_s_axi_control_BREADY,
	sum_44_s_axi_control_BVALID,
	sum_44_s_axi_control_BRESP,
	sum_45_m_axi_gmem_ARREADY,
	sum_45_m_axi_gmem_ARVALID,
	sum_45_m_axi_gmem_ARID,
	sum_45_m_axi_gmem_ARADDR,
	sum_45_m_axi_gmem_ARLEN,
	sum_45_m_axi_gmem_ARSIZE,
	sum_45_m_axi_gmem_ARBURST,
	sum_45_m_axi_gmem_ARLOCK,
	sum_45_m_axi_gmem_ARCACHE,
	sum_45_m_axi_gmem_ARPROT,
	sum_45_m_axi_gmem_ARQOS,
	sum_45_m_axi_gmem_ARREGION,
	sum_45_m_axi_gmem_ARUSER,
	sum_45_m_axi_gmem_RREADY,
	sum_45_m_axi_gmem_RVALID,
	sum_45_m_axi_gmem_RID,
	sum_45_m_axi_gmem_RDATA,
	sum_45_m_axi_gmem_RRESP,
	sum_45_m_axi_gmem_RLAST,
	sum_45_m_axi_gmem_RUSER,
	sum_45_m_axi_gmem_AWREADY,
	sum_45_m_axi_gmem_AWVALID,
	sum_45_m_axi_gmem_AWID,
	sum_45_m_axi_gmem_AWADDR,
	sum_45_m_axi_gmem_AWLEN,
	sum_45_m_axi_gmem_AWSIZE,
	sum_45_m_axi_gmem_AWBURST,
	sum_45_m_axi_gmem_AWLOCK,
	sum_45_m_axi_gmem_AWCACHE,
	sum_45_m_axi_gmem_AWPROT,
	sum_45_m_axi_gmem_AWQOS,
	sum_45_m_axi_gmem_AWREGION,
	sum_45_m_axi_gmem_AWUSER,
	sum_45_m_axi_gmem_WREADY,
	sum_45_m_axi_gmem_WVALID,
	sum_45_m_axi_gmem_WDATA,
	sum_45_m_axi_gmem_WSTRB,
	sum_45_m_axi_gmem_WLAST,
	sum_45_m_axi_gmem_WUSER,
	sum_45_m_axi_gmem_BREADY,
	sum_45_m_axi_gmem_BVALID,
	sum_45_m_axi_gmem_BID,
	sum_45_m_axi_gmem_BRESP,
	sum_45_m_axi_gmem_BUSER,
	sum_45_s_axi_control_ARREADY,
	sum_45_s_axi_control_ARVALID,
	sum_45_s_axi_control_ARADDR,
	sum_45_s_axi_control_RREADY,
	sum_45_s_axi_control_RVALID,
	sum_45_s_axi_control_RDATA,
	sum_45_s_axi_control_RRESP,
	sum_45_s_axi_control_AWREADY,
	sum_45_s_axi_control_AWVALID,
	sum_45_s_axi_control_AWADDR,
	sum_45_s_axi_control_WREADY,
	sum_45_s_axi_control_WVALID,
	sum_45_s_axi_control_WDATA,
	sum_45_s_axi_control_WSTRB,
	sum_45_s_axi_control_BREADY,
	sum_45_s_axi_control_BVALID,
	sum_45_s_axi_control_BRESP,
	sum_46_m_axi_gmem_ARREADY,
	sum_46_m_axi_gmem_ARVALID,
	sum_46_m_axi_gmem_ARID,
	sum_46_m_axi_gmem_ARADDR,
	sum_46_m_axi_gmem_ARLEN,
	sum_46_m_axi_gmem_ARSIZE,
	sum_46_m_axi_gmem_ARBURST,
	sum_46_m_axi_gmem_ARLOCK,
	sum_46_m_axi_gmem_ARCACHE,
	sum_46_m_axi_gmem_ARPROT,
	sum_46_m_axi_gmem_ARQOS,
	sum_46_m_axi_gmem_ARREGION,
	sum_46_m_axi_gmem_ARUSER,
	sum_46_m_axi_gmem_RREADY,
	sum_46_m_axi_gmem_RVALID,
	sum_46_m_axi_gmem_RID,
	sum_46_m_axi_gmem_RDATA,
	sum_46_m_axi_gmem_RRESP,
	sum_46_m_axi_gmem_RLAST,
	sum_46_m_axi_gmem_RUSER,
	sum_46_m_axi_gmem_AWREADY,
	sum_46_m_axi_gmem_AWVALID,
	sum_46_m_axi_gmem_AWID,
	sum_46_m_axi_gmem_AWADDR,
	sum_46_m_axi_gmem_AWLEN,
	sum_46_m_axi_gmem_AWSIZE,
	sum_46_m_axi_gmem_AWBURST,
	sum_46_m_axi_gmem_AWLOCK,
	sum_46_m_axi_gmem_AWCACHE,
	sum_46_m_axi_gmem_AWPROT,
	sum_46_m_axi_gmem_AWQOS,
	sum_46_m_axi_gmem_AWREGION,
	sum_46_m_axi_gmem_AWUSER,
	sum_46_m_axi_gmem_WREADY,
	sum_46_m_axi_gmem_WVALID,
	sum_46_m_axi_gmem_WDATA,
	sum_46_m_axi_gmem_WSTRB,
	sum_46_m_axi_gmem_WLAST,
	sum_46_m_axi_gmem_WUSER,
	sum_46_m_axi_gmem_BREADY,
	sum_46_m_axi_gmem_BVALID,
	sum_46_m_axi_gmem_BID,
	sum_46_m_axi_gmem_BRESP,
	sum_46_m_axi_gmem_BUSER,
	sum_46_s_axi_control_ARREADY,
	sum_46_s_axi_control_ARVALID,
	sum_46_s_axi_control_ARADDR,
	sum_46_s_axi_control_RREADY,
	sum_46_s_axi_control_RVALID,
	sum_46_s_axi_control_RDATA,
	sum_46_s_axi_control_RRESP,
	sum_46_s_axi_control_AWREADY,
	sum_46_s_axi_control_AWVALID,
	sum_46_s_axi_control_AWADDR,
	sum_46_s_axi_control_WREADY,
	sum_46_s_axi_control_WVALID,
	sum_46_s_axi_control_WDATA,
	sum_46_s_axi_control_WSTRB,
	sum_46_s_axi_control_BREADY,
	sum_46_s_axi_control_BVALID,
	sum_46_s_axi_control_BRESP,
	sum_47_m_axi_gmem_ARREADY,
	sum_47_m_axi_gmem_ARVALID,
	sum_47_m_axi_gmem_ARID,
	sum_47_m_axi_gmem_ARADDR,
	sum_47_m_axi_gmem_ARLEN,
	sum_47_m_axi_gmem_ARSIZE,
	sum_47_m_axi_gmem_ARBURST,
	sum_47_m_axi_gmem_ARLOCK,
	sum_47_m_axi_gmem_ARCACHE,
	sum_47_m_axi_gmem_ARPROT,
	sum_47_m_axi_gmem_ARQOS,
	sum_47_m_axi_gmem_ARREGION,
	sum_47_m_axi_gmem_ARUSER,
	sum_47_m_axi_gmem_RREADY,
	sum_47_m_axi_gmem_RVALID,
	sum_47_m_axi_gmem_RID,
	sum_47_m_axi_gmem_RDATA,
	sum_47_m_axi_gmem_RRESP,
	sum_47_m_axi_gmem_RLAST,
	sum_47_m_axi_gmem_RUSER,
	sum_47_m_axi_gmem_AWREADY,
	sum_47_m_axi_gmem_AWVALID,
	sum_47_m_axi_gmem_AWID,
	sum_47_m_axi_gmem_AWADDR,
	sum_47_m_axi_gmem_AWLEN,
	sum_47_m_axi_gmem_AWSIZE,
	sum_47_m_axi_gmem_AWBURST,
	sum_47_m_axi_gmem_AWLOCK,
	sum_47_m_axi_gmem_AWCACHE,
	sum_47_m_axi_gmem_AWPROT,
	sum_47_m_axi_gmem_AWQOS,
	sum_47_m_axi_gmem_AWREGION,
	sum_47_m_axi_gmem_AWUSER,
	sum_47_m_axi_gmem_WREADY,
	sum_47_m_axi_gmem_WVALID,
	sum_47_m_axi_gmem_WDATA,
	sum_47_m_axi_gmem_WSTRB,
	sum_47_m_axi_gmem_WLAST,
	sum_47_m_axi_gmem_WUSER,
	sum_47_m_axi_gmem_BREADY,
	sum_47_m_axi_gmem_BVALID,
	sum_47_m_axi_gmem_BID,
	sum_47_m_axi_gmem_BRESP,
	sum_47_m_axi_gmem_BUSER,
	sum_47_s_axi_control_ARREADY,
	sum_47_s_axi_control_ARVALID,
	sum_47_s_axi_control_ARADDR,
	sum_47_s_axi_control_RREADY,
	sum_47_s_axi_control_RVALID,
	sum_47_s_axi_control_RDATA,
	sum_47_s_axi_control_RRESP,
	sum_47_s_axi_control_AWREADY,
	sum_47_s_axi_control_AWVALID,
	sum_47_s_axi_control_AWADDR,
	sum_47_s_axi_control_WREADY,
	sum_47_s_axi_control_WVALID,
	sum_47_s_axi_control_WDATA,
	sum_47_s_axi_control_WSTRB,
	sum_47_s_axi_control_BREADY,
	sum_47_s_axi_control_BVALID,
	sum_47_s_axi_control_BRESP,
	sum_48_m_axi_gmem_ARREADY,
	sum_48_m_axi_gmem_ARVALID,
	sum_48_m_axi_gmem_ARID,
	sum_48_m_axi_gmem_ARADDR,
	sum_48_m_axi_gmem_ARLEN,
	sum_48_m_axi_gmem_ARSIZE,
	sum_48_m_axi_gmem_ARBURST,
	sum_48_m_axi_gmem_ARLOCK,
	sum_48_m_axi_gmem_ARCACHE,
	sum_48_m_axi_gmem_ARPROT,
	sum_48_m_axi_gmem_ARQOS,
	sum_48_m_axi_gmem_ARREGION,
	sum_48_m_axi_gmem_ARUSER,
	sum_48_m_axi_gmem_RREADY,
	sum_48_m_axi_gmem_RVALID,
	sum_48_m_axi_gmem_RID,
	sum_48_m_axi_gmem_RDATA,
	sum_48_m_axi_gmem_RRESP,
	sum_48_m_axi_gmem_RLAST,
	sum_48_m_axi_gmem_RUSER,
	sum_48_m_axi_gmem_AWREADY,
	sum_48_m_axi_gmem_AWVALID,
	sum_48_m_axi_gmem_AWID,
	sum_48_m_axi_gmem_AWADDR,
	sum_48_m_axi_gmem_AWLEN,
	sum_48_m_axi_gmem_AWSIZE,
	sum_48_m_axi_gmem_AWBURST,
	sum_48_m_axi_gmem_AWLOCK,
	sum_48_m_axi_gmem_AWCACHE,
	sum_48_m_axi_gmem_AWPROT,
	sum_48_m_axi_gmem_AWQOS,
	sum_48_m_axi_gmem_AWREGION,
	sum_48_m_axi_gmem_AWUSER,
	sum_48_m_axi_gmem_WREADY,
	sum_48_m_axi_gmem_WVALID,
	sum_48_m_axi_gmem_WDATA,
	sum_48_m_axi_gmem_WSTRB,
	sum_48_m_axi_gmem_WLAST,
	sum_48_m_axi_gmem_WUSER,
	sum_48_m_axi_gmem_BREADY,
	sum_48_m_axi_gmem_BVALID,
	sum_48_m_axi_gmem_BID,
	sum_48_m_axi_gmem_BRESP,
	sum_48_m_axi_gmem_BUSER,
	sum_48_s_axi_control_ARREADY,
	sum_48_s_axi_control_ARVALID,
	sum_48_s_axi_control_ARADDR,
	sum_48_s_axi_control_RREADY,
	sum_48_s_axi_control_RVALID,
	sum_48_s_axi_control_RDATA,
	sum_48_s_axi_control_RRESP,
	sum_48_s_axi_control_AWREADY,
	sum_48_s_axi_control_AWVALID,
	sum_48_s_axi_control_AWADDR,
	sum_48_s_axi_control_WREADY,
	sum_48_s_axi_control_WVALID,
	sum_48_s_axi_control_WDATA,
	sum_48_s_axi_control_WSTRB,
	sum_48_s_axi_control_BREADY,
	sum_48_s_axi_control_BVALID,
	sum_48_s_axi_control_BRESP,
	sum_49_m_axi_gmem_ARREADY,
	sum_49_m_axi_gmem_ARVALID,
	sum_49_m_axi_gmem_ARID,
	sum_49_m_axi_gmem_ARADDR,
	sum_49_m_axi_gmem_ARLEN,
	sum_49_m_axi_gmem_ARSIZE,
	sum_49_m_axi_gmem_ARBURST,
	sum_49_m_axi_gmem_ARLOCK,
	sum_49_m_axi_gmem_ARCACHE,
	sum_49_m_axi_gmem_ARPROT,
	sum_49_m_axi_gmem_ARQOS,
	sum_49_m_axi_gmem_ARREGION,
	sum_49_m_axi_gmem_ARUSER,
	sum_49_m_axi_gmem_RREADY,
	sum_49_m_axi_gmem_RVALID,
	sum_49_m_axi_gmem_RID,
	sum_49_m_axi_gmem_RDATA,
	sum_49_m_axi_gmem_RRESP,
	sum_49_m_axi_gmem_RLAST,
	sum_49_m_axi_gmem_RUSER,
	sum_49_m_axi_gmem_AWREADY,
	sum_49_m_axi_gmem_AWVALID,
	sum_49_m_axi_gmem_AWID,
	sum_49_m_axi_gmem_AWADDR,
	sum_49_m_axi_gmem_AWLEN,
	sum_49_m_axi_gmem_AWSIZE,
	sum_49_m_axi_gmem_AWBURST,
	sum_49_m_axi_gmem_AWLOCK,
	sum_49_m_axi_gmem_AWCACHE,
	sum_49_m_axi_gmem_AWPROT,
	sum_49_m_axi_gmem_AWQOS,
	sum_49_m_axi_gmem_AWREGION,
	sum_49_m_axi_gmem_AWUSER,
	sum_49_m_axi_gmem_WREADY,
	sum_49_m_axi_gmem_WVALID,
	sum_49_m_axi_gmem_WDATA,
	sum_49_m_axi_gmem_WSTRB,
	sum_49_m_axi_gmem_WLAST,
	sum_49_m_axi_gmem_WUSER,
	sum_49_m_axi_gmem_BREADY,
	sum_49_m_axi_gmem_BVALID,
	sum_49_m_axi_gmem_BID,
	sum_49_m_axi_gmem_BRESP,
	sum_49_m_axi_gmem_BUSER,
	sum_49_s_axi_control_ARREADY,
	sum_49_s_axi_control_ARVALID,
	sum_49_s_axi_control_ARADDR,
	sum_49_s_axi_control_RREADY,
	sum_49_s_axi_control_RVALID,
	sum_49_s_axi_control_RDATA,
	sum_49_s_axi_control_RRESP,
	sum_49_s_axi_control_AWREADY,
	sum_49_s_axi_control_AWVALID,
	sum_49_s_axi_control_AWADDR,
	sum_49_s_axi_control_WREADY,
	sum_49_s_axi_control_WVALID,
	sum_49_s_axi_control_WDATA,
	sum_49_s_axi_control_WSTRB,
	sum_49_s_axi_control_BREADY,
	sum_49_s_axi_control_BVALID,
	sum_49_s_axi_control_BRESP,
	sum_50_m_axi_gmem_ARREADY,
	sum_50_m_axi_gmem_ARVALID,
	sum_50_m_axi_gmem_ARID,
	sum_50_m_axi_gmem_ARADDR,
	sum_50_m_axi_gmem_ARLEN,
	sum_50_m_axi_gmem_ARSIZE,
	sum_50_m_axi_gmem_ARBURST,
	sum_50_m_axi_gmem_ARLOCK,
	sum_50_m_axi_gmem_ARCACHE,
	sum_50_m_axi_gmem_ARPROT,
	sum_50_m_axi_gmem_ARQOS,
	sum_50_m_axi_gmem_ARREGION,
	sum_50_m_axi_gmem_ARUSER,
	sum_50_m_axi_gmem_RREADY,
	sum_50_m_axi_gmem_RVALID,
	sum_50_m_axi_gmem_RID,
	sum_50_m_axi_gmem_RDATA,
	sum_50_m_axi_gmem_RRESP,
	sum_50_m_axi_gmem_RLAST,
	sum_50_m_axi_gmem_RUSER,
	sum_50_m_axi_gmem_AWREADY,
	sum_50_m_axi_gmem_AWVALID,
	sum_50_m_axi_gmem_AWID,
	sum_50_m_axi_gmem_AWADDR,
	sum_50_m_axi_gmem_AWLEN,
	sum_50_m_axi_gmem_AWSIZE,
	sum_50_m_axi_gmem_AWBURST,
	sum_50_m_axi_gmem_AWLOCK,
	sum_50_m_axi_gmem_AWCACHE,
	sum_50_m_axi_gmem_AWPROT,
	sum_50_m_axi_gmem_AWQOS,
	sum_50_m_axi_gmem_AWREGION,
	sum_50_m_axi_gmem_AWUSER,
	sum_50_m_axi_gmem_WREADY,
	sum_50_m_axi_gmem_WVALID,
	sum_50_m_axi_gmem_WDATA,
	sum_50_m_axi_gmem_WSTRB,
	sum_50_m_axi_gmem_WLAST,
	sum_50_m_axi_gmem_WUSER,
	sum_50_m_axi_gmem_BREADY,
	sum_50_m_axi_gmem_BVALID,
	sum_50_m_axi_gmem_BID,
	sum_50_m_axi_gmem_BRESP,
	sum_50_m_axi_gmem_BUSER,
	sum_50_s_axi_control_ARREADY,
	sum_50_s_axi_control_ARVALID,
	sum_50_s_axi_control_ARADDR,
	sum_50_s_axi_control_RREADY,
	sum_50_s_axi_control_RVALID,
	sum_50_s_axi_control_RDATA,
	sum_50_s_axi_control_RRESP,
	sum_50_s_axi_control_AWREADY,
	sum_50_s_axi_control_AWVALID,
	sum_50_s_axi_control_AWADDR,
	sum_50_s_axi_control_WREADY,
	sum_50_s_axi_control_WVALID,
	sum_50_s_axi_control_WDATA,
	sum_50_s_axi_control_WSTRB,
	sum_50_s_axi_control_BREADY,
	sum_50_s_axi_control_BVALID,
	sum_50_s_axi_control_BRESP,
	sum_51_m_axi_gmem_ARREADY,
	sum_51_m_axi_gmem_ARVALID,
	sum_51_m_axi_gmem_ARID,
	sum_51_m_axi_gmem_ARADDR,
	sum_51_m_axi_gmem_ARLEN,
	sum_51_m_axi_gmem_ARSIZE,
	sum_51_m_axi_gmem_ARBURST,
	sum_51_m_axi_gmem_ARLOCK,
	sum_51_m_axi_gmem_ARCACHE,
	sum_51_m_axi_gmem_ARPROT,
	sum_51_m_axi_gmem_ARQOS,
	sum_51_m_axi_gmem_ARREGION,
	sum_51_m_axi_gmem_ARUSER,
	sum_51_m_axi_gmem_RREADY,
	sum_51_m_axi_gmem_RVALID,
	sum_51_m_axi_gmem_RID,
	sum_51_m_axi_gmem_RDATA,
	sum_51_m_axi_gmem_RRESP,
	sum_51_m_axi_gmem_RLAST,
	sum_51_m_axi_gmem_RUSER,
	sum_51_m_axi_gmem_AWREADY,
	sum_51_m_axi_gmem_AWVALID,
	sum_51_m_axi_gmem_AWID,
	sum_51_m_axi_gmem_AWADDR,
	sum_51_m_axi_gmem_AWLEN,
	sum_51_m_axi_gmem_AWSIZE,
	sum_51_m_axi_gmem_AWBURST,
	sum_51_m_axi_gmem_AWLOCK,
	sum_51_m_axi_gmem_AWCACHE,
	sum_51_m_axi_gmem_AWPROT,
	sum_51_m_axi_gmem_AWQOS,
	sum_51_m_axi_gmem_AWREGION,
	sum_51_m_axi_gmem_AWUSER,
	sum_51_m_axi_gmem_WREADY,
	sum_51_m_axi_gmem_WVALID,
	sum_51_m_axi_gmem_WDATA,
	sum_51_m_axi_gmem_WSTRB,
	sum_51_m_axi_gmem_WLAST,
	sum_51_m_axi_gmem_WUSER,
	sum_51_m_axi_gmem_BREADY,
	sum_51_m_axi_gmem_BVALID,
	sum_51_m_axi_gmem_BID,
	sum_51_m_axi_gmem_BRESP,
	sum_51_m_axi_gmem_BUSER,
	sum_51_s_axi_control_ARREADY,
	sum_51_s_axi_control_ARVALID,
	sum_51_s_axi_control_ARADDR,
	sum_51_s_axi_control_RREADY,
	sum_51_s_axi_control_RVALID,
	sum_51_s_axi_control_RDATA,
	sum_51_s_axi_control_RRESP,
	sum_51_s_axi_control_AWREADY,
	sum_51_s_axi_control_AWVALID,
	sum_51_s_axi_control_AWADDR,
	sum_51_s_axi_control_WREADY,
	sum_51_s_axi_control_WVALID,
	sum_51_s_axi_control_WDATA,
	sum_51_s_axi_control_WSTRB,
	sum_51_s_axi_control_BREADY,
	sum_51_s_axi_control_BVALID,
	sum_51_s_axi_control_BRESP,
	sum_52_m_axi_gmem_ARREADY,
	sum_52_m_axi_gmem_ARVALID,
	sum_52_m_axi_gmem_ARID,
	sum_52_m_axi_gmem_ARADDR,
	sum_52_m_axi_gmem_ARLEN,
	sum_52_m_axi_gmem_ARSIZE,
	sum_52_m_axi_gmem_ARBURST,
	sum_52_m_axi_gmem_ARLOCK,
	sum_52_m_axi_gmem_ARCACHE,
	sum_52_m_axi_gmem_ARPROT,
	sum_52_m_axi_gmem_ARQOS,
	sum_52_m_axi_gmem_ARREGION,
	sum_52_m_axi_gmem_ARUSER,
	sum_52_m_axi_gmem_RREADY,
	sum_52_m_axi_gmem_RVALID,
	sum_52_m_axi_gmem_RID,
	sum_52_m_axi_gmem_RDATA,
	sum_52_m_axi_gmem_RRESP,
	sum_52_m_axi_gmem_RLAST,
	sum_52_m_axi_gmem_RUSER,
	sum_52_m_axi_gmem_AWREADY,
	sum_52_m_axi_gmem_AWVALID,
	sum_52_m_axi_gmem_AWID,
	sum_52_m_axi_gmem_AWADDR,
	sum_52_m_axi_gmem_AWLEN,
	sum_52_m_axi_gmem_AWSIZE,
	sum_52_m_axi_gmem_AWBURST,
	sum_52_m_axi_gmem_AWLOCK,
	sum_52_m_axi_gmem_AWCACHE,
	sum_52_m_axi_gmem_AWPROT,
	sum_52_m_axi_gmem_AWQOS,
	sum_52_m_axi_gmem_AWREGION,
	sum_52_m_axi_gmem_AWUSER,
	sum_52_m_axi_gmem_WREADY,
	sum_52_m_axi_gmem_WVALID,
	sum_52_m_axi_gmem_WDATA,
	sum_52_m_axi_gmem_WSTRB,
	sum_52_m_axi_gmem_WLAST,
	sum_52_m_axi_gmem_WUSER,
	sum_52_m_axi_gmem_BREADY,
	sum_52_m_axi_gmem_BVALID,
	sum_52_m_axi_gmem_BID,
	sum_52_m_axi_gmem_BRESP,
	sum_52_m_axi_gmem_BUSER,
	sum_52_s_axi_control_ARREADY,
	sum_52_s_axi_control_ARVALID,
	sum_52_s_axi_control_ARADDR,
	sum_52_s_axi_control_RREADY,
	sum_52_s_axi_control_RVALID,
	sum_52_s_axi_control_RDATA,
	sum_52_s_axi_control_RRESP,
	sum_52_s_axi_control_AWREADY,
	sum_52_s_axi_control_AWVALID,
	sum_52_s_axi_control_AWADDR,
	sum_52_s_axi_control_WREADY,
	sum_52_s_axi_control_WVALID,
	sum_52_s_axi_control_WDATA,
	sum_52_s_axi_control_WSTRB,
	sum_52_s_axi_control_BREADY,
	sum_52_s_axi_control_BVALID,
	sum_52_s_axi_control_BRESP,
	sum_53_m_axi_gmem_ARREADY,
	sum_53_m_axi_gmem_ARVALID,
	sum_53_m_axi_gmem_ARID,
	sum_53_m_axi_gmem_ARADDR,
	sum_53_m_axi_gmem_ARLEN,
	sum_53_m_axi_gmem_ARSIZE,
	sum_53_m_axi_gmem_ARBURST,
	sum_53_m_axi_gmem_ARLOCK,
	sum_53_m_axi_gmem_ARCACHE,
	sum_53_m_axi_gmem_ARPROT,
	sum_53_m_axi_gmem_ARQOS,
	sum_53_m_axi_gmem_ARREGION,
	sum_53_m_axi_gmem_ARUSER,
	sum_53_m_axi_gmem_RREADY,
	sum_53_m_axi_gmem_RVALID,
	sum_53_m_axi_gmem_RID,
	sum_53_m_axi_gmem_RDATA,
	sum_53_m_axi_gmem_RRESP,
	sum_53_m_axi_gmem_RLAST,
	sum_53_m_axi_gmem_RUSER,
	sum_53_m_axi_gmem_AWREADY,
	sum_53_m_axi_gmem_AWVALID,
	sum_53_m_axi_gmem_AWID,
	sum_53_m_axi_gmem_AWADDR,
	sum_53_m_axi_gmem_AWLEN,
	sum_53_m_axi_gmem_AWSIZE,
	sum_53_m_axi_gmem_AWBURST,
	sum_53_m_axi_gmem_AWLOCK,
	sum_53_m_axi_gmem_AWCACHE,
	sum_53_m_axi_gmem_AWPROT,
	sum_53_m_axi_gmem_AWQOS,
	sum_53_m_axi_gmem_AWREGION,
	sum_53_m_axi_gmem_AWUSER,
	sum_53_m_axi_gmem_WREADY,
	sum_53_m_axi_gmem_WVALID,
	sum_53_m_axi_gmem_WDATA,
	sum_53_m_axi_gmem_WSTRB,
	sum_53_m_axi_gmem_WLAST,
	sum_53_m_axi_gmem_WUSER,
	sum_53_m_axi_gmem_BREADY,
	sum_53_m_axi_gmem_BVALID,
	sum_53_m_axi_gmem_BID,
	sum_53_m_axi_gmem_BRESP,
	sum_53_m_axi_gmem_BUSER,
	sum_53_s_axi_control_ARREADY,
	sum_53_s_axi_control_ARVALID,
	sum_53_s_axi_control_ARADDR,
	sum_53_s_axi_control_RREADY,
	sum_53_s_axi_control_RVALID,
	sum_53_s_axi_control_RDATA,
	sum_53_s_axi_control_RRESP,
	sum_53_s_axi_control_AWREADY,
	sum_53_s_axi_control_AWVALID,
	sum_53_s_axi_control_AWADDR,
	sum_53_s_axi_control_WREADY,
	sum_53_s_axi_control_WVALID,
	sum_53_s_axi_control_WDATA,
	sum_53_s_axi_control_WSTRB,
	sum_53_s_axi_control_BREADY,
	sum_53_s_axi_control_BVALID,
	sum_53_s_axi_control_BRESP,
	sum_54_m_axi_gmem_ARREADY,
	sum_54_m_axi_gmem_ARVALID,
	sum_54_m_axi_gmem_ARID,
	sum_54_m_axi_gmem_ARADDR,
	sum_54_m_axi_gmem_ARLEN,
	sum_54_m_axi_gmem_ARSIZE,
	sum_54_m_axi_gmem_ARBURST,
	sum_54_m_axi_gmem_ARLOCK,
	sum_54_m_axi_gmem_ARCACHE,
	sum_54_m_axi_gmem_ARPROT,
	sum_54_m_axi_gmem_ARQOS,
	sum_54_m_axi_gmem_ARREGION,
	sum_54_m_axi_gmem_ARUSER,
	sum_54_m_axi_gmem_RREADY,
	sum_54_m_axi_gmem_RVALID,
	sum_54_m_axi_gmem_RID,
	sum_54_m_axi_gmem_RDATA,
	sum_54_m_axi_gmem_RRESP,
	sum_54_m_axi_gmem_RLAST,
	sum_54_m_axi_gmem_RUSER,
	sum_54_m_axi_gmem_AWREADY,
	sum_54_m_axi_gmem_AWVALID,
	sum_54_m_axi_gmem_AWID,
	sum_54_m_axi_gmem_AWADDR,
	sum_54_m_axi_gmem_AWLEN,
	sum_54_m_axi_gmem_AWSIZE,
	sum_54_m_axi_gmem_AWBURST,
	sum_54_m_axi_gmem_AWLOCK,
	sum_54_m_axi_gmem_AWCACHE,
	sum_54_m_axi_gmem_AWPROT,
	sum_54_m_axi_gmem_AWQOS,
	sum_54_m_axi_gmem_AWREGION,
	sum_54_m_axi_gmem_AWUSER,
	sum_54_m_axi_gmem_WREADY,
	sum_54_m_axi_gmem_WVALID,
	sum_54_m_axi_gmem_WDATA,
	sum_54_m_axi_gmem_WSTRB,
	sum_54_m_axi_gmem_WLAST,
	sum_54_m_axi_gmem_WUSER,
	sum_54_m_axi_gmem_BREADY,
	sum_54_m_axi_gmem_BVALID,
	sum_54_m_axi_gmem_BID,
	sum_54_m_axi_gmem_BRESP,
	sum_54_m_axi_gmem_BUSER,
	sum_54_s_axi_control_ARREADY,
	sum_54_s_axi_control_ARVALID,
	sum_54_s_axi_control_ARADDR,
	sum_54_s_axi_control_RREADY,
	sum_54_s_axi_control_RVALID,
	sum_54_s_axi_control_RDATA,
	sum_54_s_axi_control_RRESP,
	sum_54_s_axi_control_AWREADY,
	sum_54_s_axi_control_AWVALID,
	sum_54_s_axi_control_AWADDR,
	sum_54_s_axi_control_WREADY,
	sum_54_s_axi_control_WVALID,
	sum_54_s_axi_control_WDATA,
	sum_54_s_axi_control_WSTRB,
	sum_54_s_axi_control_BREADY,
	sum_54_s_axi_control_BVALID,
	sum_54_s_axi_control_BRESP,
	sum_55_m_axi_gmem_ARREADY,
	sum_55_m_axi_gmem_ARVALID,
	sum_55_m_axi_gmem_ARID,
	sum_55_m_axi_gmem_ARADDR,
	sum_55_m_axi_gmem_ARLEN,
	sum_55_m_axi_gmem_ARSIZE,
	sum_55_m_axi_gmem_ARBURST,
	sum_55_m_axi_gmem_ARLOCK,
	sum_55_m_axi_gmem_ARCACHE,
	sum_55_m_axi_gmem_ARPROT,
	sum_55_m_axi_gmem_ARQOS,
	sum_55_m_axi_gmem_ARREGION,
	sum_55_m_axi_gmem_ARUSER,
	sum_55_m_axi_gmem_RREADY,
	sum_55_m_axi_gmem_RVALID,
	sum_55_m_axi_gmem_RID,
	sum_55_m_axi_gmem_RDATA,
	sum_55_m_axi_gmem_RRESP,
	sum_55_m_axi_gmem_RLAST,
	sum_55_m_axi_gmem_RUSER,
	sum_55_m_axi_gmem_AWREADY,
	sum_55_m_axi_gmem_AWVALID,
	sum_55_m_axi_gmem_AWID,
	sum_55_m_axi_gmem_AWADDR,
	sum_55_m_axi_gmem_AWLEN,
	sum_55_m_axi_gmem_AWSIZE,
	sum_55_m_axi_gmem_AWBURST,
	sum_55_m_axi_gmem_AWLOCK,
	sum_55_m_axi_gmem_AWCACHE,
	sum_55_m_axi_gmem_AWPROT,
	sum_55_m_axi_gmem_AWQOS,
	sum_55_m_axi_gmem_AWREGION,
	sum_55_m_axi_gmem_AWUSER,
	sum_55_m_axi_gmem_WREADY,
	sum_55_m_axi_gmem_WVALID,
	sum_55_m_axi_gmem_WDATA,
	sum_55_m_axi_gmem_WSTRB,
	sum_55_m_axi_gmem_WLAST,
	sum_55_m_axi_gmem_WUSER,
	sum_55_m_axi_gmem_BREADY,
	sum_55_m_axi_gmem_BVALID,
	sum_55_m_axi_gmem_BID,
	sum_55_m_axi_gmem_BRESP,
	sum_55_m_axi_gmem_BUSER,
	sum_55_s_axi_control_ARREADY,
	sum_55_s_axi_control_ARVALID,
	sum_55_s_axi_control_ARADDR,
	sum_55_s_axi_control_RREADY,
	sum_55_s_axi_control_RVALID,
	sum_55_s_axi_control_RDATA,
	sum_55_s_axi_control_RRESP,
	sum_55_s_axi_control_AWREADY,
	sum_55_s_axi_control_AWVALID,
	sum_55_s_axi_control_AWADDR,
	sum_55_s_axi_control_WREADY,
	sum_55_s_axi_control_WVALID,
	sum_55_s_axi_control_WDATA,
	sum_55_s_axi_control_WSTRB,
	sum_55_s_axi_control_BREADY,
	sum_55_s_axi_control_BVALID,
	sum_55_s_axi_control_BRESP,
	sum_56_m_axi_gmem_ARREADY,
	sum_56_m_axi_gmem_ARVALID,
	sum_56_m_axi_gmem_ARID,
	sum_56_m_axi_gmem_ARADDR,
	sum_56_m_axi_gmem_ARLEN,
	sum_56_m_axi_gmem_ARSIZE,
	sum_56_m_axi_gmem_ARBURST,
	sum_56_m_axi_gmem_ARLOCK,
	sum_56_m_axi_gmem_ARCACHE,
	sum_56_m_axi_gmem_ARPROT,
	sum_56_m_axi_gmem_ARQOS,
	sum_56_m_axi_gmem_ARREGION,
	sum_56_m_axi_gmem_ARUSER,
	sum_56_m_axi_gmem_RREADY,
	sum_56_m_axi_gmem_RVALID,
	sum_56_m_axi_gmem_RID,
	sum_56_m_axi_gmem_RDATA,
	sum_56_m_axi_gmem_RRESP,
	sum_56_m_axi_gmem_RLAST,
	sum_56_m_axi_gmem_RUSER,
	sum_56_m_axi_gmem_AWREADY,
	sum_56_m_axi_gmem_AWVALID,
	sum_56_m_axi_gmem_AWID,
	sum_56_m_axi_gmem_AWADDR,
	sum_56_m_axi_gmem_AWLEN,
	sum_56_m_axi_gmem_AWSIZE,
	sum_56_m_axi_gmem_AWBURST,
	sum_56_m_axi_gmem_AWLOCK,
	sum_56_m_axi_gmem_AWCACHE,
	sum_56_m_axi_gmem_AWPROT,
	sum_56_m_axi_gmem_AWQOS,
	sum_56_m_axi_gmem_AWREGION,
	sum_56_m_axi_gmem_AWUSER,
	sum_56_m_axi_gmem_WREADY,
	sum_56_m_axi_gmem_WVALID,
	sum_56_m_axi_gmem_WDATA,
	sum_56_m_axi_gmem_WSTRB,
	sum_56_m_axi_gmem_WLAST,
	sum_56_m_axi_gmem_WUSER,
	sum_56_m_axi_gmem_BREADY,
	sum_56_m_axi_gmem_BVALID,
	sum_56_m_axi_gmem_BID,
	sum_56_m_axi_gmem_BRESP,
	sum_56_m_axi_gmem_BUSER,
	sum_56_s_axi_control_ARREADY,
	sum_56_s_axi_control_ARVALID,
	sum_56_s_axi_control_ARADDR,
	sum_56_s_axi_control_RREADY,
	sum_56_s_axi_control_RVALID,
	sum_56_s_axi_control_RDATA,
	sum_56_s_axi_control_RRESP,
	sum_56_s_axi_control_AWREADY,
	sum_56_s_axi_control_AWVALID,
	sum_56_s_axi_control_AWADDR,
	sum_56_s_axi_control_WREADY,
	sum_56_s_axi_control_WVALID,
	sum_56_s_axi_control_WDATA,
	sum_56_s_axi_control_WSTRB,
	sum_56_s_axi_control_BREADY,
	sum_56_s_axi_control_BVALID,
	sum_56_s_axi_control_BRESP,
	sum_57_m_axi_gmem_ARREADY,
	sum_57_m_axi_gmem_ARVALID,
	sum_57_m_axi_gmem_ARID,
	sum_57_m_axi_gmem_ARADDR,
	sum_57_m_axi_gmem_ARLEN,
	sum_57_m_axi_gmem_ARSIZE,
	sum_57_m_axi_gmem_ARBURST,
	sum_57_m_axi_gmem_ARLOCK,
	sum_57_m_axi_gmem_ARCACHE,
	sum_57_m_axi_gmem_ARPROT,
	sum_57_m_axi_gmem_ARQOS,
	sum_57_m_axi_gmem_ARREGION,
	sum_57_m_axi_gmem_ARUSER,
	sum_57_m_axi_gmem_RREADY,
	sum_57_m_axi_gmem_RVALID,
	sum_57_m_axi_gmem_RID,
	sum_57_m_axi_gmem_RDATA,
	sum_57_m_axi_gmem_RRESP,
	sum_57_m_axi_gmem_RLAST,
	sum_57_m_axi_gmem_RUSER,
	sum_57_m_axi_gmem_AWREADY,
	sum_57_m_axi_gmem_AWVALID,
	sum_57_m_axi_gmem_AWID,
	sum_57_m_axi_gmem_AWADDR,
	sum_57_m_axi_gmem_AWLEN,
	sum_57_m_axi_gmem_AWSIZE,
	sum_57_m_axi_gmem_AWBURST,
	sum_57_m_axi_gmem_AWLOCK,
	sum_57_m_axi_gmem_AWCACHE,
	sum_57_m_axi_gmem_AWPROT,
	sum_57_m_axi_gmem_AWQOS,
	sum_57_m_axi_gmem_AWREGION,
	sum_57_m_axi_gmem_AWUSER,
	sum_57_m_axi_gmem_WREADY,
	sum_57_m_axi_gmem_WVALID,
	sum_57_m_axi_gmem_WDATA,
	sum_57_m_axi_gmem_WSTRB,
	sum_57_m_axi_gmem_WLAST,
	sum_57_m_axi_gmem_WUSER,
	sum_57_m_axi_gmem_BREADY,
	sum_57_m_axi_gmem_BVALID,
	sum_57_m_axi_gmem_BID,
	sum_57_m_axi_gmem_BRESP,
	sum_57_m_axi_gmem_BUSER,
	sum_57_s_axi_control_ARREADY,
	sum_57_s_axi_control_ARVALID,
	sum_57_s_axi_control_ARADDR,
	sum_57_s_axi_control_RREADY,
	sum_57_s_axi_control_RVALID,
	sum_57_s_axi_control_RDATA,
	sum_57_s_axi_control_RRESP,
	sum_57_s_axi_control_AWREADY,
	sum_57_s_axi_control_AWVALID,
	sum_57_s_axi_control_AWADDR,
	sum_57_s_axi_control_WREADY,
	sum_57_s_axi_control_WVALID,
	sum_57_s_axi_control_WDATA,
	sum_57_s_axi_control_WSTRB,
	sum_57_s_axi_control_BREADY,
	sum_57_s_axi_control_BVALID,
	sum_57_s_axi_control_BRESP,
	sum_58_m_axi_gmem_ARREADY,
	sum_58_m_axi_gmem_ARVALID,
	sum_58_m_axi_gmem_ARID,
	sum_58_m_axi_gmem_ARADDR,
	sum_58_m_axi_gmem_ARLEN,
	sum_58_m_axi_gmem_ARSIZE,
	sum_58_m_axi_gmem_ARBURST,
	sum_58_m_axi_gmem_ARLOCK,
	sum_58_m_axi_gmem_ARCACHE,
	sum_58_m_axi_gmem_ARPROT,
	sum_58_m_axi_gmem_ARQOS,
	sum_58_m_axi_gmem_ARREGION,
	sum_58_m_axi_gmem_ARUSER,
	sum_58_m_axi_gmem_RREADY,
	sum_58_m_axi_gmem_RVALID,
	sum_58_m_axi_gmem_RID,
	sum_58_m_axi_gmem_RDATA,
	sum_58_m_axi_gmem_RRESP,
	sum_58_m_axi_gmem_RLAST,
	sum_58_m_axi_gmem_RUSER,
	sum_58_m_axi_gmem_AWREADY,
	sum_58_m_axi_gmem_AWVALID,
	sum_58_m_axi_gmem_AWID,
	sum_58_m_axi_gmem_AWADDR,
	sum_58_m_axi_gmem_AWLEN,
	sum_58_m_axi_gmem_AWSIZE,
	sum_58_m_axi_gmem_AWBURST,
	sum_58_m_axi_gmem_AWLOCK,
	sum_58_m_axi_gmem_AWCACHE,
	sum_58_m_axi_gmem_AWPROT,
	sum_58_m_axi_gmem_AWQOS,
	sum_58_m_axi_gmem_AWREGION,
	sum_58_m_axi_gmem_AWUSER,
	sum_58_m_axi_gmem_WREADY,
	sum_58_m_axi_gmem_WVALID,
	sum_58_m_axi_gmem_WDATA,
	sum_58_m_axi_gmem_WSTRB,
	sum_58_m_axi_gmem_WLAST,
	sum_58_m_axi_gmem_WUSER,
	sum_58_m_axi_gmem_BREADY,
	sum_58_m_axi_gmem_BVALID,
	sum_58_m_axi_gmem_BID,
	sum_58_m_axi_gmem_BRESP,
	sum_58_m_axi_gmem_BUSER,
	sum_58_s_axi_control_ARREADY,
	sum_58_s_axi_control_ARVALID,
	sum_58_s_axi_control_ARADDR,
	sum_58_s_axi_control_RREADY,
	sum_58_s_axi_control_RVALID,
	sum_58_s_axi_control_RDATA,
	sum_58_s_axi_control_RRESP,
	sum_58_s_axi_control_AWREADY,
	sum_58_s_axi_control_AWVALID,
	sum_58_s_axi_control_AWADDR,
	sum_58_s_axi_control_WREADY,
	sum_58_s_axi_control_WVALID,
	sum_58_s_axi_control_WDATA,
	sum_58_s_axi_control_WSTRB,
	sum_58_s_axi_control_BREADY,
	sum_58_s_axi_control_BVALID,
	sum_58_s_axi_control_BRESP,
	sum_59_m_axi_gmem_ARREADY,
	sum_59_m_axi_gmem_ARVALID,
	sum_59_m_axi_gmem_ARID,
	sum_59_m_axi_gmem_ARADDR,
	sum_59_m_axi_gmem_ARLEN,
	sum_59_m_axi_gmem_ARSIZE,
	sum_59_m_axi_gmem_ARBURST,
	sum_59_m_axi_gmem_ARLOCK,
	sum_59_m_axi_gmem_ARCACHE,
	sum_59_m_axi_gmem_ARPROT,
	sum_59_m_axi_gmem_ARQOS,
	sum_59_m_axi_gmem_ARREGION,
	sum_59_m_axi_gmem_ARUSER,
	sum_59_m_axi_gmem_RREADY,
	sum_59_m_axi_gmem_RVALID,
	sum_59_m_axi_gmem_RID,
	sum_59_m_axi_gmem_RDATA,
	sum_59_m_axi_gmem_RRESP,
	sum_59_m_axi_gmem_RLAST,
	sum_59_m_axi_gmem_RUSER,
	sum_59_m_axi_gmem_AWREADY,
	sum_59_m_axi_gmem_AWVALID,
	sum_59_m_axi_gmem_AWID,
	sum_59_m_axi_gmem_AWADDR,
	sum_59_m_axi_gmem_AWLEN,
	sum_59_m_axi_gmem_AWSIZE,
	sum_59_m_axi_gmem_AWBURST,
	sum_59_m_axi_gmem_AWLOCK,
	sum_59_m_axi_gmem_AWCACHE,
	sum_59_m_axi_gmem_AWPROT,
	sum_59_m_axi_gmem_AWQOS,
	sum_59_m_axi_gmem_AWREGION,
	sum_59_m_axi_gmem_AWUSER,
	sum_59_m_axi_gmem_WREADY,
	sum_59_m_axi_gmem_WVALID,
	sum_59_m_axi_gmem_WDATA,
	sum_59_m_axi_gmem_WSTRB,
	sum_59_m_axi_gmem_WLAST,
	sum_59_m_axi_gmem_WUSER,
	sum_59_m_axi_gmem_BREADY,
	sum_59_m_axi_gmem_BVALID,
	sum_59_m_axi_gmem_BID,
	sum_59_m_axi_gmem_BRESP,
	sum_59_m_axi_gmem_BUSER,
	sum_59_s_axi_control_ARREADY,
	sum_59_s_axi_control_ARVALID,
	sum_59_s_axi_control_ARADDR,
	sum_59_s_axi_control_RREADY,
	sum_59_s_axi_control_RVALID,
	sum_59_s_axi_control_RDATA,
	sum_59_s_axi_control_RRESP,
	sum_59_s_axi_control_AWREADY,
	sum_59_s_axi_control_AWVALID,
	sum_59_s_axi_control_AWADDR,
	sum_59_s_axi_control_WREADY,
	sum_59_s_axi_control_WVALID,
	sum_59_s_axi_control_WDATA,
	sum_59_s_axi_control_WSTRB,
	sum_59_s_axi_control_BREADY,
	sum_59_s_axi_control_BVALID,
	sum_59_s_axi_control_BRESP,
	sum_60_m_axi_gmem_ARREADY,
	sum_60_m_axi_gmem_ARVALID,
	sum_60_m_axi_gmem_ARID,
	sum_60_m_axi_gmem_ARADDR,
	sum_60_m_axi_gmem_ARLEN,
	sum_60_m_axi_gmem_ARSIZE,
	sum_60_m_axi_gmem_ARBURST,
	sum_60_m_axi_gmem_ARLOCK,
	sum_60_m_axi_gmem_ARCACHE,
	sum_60_m_axi_gmem_ARPROT,
	sum_60_m_axi_gmem_ARQOS,
	sum_60_m_axi_gmem_ARREGION,
	sum_60_m_axi_gmem_ARUSER,
	sum_60_m_axi_gmem_RREADY,
	sum_60_m_axi_gmem_RVALID,
	sum_60_m_axi_gmem_RID,
	sum_60_m_axi_gmem_RDATA,
	sum_60_m_axi_gmem_RRESP,
	sum_60_m_axi_gmem_RLAST,
	sum_60_m_axi_gmem_RUSER,
	sum_60_m_axi_gmem_AWREADY,
	sum_60_m_axi_gmem_AWVALID,
	sum_60_m_axi_gmem_AWID,
	sum_60_m_axi_gmem_AWADDR,
	sum_60_m_axi_gmem_AWLEN,
	sum_60_m_axi_gmem_AWSIZE,
	sum_60_m_axi_gmem_AWBURST,
	sum_60_m_axi_gmem_AWLOCK,
	sum_60_m_axi_gmem_AWCACHE,
	sum_60_m_axi_gmem_AWPROT,
	sum_60_m_axi_gmem_AWQOS,
	sum_60_m_axi_gmem_AWREGION,
	sum_60_m_axi_gmem_AWUSER,
	sum_60_m_axi_gmem_WREADY,
	sum_60_m_axi_gmem_WVALID,
	sum_60_m_axi_gmem_WDATA,
	sum_60_m_axi_gmem_WSTRB,
	sum_60_m_axi_gmem_WLAST,
	sum_60_m_axi_gmem_WUSER,
	sum_60_m_axi_gmem_BREADY,
	sum_60_m_axi_gmem_BVALID,
	sum_60_m_axi_gmem_BID,
	sum_60_m_axi_gmem_BRESP,
	sum_60_m_axi_gmem_BUSER,
	sum_60_s_axi_control_ARREADY,
	sum_60_s_axi_control_ARVALID,
	sum_60_s_axi_control_ARADDR,
	sum_60_s_axi_control_RREADY,
	sum_60_s_axi_control_RVALID,
	sum_60_s_axi_control_RDATA,
	sum_60_s_axi_control_RRESP,
	sum_60_s_axi_control_AWREADY,
	sum_60_s_axi_control_AWVALID,
	sum_60_s_axi_control_AWADDR,
	sum_60_s_axi_control_WREADY,
	sum_60_s_axi_control_WVALID,
	sum_60_s_axi_control_WDATA,
	sum_60_s_axi_control_WSTRB,
	sum_60_s_axi_control_BREADY,
	sum_60_s_axi_control_BVALID,
	sum_60_s_axi_control_BRESP,
	sum_61_m_axi_gmem_ARREADY,
	sum_61_m_axi_gmem_ARVALID,
	sum_61_m_axi_gmem_ARID,
	sum_61_m_axi_gmem_ARADDR,
	sum_61_m_axi_gmem_ARLEN,
	sum_61_m_axi_gmem_ARSIZE,
	sum_61_m_axi_gmem_ARBURST,
	sum_61_m_axi_gmem_ARLOCK,
	sum_61_m_axi_gmem_ARCACHE,
	sum_61_m_axi_gmem_ARPROT,
	sum_61_m_axi_gmem_ARQOS,
	sum_61_m_axi_gmem_ARREGION,
	sum_61_m_axi_gmem_ARUSER,
	sum_61_m_axi_gmem_RREADY,
	sum_61_m_axi_gmem_RVALID,
	sum_61_m_axi_gmem_RID,
	sum_61_m_axi_gmem_RDATA,
	sum_61_m_axi_gmem_RRESP,
	sum_61_m_axi_gmem_RLAST,
	sum_61_m_axi_gmem_RUSER,
	sum_61_m_axi_gmem_AWREADY,
	sum_61_m_axi_gmem_AWVALID,
	sum_61_m_axi_gmem_AWID,
	sum_61_m_axi_gmem_AWADDR,
	sum_61_m_axi_gmem_AWLEN,
	sum_61_m_axi_gmem_AWSIZE,
	sum_61_m_axi_gmem_AWBURST,
	sum_61_m_axi_gmem_AWLOCK,
	sum_61_m_axi_gmem_AWCACHE,
	sum_61_m_axi_gmem_AWPROT,
	sum_61_m_axi_gmem_AWQOS,
	sum_61_m_axi_gmem_AWREGION,
	sum_61_m_axi_gmem_AWUSER,
	sum_61_m_axi_gmem_WREADY,
	sum_61_m_axi_gmem_WVALID,
	sum_61_m_axi_gmem_WDATA,
	sum_61_m_axi_gmem_WSTRB,
	sum_61_m_axi_gmem_WLAST,
	sum_61_m_axi_gmem_WUSER,
	sum_61_m_axi_gmem_BREADY,
	sum_61_m_axi_gmem_BVALID,
	sum_61_m_axi_gmem_BID,
	sum_61_m_axi_gmem_BRESP,
	sum_61_m_axi_gmem_BUSER,
	sum_61_s_axi_control_ARREADY,
	sum_61_s_axi_control_ARVALID,
	sum_61_s_axi_control_ARADDR,
	sum_61_s_axi_control_RREADY,
	sum_61_s_axi_control_RVALID,
	sum_61_s_axi_control_RDATA,
	sum_61_s_axi_control_RRESP,
	sum_61_s_axi_control_AWREADY,
	sum_61_s_axi_control_AWVALID,
	sum_61_s_axi_control_AWADDR,
	sum_61_s_axi_control_WREADY,
	sum_61_s_axi_control_WVALID,
	sum_61_s_axi_control_WDATA,
	sum_61_s_axi_control_WSTRB,
	sum_61_s_axi_control_BREADY,
	sum_61_s_axi_control_BVALID,
	sum_61_s_axi_control_BRESP,
	sum_62_m_axi_gmem_ARREADY,
	sum_62_m_axi_gmem_ARVALID,
	sum_62_m_axi_gmem_ARID,
	sum_62_m_axi_gmem_ARADDR,
	sum_62_m_axi_gmem_ARLEN,
	sum_62_m_axi_gmem_ARSIZE,
	sum_62_m_axi_gmem_ARBURST,
	sum_62_m_axi_gmem_ARLOCK,
	sum_62_m_axi_gmem_ARCACHE,
	sum_62_m_axi_gmem_ARPROT,
	sum_62_m_axi_gmem_ARQOS,
	sum_62_m_axi_gmem_ARREGION,
	sum_62_m_axi_gmem_ARUSER,
	sum_62_m_axi_gmem_RREADY,
	sum_62_m_axi_gmem_RVALID,
	sum_62_m_axi_gmem_RID,
	sum_62_m_axi_gmem_RDATA,
	sum_62_m_axi_gmem_RRESP,
	sum_62_m_axi_gmem_RLAST,
	sum_62_m_axi_gmem_RUSER,
	sum_62_m_axi_gmem_AWREADY,
	sum_62_m_axi_gmem_AWVALID,
	sum_62_m_axi_gmem_AWID,
	sum_62_m_axi_gmem_AWADDR,
	sum_62_m_axi_gmem_AWLEN,
	sum_62_m_axi_gmem_AWSIZE,
	sum_62_m_axi_gmem_AWBURST,
	sum_62_m_axi_gmem_AWLOCK,
	sum_62_m_axi_gmem_AWCACHE,
	sum_62_m_axi_gmem_AWPROT,
	sum_62_m_axi_gmem_AWQOS,
	sum_62_m_axi_gmem_AWREGION,
	sum_62_m_axi_gmem_AWUSER,
	sum_62_m_axi_gmem_WREADY,
	sum_62_m_axi_gmem_WVALID,
	sum_62_m_axi_gmem_WDATA,
	sum_62_m_axi_gmem_WSTRB,
	sum_62_m_axi_gmem_WLAST,
	sum_62_m_axi_gmem_WUSER,
	sum_62_m_axi_gmem_BREADY,
	sum_62_m_axi_gmem_BVALID,
	sum_62_m_axi_gmem_BID,
	sum_62_m_axi_gmem_BRESP,
	sum_62_m_axi_gmem_BUSER,
	sum_62_s_axi_control_ARREADY,
	sum_62_s_axi_control_ARVALID,
	sum_62_s_axi_control_ARADDR,
	sum_62_s_axi_control_RREADY,
	sum_62_s_axi_control_RVALID,
	sum_62_s_axi_control_RDATA,
	sum_62_s_axi_control_RRESP,
	sum_62_s_axi_control_AWREADY,
	sum_62_s_axi_control_AWVALID,
	sum_62_s_axi_control_AWADDR,
	sum_62_s_axi_control_WREADY,
	sum_62_s_axi_control_WVALID,
	sum_62_s_axi_control_WDATA,
	sum_62_s_axi_control_WSTRB,
	sum_62_s_axi_control_BREADY,
	sum_62_s_axi_control_BVALID,
	sum_62_s_axi_control_BRESP,
	sum_63_m_axi_gmem_ARREADY,
	sum_63_m_axi_gmem_ARVALID,
	sum_63_m_axi_gmem_ARID,
	sum_63_m_axi_gmem_ARADDR,
	sum_63_m_axi_gmem_ARLEN,
	sum_63_m_axi_gmem_ARSIZE,
	sum_63_m_axi_gmem_ARBURST,
	sum_63_m_axi_gmem_ARLOCK,
	sum_63_m_axi_gmem_ARCACHE,
	sum_63_m_axi_gmem_ARPROT,
	sum_63_m_axi_gmem_ARQOS,
	sum_63_m_axi_gmem_ARREGION,
	sum_63_m_axi_gmem_ARUSER,
	sum_63_m_axi_gmem_RREADY,
	sum_63_m_axi_gmem_RVALID,
	sum_63_m_axi_gmem_RID,
	sum_63_m_axi_gmem_RDATA,
	sum_63_m_axi_gmem_RRESP,
	sum_63_m_axi_gmem_RLAST,
	sum_63_m_axi_gmem_RUSER,
	sum_63_m_axi_gmem_AWREADY,
	sum_63_m_axi_gmem_AWVALID,
	sum_63_m_axi_gmem_AWID,
	sum_63_m_axi_gmem_AWADDR,
	sum_63_m_axi_gmem_AWLEN,
	sum_63_m_axi_gmem_AWSIZE,
	sum_63_m_axi_gmem_AWBURST,
	sum_63_m_axi_gmem_AWLOCK,
	sum_63_m_axi_gmem_AWCACHE,
	sum_63_m_axi_gmem_AWPROT,
	sum_63_m_axi_gmem_AWQOS,
	sum_63_m_axi_gmem_AWREGION,
	sum_63_m_axi_gmem_AWUSER,
	sum_63_m_axi_gmem_WREADY,
	sum_63_m_axi_gmem_WVALID,
	sum_63_m_axi_gmem_WDATA,
	sum_63_m_axi_gmem_WSTRB,
	sum_63_m_axi_gmem_WLAST,
	sum_63_m_axi_gmem_WUSER,
	sum_63_m_axi_gmem_BREADY,
	sum_63_m_axi_gmem_BVALID,
	sum_63_m_axi_gmem_BID,
	sum_63_m_axi_gmem_BRESP,
	sum_63_m_axi_gmem_BUSER,
	sum_63_s_axi_control_ARREADY,
	sum_63_s_axi_control_ARVALID,
	sum_63_s_axi_control_ARADDR,
	sum_63_s_axi_control_RREADY,
	sum_63_s_axi_control_RVALID,
	sum_63_s_axi_control_RDATA,
	sum_63_s_axi_control_RRESP,
	sum_63_s_axi_control_AWREADY,
	sum_63_s_axi_control_AWVALID,
	sum_63_s_axi_control_AWADDR,
	sum_63_s_axi_control_WREADY,
	sum_63_s_axi_control_WVALID,
	sum_63_s_axi_control_WDATA,
	sum_63_s_axi_control_WSTRB,
	sum_63_s_axi_control_BREADY,
	sum_63_s_axi_control_BVALID,
	sum_63_s_axi_control_BRESP,
	sum_schedulerAXI_0_ARREADY,
	sum_schedulerAXI_0_ARVALID,
	sum_schedulerAXI_0_ARID,
	sum_schedulerAXI_0_ARADDR,
	sum_schedulerAXI_0_ARLEN,
	sum_schedulerAXI_0_ARSIZE,
	sum_schedulerAXI_0_ARBURST,
	sum_schedulerAXI_0_ARLOCK,
	sum_schedulerAXI_0_ARCACHE,
	sum_schedulerAXI_0_ARPROT,
	sum_schedulerAXI_0_ARQOS,
	sum_schedulerAXI_0_ARREGION,
	sum_schedulerAXI_0_RREADY,
	sum_schedulerAXI_0_RVALID,
	sum_schedulerAXI_0_RID,
	sum_schedulerAXI_0_RDATA,
	sum_schedulerAXI_0_RRESP,
	sum_schedulerAXI_0_RLAST,
	sum_schedulerAXI_0_AWREADY,
	sum_schedulerAXI_0_AWVALID,
	sum_schedulerAXI_0_AWID,
	sum_schedulerAXI_0_AWADDR,
	sum_schedulerAXI_0_AWLEN,
	sum_schedulerAXI_0_AWSIZE,
	sum_schedulerAXI_0_AWBURST,
	sum_schedulerAXI_0_AWLOCK,
	sum_schedulerAXI_0_AWCACHE,
	sum_schedulerAXI_0_AWPROT,
	sum_schedulerAXI_0_AWQOS,
	sum_schedulerAXI_0_AWREGION,
	sum_schedulerAXI_0_WREADY,
	sum_schedulerAXI_0_WVALID,
	sum_schedulerAXI_0_WDATA,
	sum_schedulerAXI_0_WSTRB,
	sum_schedulerAXI_0_WLAST,
	sum_schedulerAXI_0_BREADY,
	sum_schedulerAXI_0_BVALID,
	sum_schedulerAXI_0_BID,
	sum_schedulerAXI_0_BRESP,
	sum_closureAllocatorAXI_0_ARREADY,
	sum_closureAllocatorAXI_0_ARVALID,
	sum_closureAllocatorAXI_0_ARID,
	sum_closureAllocatorAXI_0_ARADDR,
	sum_closureAllocatorAXI_0_ARLEN,
	sum_closureAllocatorAXI_0_ARSIZE,
	sum_closureAllocatorAXI_0_ARBURST,
	sum_closureAllocatorAXI_0_ARLOCK,
	sum_closureAllocatorAXI_0_ARCACHE,
	sum_closureAllocatorAXI_0_ARPROT,
	sum_closureAllocatorAXI_0_ARQOS,
	sum_closureAllocatorAXI_0_ARREGION,
	sum_closureAllocatorAXI_0_RREADY,
	sum_closureAllocatorAXI_0_RVALID,
	sum_closureAllocatorAXI_0_RID,
	sum_closureAllocatorAXI_0_RDATA,
	sum_closureAllocatorAXI_0_RRESP,
	sum_closureAllocatorAXI_0_RLAST,
	sum_closureAllocatorAXI_0_AWREADY,
	sum_closureAllocatorAXI_0_AWVALID,
	sum_closureAllocatorAXI_0_AWID,
	sum_closureAllocatorAXI_0_AWADDR,
	sum_closureAllocatorAXI_0_AWLEN,
	sum_closureAllocatorAXI_0_AWSIZE,
	sum_closureAllocatorAXI_0_AWBURST,
	sum_closureAllocatorAXI_0_AWLOCK,
	sum_closureAllocatorAXI_0_AWCACHE,
	sum_closureAllocatorAXI_0_AWPROT,
	sum_closureAllocatorAXI_0_AWQOS,
	sum_closureAllocatorAXI_0_AWREGION,
	sum_closureAllocatorAXI_0_WREADY,
	sum_closureAllocatorAXI_0_WVALID,
	sum_closureAllocatorAXI_0_WDATA,
	sum_closureAllocatorAXI_0_WSTRB,
	sum_closureAllocatorAXI_0_WLAST,
	sum_closureAllocatorAXI_0_BREADY,
	sum_closureAllocatorAXI_0_BVALID,
	sum_closureAllocatorAXI_0_BID,
	sum_closureAllocatorAXI_0_BRESP,
	sum_argumentNotifierAXI_0_ARREADY,
	sum_argumentNotifierAXI_0_ARVALID,
	sum_argumentNotifierAXI_0_ARID,
	sum_argumentNotifierAXI_0_ARADDR,
	sum_argumentNotifierAXI_0_ARLEN,
	sum_argumentNotifierAXI_0_ARSIZE,
	sum_argumentNotifierAXI_0_ARBURST,
	sum_argumentNotifierAXI_0_ARLOCK,
	sum_argumentNotifierAXI_0_ARCACHE,
	sum_argumentNotifierAXI_0_ARPROT,
	sum_argumentNotifierAXI_0_ARQOS,
	sum_argumentNotifierAXI_0_ARREGION,
	sum_argumentNotifierAXI_0_RREADY,
	sum_argumentNotifierAXI_0_RVALID,
	sum_argumentNotifierAXI_0_RID,
	sum_argumentNotifierAXI_0_RDATA,
	sum_argumentNotifierAXI_0_RRESP,
	sum_argumentNotifierAXI_0_RLAST,
	sum_argumentNotifierAXI_0_AWREADY,
	sum_argumentNotifierAXI_0_AWVALID,
	sum_argumentNotifierAXI_0_AWID,
	sum_argumentNotifierAXI_0_AWADDR,
	sum_argumentNotifierAXI_0_AWLEN,
	sum_argumentNotifierAXI_0_AWSIZE,
	sum_argumentNotifierAXI_0_AWBURST,
	sum_argumentNotifierAXI_0_AWLOCK,
	sum_argumentNotifierAXI_0_AWCACHE,
	sum_argumentNotifierAXI_0_AWPROT,
	sum_argumentNotifierAXI_0_AWQOS,
	sum_argumentNotifierAXI_0_AWREGION,
	sum_argumentNotifierAXI_0_WREADY,
	sum_argumentNotifierAXI_0_WVALID,
	sum_argumentNotifierAXI_0_WDATA,
	sum_argumentNotifierAXI_0_WSTRB,
	sum_argumentNotifierAXI_0_WLAST,
	sum_argumentNotifierAXI_0_BREADY,
	sum_argumentNotifierAXI_0_BVALID,
	sum_argumentNotifierAXI_0_BID,
	sum_argumentNotifierAXI_0_BRESP
);
	input clock;
	input reset;
	output wire s_axil_mgmt_hardcilk_ARREADY;
	input s_axil_mgmt_hardcilk_ARVALID;
	input [13:0] s_axil_mgmt_hardcilk_ARADDR;
	input [2:0] s_axil_mgmt_hardcilk_ARPROT;
	input s_axil_mgmt_hardcilk_RREADY;
	output wire s_axil_mgmt_hardcilk_RVALID;
	output wire [63:0] s_axil_mgmt_hardcilk_RDATA;
	output wire [1:0] s_axil_mgmt_hardcilk_RRESP;
	output wire s_axil_mgmt_hardcilk_AWREADY;
	input s_axil_mgmt_hardcilk_AWVALID;
	input [13:0] s_axil_mgmt_hardcilk_AWADDR;
	input [2:0] s_axil_mgmt_hardcilk_AWPROT;
	output wire s_axil_mgmt_hardcilk_WREADY;
	input s_axil_mgmt_hardcilk_WVALID;
	input [63:0] s_axil_mgmt_hardcilk_WDATA;
	input [7:0] s_axil_mgmt_hardcilk_WSTRB;
	input s_axil_mgmt_hardcilk_BREADY;
	output wire s_axil_mgmt_hardcilk_BVALID;
	output wire [1:0] s_axil_mgmt_hardcilk_BRESP;
	input fib_0_m_axi_gmem_ARREADY;
	output wire fib_0_m_axi_gmem_ARVALID;
	output wire fib_0_m_axi_gmem_ARID;
	output wire [63:0] fib_0_m_axi_gmem_ARADDR;
	output wire [7:0] fib_0_m_axi_gmem_ARLEN;
	output wire [2:0] fib_0_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_0_m_axi_gmem_ARBURST;
	output wire fib_0_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_0_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_0_m_axi_gmem_ARPROT;
	output wire [3:0] fib_0_m_axi_gmem_ARQOS;
	output wire [3:0] fib_0_m_axi_gmem_ARREGION;
	output wire fib_0_m_axi_gmem_ARUSER;
	output wire fib_0_m_axi_gmem_RREADY;
	input fib_0_m_axi_gmem_RVALID;
	input fib_0_m_axi_gmem_RID;
	input [63:0] fib_0_m_axi_gmem_RDATA;
	input [1:0] fib_0_m_axi_gmem_RRESP;
	input fib_0_m_axi_gmem_RLAST;
	input fib_0_m_axi_gmem_RUSER;
	input fib_0_m_axi_gmem_AWREADY;
	output wire fib_0_m_axi_gmem_AWVALID;
	output wire fib_0_m_axi_gmem_AWID;
	output wire [63:0] fib_0_m_axi_gmem_AWADDR;
	output wire [7:0] fib_0_m_axi_gmem_AWLEN;
	output wire [2:0] fib_0_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_0_m_axi_gmem_AWBURST;
	output wire fib_0_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_0_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_0_m_axi_gmem_AWPROT;
	output wire [3:0] fib_0_m_axi_gmem_AWQOS;
	output wire [3:0] fib_0_m_axi_gmem_AWREGION;
	output wire fib_0_m_axi_gmem_AWUSER;
	input fib_0_m_axi_gmem_WREADY;
	output wire fib_0_m_axi_gmem_WVALID;
	output wire [63:0] fib_0_m_axi_gmem_WDATA;
	output wire [7:0] fib_0_m_axi_gmem_WSTRB;
	output wire fib_0_m_axi_gmem_WLAST;
	output wire fib_0_m_axi_gmem_WUSER;
	output wire fib_0_m_axi_gmem_BREADY;
	input fib_0_m_axi_gmem_BVALID;
	input fib_0_m_axi_gmem_BID;
	input [1:0] fib_0_m_axi_gmem_BRESP;
	input fib_0_m_axi_gmem_BUSER;
	output wire fib_0_s_axi_control_ARREADY;
	input fib_0_s_axi_control_ARVALID;
	input [4:0] fib_0_s_axi_control_ARADDR;
	input fib_0_s_axi_control_RREADY;
	output wire fib_0_s_axi_control_RVALID;
	output wire [31:0] fib_0_s_axi_control_RDATA;
	output wire [1:0] fib_0_s_axi_control_RRESP;
	output wire fib_0_s_axi_control_AWREADY;
	input fib_0_s_axi_control_AWVALID;
	input [4:0] fib_0_s_axi_control_AWADDR;
	output wire fib_0_s_axi_control_WREADY;
	input fib_0_s_axi_control_WVALID;
	input [31:0] fib_0_s_axi_control_WDATA;
	input [3:0] fib_0_s_axi_control_WSTRB;
	input fib_0_s_axi_control_BREADY;
	output wire fib_0_s_axi_control_BVALID;
	output wire [1:0] fib_0_s_axi_control_BRESP;
	input fib_1_m_axi_gmem_ARREADY;
	output wire fib_1_m_axi_gmem_ARVALID;
	output wire fib_1_m_axi_gmem_ARID;
	output wire [63:0] fib_1_m_axi_gmem_ARADDR;
	output wire [7:0] fib_1_m_axi_gmem_ARLEN;
	output wire [2:0] fib_1_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_1_m_axi_gmem_ARBURST;
	output wire fib_1_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_1_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_1_m_axi_gmem_ARPROT;
	output wire [3:0] fib_1_m_axi_gmem_ARQOS;
	output wire [3:0] fib_1_m_axi_gmem_ARREGION;
	output wire fib_1_m_axi_gmem_ARUSER;
	output wire fib_1_m_axi_gmem_RREADY;
	input fib_1_m_axi_gmem_RVALID;
	input fib_1_m_axi_gmem_RID;
	input [63:0] fib_1_m_axi_gmem_RDATA;
	input [1:0] fib_1_m_axi_gmem_RRESP;
	input fib_1_m_axi_gmem_RLAST;
	input fib_1_m_axi_gmem_RUSER;
	input fib_1_m_axi_gmem_AWREADY;
	output wire fib_1_m_axi_gmem_AWVALID;
	output wire fib_1_m_axi_gmem_AWID;
	output wire [63:0] fib_1_m_axi_gmem_AWADDR;
	output wire [7:0] fib_1_m_axi_gmem_AWLEN;
	output wire [2:0] fib_1_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_1_m_axi_gmem_AWBURST;
	output wire fib_1_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_1_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_1_m_axi_gmem_AWPROT;
	output wire [3:0] fib_1_m_axi_gmem_AWQOS;
	output wire [3:0] fib_1_m_axi_gmem_AWREGION;
	output wire fib_1_m_axi_gmem_AWUSER;
	input fib_1_m_axi_gmem_WREADY;
	output wire fib_1_m_axi_gmem_WVALID;
	output wire [63:0] fib_1_m_axi_gmem_WDATA;
	output wire [7:0] fib_1_m_axi_gmem_WSTRB;
	output wire fib_1_m_axi_gmem_WLAST;
	output wire fib_1_m_axi_gmem_WUSER;
	output wire fib_1_m_axi_gmem_BREADY;
	input fib_1_m_axi_gmem_BVALID;
	input fib_1_m_axi_gmem_BID;
	input [1:0] fib_1_m_axi_gmem_BRESP;
	input fib_1_m_axi_gmem_BUSER;
	output wire fib_1_s_axi_control_ARREADY;
	input fib_1_s_axi_control_ARVALID;
	input [4:0] fib_1_s_axi_control_ARADDR;
	input fib_1_s_axi_control_RREADY;
	output wire fib_1_s_axi_control_RVALID;
	output wire [31:0] fib_1_s_axi_control_RDATA;
	output wire [1:0] fib_1_s_axi_control_RRESP;
	output wire fib_1_s_axi_control_AWREADY;
	input fib_1_s_axi_control_AWVALID;
	input [4:0] fib_1_s_axi_control_AWADDR;
	output wire fib_1_s_axi_control_WREADY;
	input fib_1_s_axi_control_WVALID;
	input [31:0] fib_1_s_axi_control_WDATA;
	input [3:0] fib_1_s_axi_control_WSTRB;
	input fib_1_s_axi_control_BREADY;
	output wire fib_1_s_axi_control_BVALID;
	output wire [1:0] fib_1_s_axi_control_BRESP;
	input fib_2_m_axi_gmem_ARREADY;
	output wire fib_2_m_axi_gmem_ARVALID;
	output wire fib_2_m_axi_gmem_ARID;
	output wire [63:0] fib_2_m_axi_gmem_ARADDR;
	output wire [7:0] fib_2_m_axi_gmem_ARLEN;
	output wire [2:0] fib_2_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_2_m_axi_gmem_ARBURST;
	output wire fib_2_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_2_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_2_m_axi_gmem_ARPROT;
	output wire [3:0] fib_2_m_axi_gmem_ARQOS;
	output wire [3:0] fib_2_m_axi_gmem_ARREGION;
	output wire fib_2_m_axi_gmem_ARUSER;
	output wire fib_2_m_axi_gmem_RREADY;
	input fib_2_m_axi_gmem_RVALID;
	input fib_2_m_axi_gmem_RID;
	input [63:0] fib_2_m_axi_gmem_RDATA;
	input [1:0] fib_2_m_axi_gmem_RRESP;
	input fib_2_m_axi_gmem_RLAST;
	input fib_2_m_axi_gmem_RUSER;
	input fib_2_m_axi_gmem_AWREADY;
	output wire fib_2_m_axi_gmem_AWVALID;
	output wire fib_2_m_axi_gmem_AWID;
	output wire [63:0] fib_2_m_axi_gmem_AWADDR;
	output wire [7:0] fib_2_m_axi_gmem_AWLEN;
	output wire [2:0] fib_2_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_2_m_axi_gmem_AWBURST;
	output wire fib_2_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_2_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_2_m_axi_gmem_AWPROT;
	output wire [3:0] fib_2_m_axi_gmem_AWQOS;
	output wire [3:0] fib_2_m_axi_gmem_AWREGION;
	output wire fib_2_m_axi_gmem_AWUSER;
	input fib_2_m_axi_gmem_WREADY;
	output wire fib_2_m_axi_gmem_WVALID;
	output wire [63:0] fib_2_m_axi_gmem_WDATA;
	output wire [7:0] fib_2_m_axi_gmem_WSTRB;
	output wire fib_2_m_axi_gmem_WLAST;
	output wire fib_2_m_axi_gmem_WUSER;
	output wire fib_2_m_axi_gmem_BREADY;
	input fib_2_m_axi_gmem_BVALID;
	input fib_2_m_axi_gmem_BID;
	input [1:0] fib_2_m_axi_gmem_BRESP;
	input fib_2_m_axi_gmem_BUSER;
	output wire fib_2_s_axi_control_ARREADY;
	input fib_2_s_axi_control_ARVALID;
	input [4:0] fib_2_s_axi_control_ARADDR;
	input fib_2_s_axi_control_RREADY;
	output wire fib_2_s_axi_control_RVALID;
	output wire [31:0] fib_2_s_axi_control_RDATA;
	output wire [1:0] fib_2_s_axi_control_RRESP;
	output wire fib_2_s_axi_control_AWREADY;
	input fib_2_s_axi_control_AWVALID;
	input [4:0] fib_2_s_axi_control_AWADDR;
	output wire fib_2_s_axi_control_WREADY;
	input fib_2_s_axi_control_WVALID;
	input [31:0] fib_2_s_axi_control_WDATA;
	input [3:0] fib_2_s_axi_control_WSTRB;
	input fib_2_s_axi_control_BREADY;
	output wire fib_2_s_axi_control_BVALID;
	output wire [1:0] fib_2_s_axi_control_BRESP;
	input fib_3_m_axi_gmem_ARREADY;
	output wire fib_3_m_axi_gmem_ARVALID;
	output wire fib_3_m_axi_gmem_ARID;
	output wire [63:0] fib_3_m_axi_gmem_ARADDR;
	output wire [7:0] fib_3_m_axi_gmem_ARLEN;
	output wire [2:0] fib_3_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_3_m_axi_gmem_ARBURST;
	output wire fib_3_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_3_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_3_m_axi_gmem_ARPROT;
	output wire [3:0] fib_3_m_axi_gmem_ARQOS;
	output wire [3:0] fib_3_m_axi_gmem_ARREGION;
	output wire fib_3_m_axi_gmem_ARUSER;
	output wire fib_3_m_axi_gmem_RREADY;
	input fib_3_m_axi_gmem_RVALID;
	input fib_3_m_axi_gmem_RID;
	input [63:0] fib_3_m_axi_gmem_RDATA;
	input [1:0] fib_3_m_axi_gmem_RRESP;
	input fib_3_m_axi_gmem_RLAST;
	input fib_3_m_axi_gmem_RUSER;
	input fib_3_m_axi_gmem_AWREADY;
	output wire fib_3_m_axi_gmem_AWVALID;
	output wire fib_3_m_axi_gmem_AWID;
	output wire [63:0] fib_3_m_axi_gmem_AWADDR;
	output wire [7:0] fib_3_m_axi_gmem_AWLEN;
	output wire [2:0] fib_3_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_3_m_axi_gmem_AWBURST;
	output wire fib_3_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_3_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_3_m_axi_gmem_AWPROT;
	output wire [3:0] fib_3_m_axi_gmem_AWQOS;
	output wire [3:0] fib_3_m_axi_gmem_AWREGION;
	output wire fib_3_m_axi_gmem_AWUSER;
	input fib_3_m_axi_gmem_WREADY;
	output wire fib_3_m_axi_gmem_WVALID;
	output wire [63:0] fib_3_m_axi_gmem_WDATA;
	output wire [7:0] fib_3_m_axi_gmem_WSTRB;
	output wire fib_3_m_axi_gmem_WLAST;
	output wire fib_3_m_axi_gmem_WUSER;
	output wire fib_3_m_axi_gmem_BREADY;
	input fib_3_m_axi_gmem_BVALID;
	input fib_3_m_axi_gmem_BID;
	input [1:0] fib_3_m_axi_gmem_BRESP;
	input fib_3_m_axi_gmem_BUSER;
	output wire fib_3_s_axi_control_ARREADY;
	input fib_3_s_axi_control_ARVALID;
	input [4:0] fib_3_s_axi_control_ARADDR;
	input fib_3_s_axi_control_RREADY;
	output wire fib_3_s_axi_control_RVALID;
	output wire [31:0] fib_3_s_axi_control_RDATA;
	output wire [1:0] fib_3_s_axi_control_RRESP;
	output wire fib_3_s_axi_control_AWREADY;
	input fib_3_s_axi_control_AWVALID;
	input [4:0] fib_3_s_axi_control_AWADDR;
	output wire fib_3_s_axi_control_WREADY;
	input fib_3_s_axi_control_WVALID;
	input [31:0] fib_3_s_axi_control_WDATA;
	input [3:0] fib_3_s_axi_control_WSTRB;
	input fib_3_s_axi_control_BREADY;
	output wire fib_3_s_axi_control_BVALID;
	output wire [1:0] fib_3_s_axi_control_BRESP;
	input fib_4_m_axi_gmem_ARREADY;
	output wire fib_4_m_axi_gmem_ARVALID;
	output wire fib_4_m_axi_gmem_ARID;
	output wire [63:0] fib_4_m_axi_gmem_ARADDR;
	output wire [7:0] fib_4_m_axi_gmem_ARLEN;
	output wire [2:0] fib_4_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_4_m_axi_gmem_ARBURST;
	output wire fib_4_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_4_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_4_m_axi_gmem_ARPROT;
	output wire [3:0] fib_4_m_axi_gmem_ARQOS;
	output wire [3:0] fib_4_m_axi_gmem_ARREGION;
	output wire fib_4_m_axi_gmem_ARUSER;
	output wire fib_4_m_axi_gmem_RREADY;
	input fib_4_m_axi_gmem_RVALID;
	input fib_4_m_axi_gmem_RID;
	input [63:0] fib_4_m_axi_gmem_RDATA;
	input [1:0] fib_4_m_axi_gmem_RRESP;
	input fib_4_m_axi_gmem_RLAST;
	input fib_4_m_axi_gmem_RUSER;
	input fib_4_m_axi_gmem_AWREADY;
	output wire fib_4_m_axi_gmem_AWVALID;
	output wire fib_4_m_axi_gmem_AWID;
	output wire [63:0] fib_4_m_axi_gmem_AWADDR;
	output wire [7:0] fib_4_m_axi_gmem_AWLEN;
	output wire [2:0] fib_4_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_4_m_axi_gmem_AWBURST;
	output wire fib_4_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_4_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_4_m_axi_gmem_AWPROT;
	output wire [3:0] fib_4_m_axi_gmem_AWQOS;
	output wire [3:0] fib_4_m_axi_gmem_AWREGION;
	output wire fib_4_m_axi_gmem_AWUSER;
	input fib_4_m_axi_gmem_WREADY;
	output wire fib_4_m_axi_gmem_WVALID;
	output wire [63:0] fib_4_m_axi_gmem_WDATA;
	output wire [7:0] fib_4_m_axi_gmem_WSTRB;
	output wire fib_4_m_axi_gmem_WLAST;
	output wire fib_4_m_axi_gmem_WUSER;
	output wire fib_4_m_axi_gmem_BREADY;
	input fib_4_m_axi_gmem_BVALID;
	input fib_4_m_axi_gmem_BID;
	input [1:0] fib_4_m_axi_gmem_BRESP;
	input fib_4_m_axi_gmem_BUSER;
	output wire fib_4_s_axi_control_ARREADY;
	input fib_4_s_axi_control_ARVALID;
	input [4:0] fib_4_s_axi_control_ARADDR;
	input fib_4_s_axi_control_RREADY;
	output wire fib_4_s_axi_control_RVALID;
	output wire [31:0] fib_4_s_axi_control_RDATA;
	output wire [1:0] fib_4_s_axi_control_RRESP;
	output wire fib_4_s_axi_control_AWREADY;
	input fib_4_s_axi_control_AWVALID;
	input [4:0] fib_4_s_axi_control_AWADDR;
	output wire fib_4_s_axi_control_WREADY;
	input fib_4_s_axi_control_WVALID;
	input [31:0] fib_4_s_axi_control_WDATA;
	input [3:0] fib_4_s_axi_control_WSTRB;
	input fib_4_s_axi_control_BREADY;
	output wire fib_4_s_axi_control_BVALID;
	output wire [1:0] fib_4_s_axi_control_BRESP;
	input fib_5_m_axi_gmem_ARREADY;
	output wire fib_5_m_axi_gmem_ARVALID;
	output wire fib_5_m_axi_gmem_ARID;
	output wire [63:0] fib_5_m_axi_gmem_ARADDR;
	output wire [7:0] fib_5_m_axi_gmem_ARLEN;
	output wire [2:0] fib_5_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_5_m_axi_gmem_ARBURST;
	output wire fib_5_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_5_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_5_m_axi_gmem_ARPROT;
	output wire [3:0] fib_5_m_axi_gmem_ARQOS;
	output wire [3:0] fib_5_m_axi_gmem_ARREGION;
	output wire fib_5_m_axi_gmem_ARUSER;
	output wire fib_5_m_axi_gmem_RREADY;
	input fib_5_m_axi_gmem_RVALID;
	input fib_5_m_axi_gmem_RID;
	input [63:0] fib_5_m_axi_gmem_RDATA;
	input [1:0] fib_5_m_axi_gmem_RRESP;
	input fib_5_m_axi_gmem_RLAST;
	input fib_5_m_axi_gmem_RUSER;
	input fib_5_m_axi_gmem_AWREADY;
	output wire fib_5_m_axi_gmem_AWVALID;
	output wire fib_5_m_axi_gmem_AWID;
	output wire [63:0] fib_5_m_axi_gmem_AWADDR;
	output wire [7:0] fib_5_m_axi_gmem_AWLEN;
	output wire [2:0] fib_5_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_5_m_axi_gmem_AWBURST;
	output wire fib_5_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_5_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_5_m_axi_gmem_AWPROT;
	output wire [3:0] fib_5_m_axi_gmem_AWQOS;
	output wire [3:0] fib_5_m_axi_gmem_AWREGION;
	output wire fib_5_m_axi_gmem_AWUSER;
	input fib_5_m_axi_gmem_WREADY;
	output wire fib_5_m_axi_gmem_WVALID;
	output wire [63:0] fib_5_m_axi_gmem_WDATA;
	output wire [7:0] fib_5_m_axi_gmem_WSTRB;
	output wire fib_5_m_axi_gmem_WLAST;
	output wire fib_5_m_axi_gmem_WUSER;
	output wire fib_5_m_axi_gmem_BREADY;
	input fib_5_m_axi_gmem_BVALID;
	input fib_5_m_axi_gmem_BID;
	input [1:0] fib_5_m_axi_gmem_BRESP;
	input fib_5_m_axi_gmem_BUSER;
	output wire fib_5_s_axi_control_ARREADY;
	input fib_5_s_axi_control_ARVALID;
	input [4:0] fib_5_s_axi_control_ARADDR;
	input fib_5_s_axi_control_RREADY;
	output wire fib_5_s_axi_control_RVALID;
	output wire [31:0] fib_5_s_axi_control_RDATA;
	output wire [1:0] fib_5_s_axi_control_RRESP;
	output wire fib_5_s_axi_control_AWREADY;
	input fib_5_s_axi_control_AWVALID;
	input [4:0] fib_5_s_axi_control_AWADDR;
	output wire fib_5_s_axi_control_WREADY;
	input fib_5_s_axi_control_WVALID;
	input [31:0] fib_5_s_axi_control_WDATA;
	input [3:0] fib_5_s_axi_control_WSTRB;
	input fib_5_s_axi_control_BREADY;
	output wire fib_5_s_axi_control_BVALID;
	output wire [1:0] fib_5_s_axi_control_BRESP;
	input fib_6_m_axi_gmem_ARREADY;
	output wire fib_6_m_axi_gmem_ARVALID;
	output wire fib_6_m_axi_gmem_ARID;
	output wire [63:0] fib_6_m_axi_gmem_ARADDR;
	output wire [7:0] fib_6_m_axi_gmem_ARLEN;
	output wire [2:0] fib_6_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_6_m_axi_gmem_ARBURST;
	output wire fib_6_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_6_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_6_m_axi_gmem_ARPROT;
	output wire [3:0] fib_6_m_axi_gmem_ARQOS;
	output wire [3:0] fib_6_m_axi_gmem_ARREGION;
	output wire fib_6_m_axi_gmem_ARUSER;
	output wire fib_6_m_axi_gmem_RREADY;
	input fib_6_m_axi_gmem_RVALID;
	input fib_6_m_axi_gmem_RID;
	input [63:0] fib_6_m_axi_gmem_RDATA;
	input [1:0] fib_6_m_axi_gmem_RRESP;
	input fib_6_m_axi_gmem_RLAST;
	input fib_6_m_axi_gmem_RUSER;
	input fib_6_m_axi_gmem_AWREADY;
	output wire fib_6_m_axi_gmem_AWVALID;
	output wire fib_6_m_axi_gmem_AWID;
	output wire [63:0] fib_6_m_axi_gmem_AWADDR;
	output wire [7:0] fib_6_m_axi_gmem_AWLEN;
	output wire [2:0] fib_6_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_6_m_axi_gmem_AWBURST;
	output wire fib_6_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_6_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_6_m_axi_gmem_AWPROT;
	output wire [3:0] fib_6_m_axi_gmem_AWQOS;
	output wire [3:0] fib_6_m_axi_gmem_AWREGION;
	output wire fib_6_m_axi_gmem_AWUSER;
	input fib_6_m_axi_gmem_WREADY;
	output wire fib_6_m_axi_gmem_WVALID;
	output wire [63:0] fib_6_m_axi_gmem_WDATA;
	output wire [7:0] fib_6_m_axi_gmem_WSTRB;
	output wire fib_6_m_axi_gmem_WLAST;
	output wire fib_6_m_axi_gmem_WUSER;
	output wire fib_6_m_axi_gmem_BREADY;
	input fib_6_m_axi_gmem_BVALID;
	input fib_6_m_axi_gmem_BID;
	input [1:0] fib_6_m_axi_gmem_BRESP;
	input fib_6_m_axi_gmem_BUSER;
	output wire fib_6_s_axi_control_ARREADY;
	input fib_6_s_axi_control_ARVALID;
	input [4:0] fib_6_s_axi_control_ARADDR;
	input fib_6_s_axi_control_RREADY;
	output wire fib_6_s_axi_control_RVALID;
	output wire [31:0] fib_6_s_axi_control_RDATA;
	output wire [1:0] fib_6_s_axi_control_RRESP;
	output wire fib_6_s_axi_control_AWREADY;
	input fib_6_s_axi_control_AWVALID;
	input [4:0] fib_6_s_axi_control_AWADDR;
	output wire fib_6_s_axi_control_WREADY;
	input fib_6_s_axi_control_WVALID;
	input [31:0] fib_6_s_axi_control_WDATA;
	input [3:0] fib_6_s_axi_control_WSTRB;
	input fib_6_s_axi_control_BREADY;
	output wire fib_6_s_axi_control_BVALID;
	output wire [1:0] fib_6_s_axi_control_BRESP;
	input fib_7_m_axi_gmem_ARREADY;
	output wire fib_7_m_axi_gmem_ARVALID;
	output wire fib_7_m_axi_gmem_ARID;
	output wire [63:0] fib_7_m_axi_gmem_ARADDR;
	output wire [7:0] fib_7_m_axi_gmem_ARLEN;
	output wire [2:0] fib_7_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_7_m_axi_gmem_ARBURST;
	output wire fib_7_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_7_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_7_m_axi_gmem_ARPROT;
	output wire [3:0] fib_7_m_axi_gmem_ARQOS;
	output wire [3:0] fib_7_m_axi_gmem_ARREGION;
	output wire fib_7_m_axi_gmem_ARUSER;
	output wire fib_7_m_axi_gmem_RREADY;
	input fib_7_m_axi_gmem_RVALID;
	input fib_7_m_axi_gmem_RID;
	input [63:0] fib_7_m_axi_gmem_RDATA;
	input [1:0] fib_7_m_axi_gmem_RRESP;
	input fib_7_m_axi_gmem_RLAST;
	input fib_7_m_axi_gmem_RUSER;
	input fib_7_m_axi_gmem_AWREADY;
	output wire fib_7_m_axi_gmem_AWVALID;
	output wire fib_7_m_axi_gmem_AWID;
	output wire [63:0] fib_7_m_axi_gmem_AWADDR;
	output wire [7:0] fib_7_m_axi_gmem_AWLEN;
	output wire [2:0] fib_7_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_7_m_axi_gmem_AWBURST;
	output wire fib_7_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_7_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_7_m_axi_gmem_AWPROT;
	output wire [3:0] fib_7_m_axi_gmem_AWQOS;
	output wire [3:0] fib_7_m_axi_gmem_AWREGION;
	output wire fib_7_m_axi_gmem_AWUSER;
	input fib_7_m_axi_gmem_WREADY;
	output wire fib_7_m_axi_gmem_WVALID;
	output wire [63:0] fib_7_m_axi_gmem_WDATA;
	output wire [7:0] fib_7_m_axi_gmem_WSTRB;
	output wire fib_7_m_axi_gmem_WLAST;
	output wire fib_7_m_axi_gmem_WUSER;
	output wire fib_7_m_axi_gmem_BREADY;
	input fib_7_m_axi_gmem_BVALID;
	input fib_7_m_axi_gmem_BID;
	input [1:0] fib_7_m_axi_gmem_BRESP;
	input fib_7_m_axi_gmem_BUSER;
	output wire fib_7_s_axi_control_ARREADY;
	input fib_7_s_axi_control_ARVALID;
	input [4:0] fib_7_s_axi_control_ARADDR;
	input fib_7_s_axi_control_RREADY;
	output wire fib_7_s_axi_control_RVALID;
	output wire [31:0] fib_7_s_axi_control_RDATA;
	output wire [1:0] fib_7_s_axi_control_RRESP;
	output wire fib_7_s_axi_control_AWREADY;
	input fib_7_s_axi_control_AWVALID;
	input [4:0] fib_7_s_axi_control_AWADDR;
	output wire fib_7_s_axi_control_WREADY;
	input fib_7_s_axi_control_WVALID;
	input [31:0] fib_7_s_axi_control_WDATA;
	input [3:0] fib_7_s_axi_control_WSTRB;
	input fib_7_s_axi_control_BREADY;
	output wire fib_7_s_axi_control_BVALID;
	output wire [1:0] fib_7_s_axi_control_BRESP;
	input fib_8_m_axi_gmem_ARREADY;
	output wire fib_8_m_axi_gmem_ARVALID;
	output wire fib_8_m_axi_gmem_ARID;
	output wire [63:0] fib_8_m_axi_gmem_ARADDR;
	output wire [7:0] fib_8_m_axi_gmem_ARLEN;
	output wire [2:0] fib_8_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_8_m_axi_gmem_ARBURST;
	output wire fib_8_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_8_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_8_m_axi_gmem_ARPROT;
	output wire [3:0] fib_8_m_axi_gmem_ARQOS;
	output wire [3:0] fib_8_m_axi_gmem_ARREGION;
	output wire fib_8_m_axi_gmem_ARUSER;
	output wire fib_8_m_axi_gmem_RREADY;
	input fib_8_m_axi_gmem_RVALID;
	input fib_8_m_axi_gmem_RID;
	input [63:0] fib_8_m_axi_gmem_RDATA;
	input [1:0] fib_8_m_axi_gmem_RRESP;
	input fib_8_m_axi_gmem_RLAST;
	input fib_8_m_axi_gmem_RUSER;
	input fib_8_m_axi_gmem_AWREADY;
	output wire fib_8_m_axi_gmem_AWVALID;
	output wire fib_8_m_axi_gmem_AWID;
	output wire [63:0] fib_8_m_axi_gmem_AWADDR;
	output wire [7:0] fib_8_m_axi_gmem_AWLEN;
	output wire [2:0] fib_8_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_8_m_axi_gmem_AWBURST;
	output wire fib_8_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_8_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_8_m_axi_gmem_AWPROT;
	output wire [3:0] fib_8_m_axi_gmem_AWQOS;
	output wire [3:0] fib_8_m_axi_gmem_AWREGION;
	output wire fib_8_m_axi_gmem_AWUSER;
	input fib_8_m_axi_gmem_WREADY;
	output wire fib_8_m_axi_gmem_WVALID;
	output wire [63:0] fib_8_m_axi_gmem_WDATA;
	output wire [7:0] fib_8_m_axi_gmem_WSTRB;
	output wire fib_8_m_axi_gmem_WLAST;
	output wire fib_8_m_axi_gmem_WUSER;
	output wire fib_8_m_axi_gmem_BREADY;
	input fib_8_m_axi_gmem_BVALID;
	input fib_8_m_axi_gmem_BID;
	input [1:0] fib_8_m_axi_gmem_BRESP;
	input fib_8_m_axi_gmem_BUSER;
	output wire fib_8_s_axi_control_ARREADY;
	input fib_8_s_axi_control_ARVALID;
	input [4:0] fib_8_s_axi_control_ARADDR;
	input fib_8_s_axi_control_RREADY;
	output wire fib_8_s_axi_control_RVALID;
	output wire [31:0] fib_8_s_axi_control_RDATA;
	output wire [1:0] fib_8_s_axi_control_RRESP;
	output wire fib_8_s_axi_control_AWREADY;
	input fib_8_s_axi_control_AWVALID;
	input [4:0] fib_8_s_axi_control_AWADDR;
	output wire fib_8_s_axi_control_WREADY;
	input fib_8_s_axi_control_WVALID;
	input [31:0] fib_8_s_axi_control_WDATA;
	input [3:0] fib_8_s_axi_control_WSTRB;
	input fib_8_s_axi_control_BREADY;
	output wire fib_8_s_axi_control_BVALID;
	output wire [1:0] fib_8_s_axi_control_BRESP;
	input fib_9_m_axi_gmem_ARREADY;
	output wire fib_9_m_axi_gmem_ARVALID;
	output wire fib_9_m_axi_gmem_ARID;
	output wire [63:0] fib_9_m_axi_gmem_ARADDR;
	output wire [7:0] fib_9_m_axi_gmem_ARLEN;
	output wire [2:0] fib_9_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_9_m_axi_gmem_ARBURST;
	output wire fib_9_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_9_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_9_m_axi_gmem_ARPROT;
	output wire [3:0] fib_9_m_axi_gmem_ARQOS;
	output wire [3:0] fib_9_m_axi_gmem_ARREGION;
	output wire fib_9_m_axi_gmem_ARUSER;
	output wire fib_9_m_axi_gmem_RREADY;
	input fib_9_m_axi_gmem_RVALID;
	input fib_9_m_axi_gmem_RID;
	input [63:0] fib_9_m_axi_gmem_RDATA;
	input [1:0] fib_9_m_axi_gmem_RRESP;
	input fib_9_m_axi_gmem_RLAST;
	input fib_9_m_axi_gmem_RUSER;
	input fib_9_m_axi_gmem_AWREADY;
	output wire fib_9_m_axi_gmem_AWVALID;
	output wire fib_9_m_axi_gmem_AWID;
	output wire [63:0] fib_9_m_axi_gmem_AWADDR;
	output wire [7:0] fib_9_m_axi_gmem_AWLEN;
	output wire [2:0] fib_9_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_9_m_axi_gmem_AWBURST;
	output wire fib_9_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_9_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_9_m_axi_gmem_AWPROT;
	output wire [3:0] fib_9_m_axi_gmem_AWQOS;
	output wire [3:0] fib_9_m_axi_gmem_AWREGION;
	output wire fib_9_m_axi_gmem_AWUSER;
	input fib_9_m_axi_gmem_WREADY;
	output wire fib_9_m_axi_gmem_WVALID;
	output wire [63:0] fib_9_m_axi_gmem_WDATA;
	output wire [7:0] fib_9_m_axi_gmem_WSTRB;
	output wire fib_9_m_axi_gmem_WLAST;
	output wire fib_9_m_axi_gmem_WUSER;
	output wire fib_9_m_axi_gmem_BREADY;
	input fib_9_m_axi_gmem_BVALID;
	input fib_9_m_axi_gmem_BID;
	input [1:0] fib_9_m_axi_gmem_BRESP;
	input fib_9_m_axi_gmem_BUSER;
	output wire fib_9_s_axi_control_ARREADY;
	input fib_9_s_axi_control_ARVALID;
	input [4:0] fib_9_s_axi_control_ARADDR;
	input fib_9_s_axi_control_RREADY;
	output wire fib_9_s_axi_control_RVALID;
	output wire [31:0] fib_9_s_axi_control_RDATA;
	output wire [1:0] fib_9_s_axi_control_RRESP;
	output wire fib_9_s_axi_control_AWREADY;
	input fib_9_s_axi_control_AWVALID;
	input [4:0] fib_9_s_axi_control_AWADDR;
	output wire fib_9_s_axi_control_WREADY;
	input fib_9_s_axi_control_WVALID;
	input [31:0] fib_9_s_axi_control_WDATA;
	input [3:0] fib_9_s_axi_control_WSTRB;
	input fib_9_s_axi_control_BREADY;
	output wire fib_9_s_axi_control_BVALID;
	output wire [1:0] fib_9_s_axi_control_BRESP;
	input fib_10_m_axi_gmem_ARREADY;
	output wire fib_10_m_axi_gmem_ARVALID;
	output wire fib_10_m_axi_gmem_ARID;
	output wire [63:0] fib_10_m_axi_gmem_ARADDR;
	output wire [7:0] fib_10_m_axi_gmem_ARLEN;
	output wire [2:0] fib_10_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_10_m_axi_gmem_ARBURST;
	output wire fib_10_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_10_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_10_m_axi_gmem_ARPROT;
	output wire [3:0] fib_10_m_axi_gmem_ARQOS;
	output wire [3:0] fib_10_m_axi_gmem_ARREGION;
	output wire fib_10_m_axi_gmem_ARUSER;
	output wire fib_10_m_axi_gmem_RREADY;
	input fib_10_m_axi_gmem_RVALID;
	input fib_10_m_axi_gmem_RID;
	input [63:0] fib_10_m_axi_gmem_RDATA;
	input [1:0] fib_10_m_axi_gmem_RRESP;
	input fib_10_m_axi_gmem_RLAST;
	input fib_10_m_axi_gmem_RUSER;
	input fib_10_m_axi_gmem_AWREADY;
	output wire fib_10_m_axi_gmem_AWVALID;
	output wire fib_10_m_axi_gmem_AWID;
	output wire [63:0] fib_10_m_axi_gmem_AWADDR;
	output wire [7:0] fib_10_m_axi_gmem_AWLEN;
	output wire [2:0] fib_10_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_10_m_axi_gmem_AWBURST;
	output wire fib_10_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_10_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_10_m_axi_gmem_AWPROT;
	output wire [3:0] fib_10_m_axi_gmem_AWQOS;
	output wire [3:0] fib_10_m_axi_gmem_AWREGION;
	output wire fib_10_m_axi_gmem_AWUSER;
	input fib_10_m_axi_gmem_WREADY;
	output wire fib_10_m_axi_gmem_WVALID;
	output wire [63:0] fib_10_m_axi_gmem_WDATA;
	output wire [7:0] fib_10_m_axi_gmem_WSTRB;
	output wire fib_10_m_axi_gmem_WLAST;
	output wire fib_10_m_axi_gmem_WUSER;
	output wire fib_10_m_axi_gmem_BREADY;
	input fib_10_m_axi_gmem_BVALID;
	input fib_10_m_axi_gmem_BID;
	input [1:0] fib_10_m_axi_gmem_BRESP;
	input fib_10_m_axi_gmem_BUSER;
	output wire fib_10_s_axi_control_ARREADY;
	input fib_10_s_axi_control_ARVALID;
	input [4:0] fib_10_s_axi_control_ARADDR;
	input fib_10_s_axi_control_RREADY;
	output wire fib_10_s_axi_control_RVALID;
	output wire [31:0] fib_10_s_axi_control_RDATA;
	output wire [1:0] fib_10_s_axi_control_RRESP;
	output wire fib_10_s_axi_control_AWREADY;
	input fib_10_s_axi_control_AWVALID;
	input [4:0] fib_10_s_axi_control_AWADDR;
	output wire fib_10_s_axi_control_WREADY;
	input fib_10_s_axi_control_WVALID;
	input [31:0] fib_10_s_axi_control_WDATA;
	input [3:0] fib_10_s_axi_control_WSTRB;
	input fib_10_s_axi_control_BREADY;
	output wire fib_10_s_axi_control_BVALID;
	output wire [1:0] fib_10_s_axi_control_BRESP;
	input fib_11_m_axi_gmem_ARREADY;
	output wire fib_11_m_axi_gmem_ARVALID;
	output wire fib_11_m_axi_gmem_ARID;
	output wire [63:0] fib_11_m_axi_gmem_ARADDR;
	output wire [7:0] fib_11_m_axi_gmem_ARLEN;
	output wire [2:0] fib_11_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_11_m_axi_gmem_ARBURST;
	output wire fib_11_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_11_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_11_m_axi_gmem_ARPROT;
	output wire [3:0] fib_11_m_axi_gmem_ARQOS;
	output wire [3:0] fib_11_m_axi_gmem_ARREGION;
	output wire fib_11_m_axi_gmem_ARUSER;
	output wire fib_11_m_axi_gmem_RREADY;
	input fib_11_m_axi_gmem_RVALID;
	input fib_11_m_axi_gmem_RID;
	input [63:0] fib_11_m_axi_gmem_RDATA;
	input [1:0] fib_11_m_axi_gmem_RRESP;
	input fib_11_m_axi_gmem_RLAST;
	input fib_11_m_axi_gmem_RUSER;
	input fib_11_m_axi_gmem_AWREADY;
	output wire fib_11_m_axi_gmem_AWVALID;
	output wire fib_11_m_axi_gmem_AWID;
	output wire [63:0] fib_11_m_axi_gmem_AWADDR;
	output wire [7:0] fib_11_m_axi_gmem_AWLEN;
	output wire [2:0] fib_11_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_11_m_axi_gmem_AWBURST;
	output wire fib_11_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_11_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_11_m_axi_gmem_AWPROT;
	output wire [3:0] fib_11_m_axi_gmem_AWQOS;
	output wire [3:0] fib_11_m_axi_gmem_AWREGION;
	output wire fib_11_m_axi_gmem_AWUSER;
	input fib_11_m_axi_gmem_WREADY;
	output wire fib_11_m_axi_gmem_WVALID;
	output wire [63:0] fib_11_m_axi_gmem_WDATA;
	output wire [7:0] fib_11_m_axi_gmem_WSTRB;
	output wire fib_11_m_axi_gmem_WLAST;
	output wire fib_11_m_axi_gmem_WUSER;
	output wire fib_11_m_axi_gmem_BREADY;
	input fib_11_m_axi_gmem_BVALID;
	input fib_11_m_axi_gmem_BID;
	input [1:0] fib_11_m_axi_gmem_BRESP;
	input fib_11_m_axi_gmem_BUSER;
	output wire fib_11_s_axi_control_ARREADY;
	input fib_11_s_axi_control_ARVALID;
	input [4:0] fib_11_s_axi_control_ARADDR;
	input fib_11_s_axi_control_RREADY;
	output wire fib_11_s_axi_control_RVALID;
	output wire [31:0] fib_11_s_axi_control_RDATA;
	output wire [1:0] fib_11_s_axi_control_RRESP;
	output wire fib_11_s_axi_control_AWREADY;
	input fib_11_s_axi_control_AWVALID;
	input [4:0] fib_11_s_axi_control_AWADDR;
	output wire fib_11_s_axi_control_WREADY;
	input fib_11_s_axi_control_WVALID;
	input [31:0] fib_11_s_axi_control_WDATA;
	input [3:0] fib_11_s_axi_control_WSTRB;
	input fib_11_s_axi_control_BREADY;
	output wire fib_11_s_axi_control_BVALID;
	output wire [1:0] fib_11_s_axi_control_BRESP;
	input fib_12_m_axi_gmem_ARREADY;
	output wire fib_12_m_axi_gmem_ARVALID;
	output wire fib_12_m_axi_gmem_ARID;
	output wire [63:0] fib_12_m_axi_gmem_ARADDR;
	output wire [7:0] fib_12_m_axi_gmem_ARLEN;
	output wire [2:0] fib_12_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_12_m_axi_gmem_ARBURST;
	output wire fib_12_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_12_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_12_m_axi_gmem_ARPROT;
	output wire [3:0] fib_12_m_axi_gmem_ARQOS;
	output wire [3:0] fib_12_m_axi_gmem_ARREGION;
	output wire fib_12_m_axi_gmem_ARUSER;
	output wire fib_12_m_axi_gmem_RREADY;
	input fib_12_m_axi_gmem_RVALID;
	input fib_12_m_axi_gmem_RID;
	input [63:0] fib_12_m_axi_gmem_RDATA;
	input [1:0] fib_12_m_axi_gmem_RRESP;
	input fib_12_m_axi_gmem_RLAST;
	input fib_12_m_axi_gmem_RUSER;
	input fib_12_m_axi_gmem_AWREADY;
	output wire fib_12_m_axi_gmem_AWVALID;
	output wire fib_12_m_axi_gmem_AWID;
	output wire [63:0] fib_12_m_axi_gmem_AWADDR;
	output wire [7:0] fib_12_m_axi_gmem_AWLEN;
	output wire [2:0] fib_12_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_12_m_axi_gmem_AWBURST;
	output wire fib_12_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_12_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_12_m_axi_gmem_AWPROT;
	output wire [3:0] fib_12_m_axi_gmem_AWQOS;
	output wire [3:0] fib_12_m_axi_gmem_AWREGION;
	output wire fib_12_m_axi_gmem_AWUSER;
	input fib_12_m_axi_gmem_WREADY;
	output wire fib_12_m_axi_gmem_WVALID;
	output wire [63:0] fib_12_m_axi_gmem_WDATA;
	output wire [7:0] fib_12_m_axi_gmem_WSTRB;
	output wire fib_12_m_axi_gmem_WLAST;
	output wire fib_12_m_axi_gmem_WUSER;
	output wire fib_12_m_axi_gmem_BREADY;
	input fib_12_m_axi_gmem_BVALID;
	input fib_12_m_axi_gmem_BID;
	input [1:0] fib_12_m_axi_gmem_BRESP;
	input fib_12_m_axi_gmem_BUSER;
	output wire fib_12_s_axi_control_ARREADY;
	input fib_12_s_axi_control_ARVALID;
	input [4:0] fib_12_s_axi_control_ARADDR;
	input fib_12_s_axi_control_RREADY;
	output wire fib_12_s_axi_control_RVALID;
	output wire [31:0] fib_12_s_axi_control_RDATA;
	output wire [1:0] fib_12_s_axi_control_RRESP;
	output wire fib_12_s_axi_control_AWREADY;
	input fib_12_s_axi_control_AWVALID;
	input [4:0] fib_12_s_axi_control_AWADDR;
	output wire fib_12_s_axi_control_WREADY;
	input fib_12_s_axi_control_WVALID;
	input [31:0] fib_12_s_axi_control_WDATA;
	input [3:0] fib_12_s_axi_control_WSTRB;
	input fib_12_s_axi_control_BREADY;
	output wire fib_12_s_axi_control_BVALID;
	output wire [1:0] fib_12_s_axi_control_BRESP;
	input fib_13_m_axi_gmem_ARREADY;
	output wire fib_13_m_axi_gmem_ARVALID;
	output wire fib_13_m_axi_gmem_ARID;
	output wire [63:0] fib_13_m_axi_gmem_ARADDR;
	output wire [7:0] fib_13_m_axi_gmem_ARLEN;
	output wire [2:0] fib_13_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_13_m_axi_gmem_ARBURST;
	output wire fib_13_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_13_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_13_m_axi_gmem_ARPROT;
	output wire [3:0] fib_13_m_axi_gmem_ARQOS;
	output wire [3:0] fib_13_m_axi_gmem_ARREGION;
	output wire fib_13_m_axi_gmem_ARUSER;
	output wire fib_13_m_axi_gmem_RREADY;
	input fib_13_m_axi_gmem_RVALID;
	input fib_13_m_axi_gmem_RID;
	input [63:0] fib_13_m_axi_gmem_RDATA;
	input [1:0] fib_13_m_axi_gmem_RRESP;
	input fib_13_m_axi_gmem_RLAST;
	input fib_13_m_axi_gmem_RUSER;
	input fib_13_m_axi_gmem_AWREADY;
	output wire fib_13_m_axi_gmem_AWVALID;
	output wire fib_13_m_axi_gmem_AWID;
	output wire [63:0] fib_13_m_axi_gmem_AWADDR;
	output wire [7:0] fib_13_m_axi_gmem_AWLEN;
	output wire [2:0] fib_13_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_13_m_axi_gmem_AWBURST;
	output wire fib_13_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_13_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_13_m_axi_gmem_AWPROT;
	output wire [3:0] fib_13_m_axi_gmem_AWQOS;
	output wire [3:0] fib_13_m_axi_gmem_AWREGION;
	output wire fib_13_m_axi_gmem_AWUSER;
	input fib_13_m_axi_gmem_WREADY;
	output wire fib_13_m_axi_gmem_WVALID;
	output wire [63:0] fib_13_m_axi_gmem_WDATA;
	output wire [7:0] fib_13_m_axi_gmem_WSTRB;
	output wire fib_13_m_axi_gmem_WLAST;
	output wire fib_13_m_axi_gmem_WUSER;
	output wire fib_13_m_axi_gmem_BREADY;
	input fib_13_m_axi_gmem_BVALID;
	input fib_13_m_axi_gmem_BID;
	input [1:0] fib_13_m_axi_gmem_BRESP;
	input fib_13_m_axi_gmem_BUSER;
	output wire fib_13_s_axi_control_ARREADY;
	input fib_13_s_axi_control_ARVALID;
	input [4:0] fib_13_s_axi_control_ARADDR;
	input fib_13_s_axi_control_RREADY;
	output wire fib_13_s_axi_control_RVALID;
	output wire [31:0] fib_13_s_axi_control_RDATA;
	output wire [1:0] fib_13_s_axi_control_RRESP;
	output wire fib_13_s_axi_control_AWREADY;
	input fib_13_s_axi_control_AWVALID;
	input [4:0] fib_13_s_axi_control_AWADDR;
	output wire fib_13_s_axi_control_WREADY;
	input fib_13_s_axi_control_WVALID;
	input [31:0] fib_13_s_axi_control_WDATA;
	input [3:0] fib_13_s_axi_control_WSTRB;
	input fib_13_s_axi_control_BREADY;
	output wire fib_13_s_axi_control_BVALID;
	output wire [1:0] fib_13_s_axi_control_BRESP;
	input fib_14_m_axi_gmem_ARREADY;
	output wire fib_14_m_axi_gmem_ARVALID;
	output wire fib_14_m_axi_gmem_ARID;
	output wire [63:0] fib_14_m_axi_gmem_ARADDR;
	output wire [7:0] fib_14_m_axi_gmem_ARLEN;
	output wire [2:0] fib_14_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_14_m_axi_gmem_ARBURST;
	output wire fib_14_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_14_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_14_m_axi_gmem_ARPROT;
	output wire [3:0] fib_14_m_axi_gmem_ARQOS;
	output wire [3:0] fib_14_m_axi_gmem_ARREGION;
	output wire fib_14_m_axi_gmem_ARUSER;
	output wire fib_14_m_axi_gmem_RREADY;
	input fib_14_m_axi_gmem_RVALID;
	input fib_14_m_axi_gmem_RID;
	input [63:0] fib_14_m_axi_gmem_RDATA;
	input [1:0] fib_14_m_axi_gmem_RRESP;
	input fib_14_m_axi_gmem_RLAST;
	input fib_14_m_axi_gmem_RUSER;
	input fib_14_m_axi_gmem_AWREADY;
	output wire fib_14_m_axi_gmem_AWVALID;
	output wire fib_14_m_axi_gmem_AWID;
	output wire [63:0] fib_14_m_axi_gmem_AWADDR;
	output wire [7:0] fib_14_m_axi_gmem_AWLEN;
	output wire [2:0] fib_14_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_14_m_axi_gmem_AWBURST;
	output wire fib_14_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_14_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_14_m_axi_gmem_AWPROT;
	output wire [3:0] fib_14_m_axi_gmem_AWQOS;
	output wire [3:0] fib_14_m_axi_gmem_AWREGION;
	output wire fib_14_m_axi_gmem_AWUSER;
	input fib_14_m_axi_gmem_WREADY;
	output wire fib_14_m_axi_gmem_WVALID;
	output wire [63:0] fib_14_m_axi_gmem_WDATA;
	output wire [7:0] fib_14_m_axi_gmem_WSTRB;
	output wire fib_14_m_axi_gmem_WLAST;
	output wire fib_14_m_axi_gmem_WUSER;
	output wire fib_14_m_axi_gmem_BREADY;
	input fib_14_m_axi_gmem_BVALID;
	input fib_14_m_axi_gmem_BID;
	input [1:0] fib_14_m_axi_gmem_BRESP;
	input fib_14_m_axi_gmem_BUSER;
	output wire fib_14_s_axi_control_ARREADY;
	input fib_14_s_axi_control_ARVALID;
	input [4:0] fib_14_s_axi_control_ARADDR;
	input fib_14_s_axi_control_RREADY;
	output wire fib_14_s_axi_control_RVALID;
	output wire [31:0] fib_14_s_axi_control_RDATA;
	output wire [1:0] fib_14_s_axi_control_RRESP;
	output wire fib_14_s_axi_control_AWREADY;
	input fib_14_s_axi_control_AWVALID;
	input [4:0] fib_14_s_axi_control_AWADDR;
	output wire fib_14_s_axi_control_WREADY;
	input fib_14_s_axi_control_WVALID;
	input [31:0] fib_14_s_axi_control_WDATA;
	input [3:0] fib_14_s_axi_control_WSTRB;
	input fib_14_s_axi_control_BREADY;
	output wire fib_14_s_axi_control_BVALID;
	output wire [1:0] fib_14_s_axi_control_BRESP;
	input fib_15_m_axi_gmem_ARREADY;
	output wire fib_15_m_axi_gmem_ARVALID;
	output wire fib_15_m_axi_gmem_ARID;
	output wire [63:0] fib_15_m_axi_gmem_ARADDR;
	output wire [7:0] fib_15_m_axi_gmem_ARLEN;
	output wire [2:0] fib_15_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_15_m_axi_gmem_ARBURST;
	output wire fib_15_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_15_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_15_m_axi_gmem_ARPROT;
	output wire [3:0] fib_15_m_axi_gmem_ARQOS;
	output wire [3:0] fib_15_m_axi_gmem_ARREGION;
	output wire fib_15_m_axi_gmem_ARUSER;
	output wire fib_15_m_axi_gmem_RREADY;
	input fib_15_m_axi_gmem_RVALID;
	input fib_15_m_axi_gmem_RID;
	input [63:0] fib_15_m_axi_gmem_RDATA;
	input [1:0] fib_15_m_axi_gmem_RRESP;
	input fib_15_m_axi_gmem_RLAST;
	input fib_15_m_axi_gmem_RUSER;
	input fib_15_m_axi_gmem_AWREADY;
	output wire fib_15_m_axi_gmem_AWVALID;
	output wire fib_15_m_axi_gmem_AWID;
	output wire [63:0] fib_15_m_axi_gmem_AWADDR;
	output wire [7:0] fib_15_m_axi_gmem_AWLEN;
	output wire [2:0] fib_15_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_15_m_axi_gmem_AWBURST;
	output wire fib_15_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_15_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_15_m_axi_gmem_AWPROT;
	output wire [3:0] fib_15_m_axi_gmem_AWQOS;
	output wire [3:0] fib_15_m_axi_gmem_AWREGION;
	output wire fib_15_m_axi_gmem_AWUSER;
	input fib_15_m_axi_gmem_WREADY;
	output wire fib_15_m_axi_gmem_WVALID;
	output wire [63:0] fib_15_m_axi_gmem_WDATA;
	output wire [7:0] fib_15_m_axi_gmem_WSTRB;
	output wire fib_15_m_axi_gmem_WLAST;
	output wire fib_15_m_axi_gmem_WUSER;
	output wire fib_15_m_axi_gmem_BREADY;
	input fib_15_m_axi_gmem_BVALID;
	input fib_15_m_axi_gmem_BID;
	input [1:0] fib_15_m_axi_gmem_BRESP;
	input fib_15_m_axi_gmem_BUSER;
	output wire fib_15_s_axi_control_ARREADY;
	input fib_15_s_axi_control_ARVALID;
	input [4:0] fib_15_s_axi_control_ARADDR;
	input fib_15_s_axi_control_RREADY;
	output wire fib_15_s_axi_control_RVALID;
	output wire [31:0] fib_15_s_axi_control_RDATA;
	output wire [1:0] fib_15_s_axi_control_RRESP;
	output wire fib_15_s_axi_control_AWREADY;
	input fib_15_s_axi_control_AWVALID;
	input [4:0] fib_15_s_axi_control_AWADDR;
	output wire fib_15_s_axi_control_WREADY;
	input fib_15_s_axi_control_WVALID;
	input [31:0] fib_15_s_axi_control_WDATA;
	input [3:0] fib_15_s_axi_control_WSTRB;
	input fib_15_s_axi_control_BREADY;
	output wire fib_15_s_axi_control_BVALID;
	output wire [1:0] fib_15_s_axi_control_BRESP;
	input fib_16_m_axi_gmem_ARREADY;
	output wire fib_16_m_axi_gmem_ARVALID;
	output wire fib_16_m_axi_gmem_ARID;
	output wire [63:0] fib_16_m_axi_gmem_ARADDR;
	output wire [7:0] fib_16_m_axi_gmem_ARLEN;
	output wire [2:0] fib_16_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_16_m_axi_gmem_ARBURST;
	output wire fib_16_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_16_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_16_m_axi_gmem_ARPROT;
	output wire [3:0] fib_16_m_axi_gmem_ARQOS;
	output wire [3:0] fib_16_m_axi_gmem_ARREGION;
	output wire fib_16_m_axi_gmem_ARUSER;
	output wire fib_16_m_axi_gmem_RREADY;
	input fib_16_m_axi_gmem_RVALID;
	input fib_16_m_axi_gmem_RID;
	input [63:0] fib_16_m_axi_gmem_RDATA;
	input [1:0] fib_16_m_axi_gmem_RRESP;
	input fib_16_m_axi_gmem_RLAST;
	input fib_16_m_axi_gmem_RUSER;
	input fib_16_m_axi_gmem_AWREADY;
	output wire fib_16_m_axi_gmem_AWVALID;
	output wire fib_16_m_axi_gmem_AWID;
	output wire [63:0] fib_16_m_axi_gmem_AWADDR;
	output wire [7:0] fib_16_m_axi_gmem_AWLEN;
	output wire [2:0] fib_16_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_16_m_axi_gmem_AWBURST;
	output wire fib_16_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_16_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_16_m_axi_gmem_AWPROT;
	output wire [3:0] fib_16_m_axi_gmem_AWQOS;
	output wire [3:0] fib_16_m_axi_gmem_AWREGION;
	output wire fib_16_m_axi_gmem_AWUSER;
	input fib_16_m_axi_gmem_WREADY;
	output wire fib_16_m_axi_gmem_WVALID;
	output wire [63:0] fib_16_m_axi_gmem_WDATA;
	output wire [7:0] fib_16_m_axi_gmem_WSTRB;
	output wire fib_16_m_axi_gmem_WLAST;
	output wire fib_16_m_axi_gmem_WUSER;
	output wire fib_16_m_axi_gmem_BREADY;
	input fib_16_m_axi_gmem_BVALID;
	input fib_16_m_axi_gmem_BID;
	input [1:0] fib_16_m_axi_gmem_BRESP;
	input fib_16_m_axi_gmem_BUSER;
	output wire fib_16_s_axi_control_ARREADY;
	input fib_16_s_axi_control_ARVALID;
	input [4:0] fib_16_s_axi_control_ARADDR;
	input fib_16_s_axi_control_RREADY;
	output wire fib_16_s_axi_control_RVALID;
	output wire [31:0] fib_16_s_axi_control_RDATA;
	output wire [1:0] fib_16_s_axi_control_RRESP;
	output wire fib_16_s_axi_control_AWREADY;
	input fib_16_s_axi_control_AWVALID;
	input [4:0] fib_16_s_axi_control_AWADDR;
	output wire fib_16_s_axi_control_WREADY;
	input fib_16_s_axi_control_WVALID;
	input [31:0] fib_16_s_axi_control_WDATA;
	input [3:0] fib_16_s_axi_control_WSTRB;
	input fib_16_s_axi_control_BREADY;
	output wire fib_16_s_axi_control_BVALID;
	output wire [1:0] fib_16_s_axi_control_BRESP;
	input fib_17_m_axi_gmem_ARREADY;
	output wire fib_17_m_axi_gmem_ARVALID;
	output wire fib_17_m_axi_gmem_ARID;
	output wire [63:0] fib_17_m_axi_gmem_ARADDR;
	output wire [7:0] fib_17_m_axi_gmem_ARLEN;
	output wire [2:0] fib_17_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_17_m_axi_gmem_ARBURST;
	output wire fib_17_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_17_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_17_m_axi_gmem_ARPROT;
	output wire [3:0] fib_17_m_axi_gmem_ARQOS;
	output wire [3:0] fib_17_m_axi_gmem_ARREGION;
	output wire fib_17_m_axi_gmem_ARUSER;
	output wire fib_17_m_axi_gmem_RREADY;
	input fib_17_m_axi_gmem_RVALID;
	input fib_17_m_axi_gmem_RID;
	input [63:0] fib_17_m_axi_gmem_RDATA;
	input [1:0] fib_17_m_axi_gmem_RRESP;
	input fib_17_m_axi_gmem_RLAST;
	input fib_17_m_axi_gmem_RUSER;
	input fib_17_m_axi_gmem_AWREADY;
	output wire fib_17_m_axi_gmem_AWVALID;
	output wire fib_17_m_axi_gmem_AWID;
	output wire [63:0] fib_17_m_axi_gmem_AWADDR;
	output wire [7:0] fib_17_m_axi_gmem_AWLEN;
	output wire [2:0] fib_17_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_17_m_axi_gmem_AWBURST;
	output wire fib_17_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_17_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_17_m_axi_gmem_AWPROT;
	output wire [3:0] fib_17_m_axi_gmem_AWQOS;
	output wire [3:0] fib_17_m_axi_gmem_AWREGION;
	output wire fib_17_m_axi_gmem_AWUSER;
	input fib_17_m_axi_gmem_WREADY;
	output wire fib_17_m_axi_gmem_WVALID;
	output wire [63:0] fib_17_m_axi_gmem_WDATA;
	output wire [7:0] fib_17_m_axi_gmem_WSTRB;
	output wire fib_17_m_axi_gmem_WLAST;
	output wire fib_17_m_axi_gmem_WUSER;
	output wire fib_17_m_axi_gmem_BREADY;
	input fib_17_m_axi_gmem_BVALID;
	input fib_17_m_axi_gmem_BID;
	input [1:0] fib_17_m_axi_gmem_BRESP;
	input fib_17_m_axi_gmem_BUSER;
	output wire fib_17_s_axi_control_ARREADY;
	input fib_17_s_axi_control_ARVALID;
	input [4:0] fib_17_s_axi_control_ARADDR;
	input fib_17_s_axi_control_RREADY;
	output wire fib_17_s_axi_control_RVALID;
	output wire [31:0] fib_17_s_axi_control_RDATA;
	output wire [1:0] fib_17_s_axi_control_RRESP;
	output wire fib_17_s_axi_control_AWREADY;
	input fib_17_s_axi_control_AWVALID;
	input [4:0] fib_17_s_axi_control_AWADDR;
	output wire fib_17_s_axi_control_WREADY;
	input fib_17_s_axi_control_WVALID;
	input [31:0] fib_17_s_axi_control_WDATA;
	input [3:0] fib_17_s_axi_control_WSTRB;
	input fib_17_s_axi_control_BREADY;
	output wire fib_17_s_axi_control_BVALID;
	output wire [1:0] fib_17_s_axi_control_BRESP;
	input fib_18_m_axi_gmem_ARREADY;
	output wire fib_18_m_axi_gmem_ARVALID;
	output wire fib_18_m_axi_gmem_ARID;
	output wire [63:0] fib_18_m_axi_gmem_ARADDR;
	output wire [7:0] fib_18_m_axi_gmem_ARLEN;
	output wire [2:0] fib_18_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_18_m_axi_gmem_ARBURST;
	output wire fib_18_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_18_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_18_m_axi_gmem_ARPROT;
	output wire [3:0] fib_18_m_axi_gmem_ARQOS;
	output wire [3:0] fib_18_m_axi_gmem_ARREGION;
	output wire fib_18_m_axi_gmem_ARUSER;
	output wire fib_18_m_axi_gmem_RREADY;
	input fib_18_m_axi_gmem_RVALID;
	input fib_18_m_axi_gmem_RID;
	input [63:0] fib_18_m_axi_gmem_RDATA;
	input [1:0] fib_18_m_axi_gmem_RRESP;
	input fib_18_m_axi_gmem_RLAST;
	input fib_18_m_axi_gmem_RUSER;
	input fib_18_m_axi_gmem_AWREADY;
	output wire fib_18_m_axi_gmem_AWVALID;
	output wire fib_18_m_axi_gmem_AWID;
	output wire [63:0] fib_18_m_axi_gmem_AWADDR;
	output wire [7:0] fib_18_m_axi_gmem_AWLEN;
	output wire [2:0] fib_18_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_18_m_axi_gmem_AWBURST;
	output wire fib_18_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_18_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_18_m_axi_gmem_AWPROT;
	output wire [3:0] fib_18_m_axi_gmem_AWQOS;
	output wire [3:0] fib_18_m_axi_gmem_AWREGION;
	output wire fib_18_m_axi_gmem_AWUSER;
	input fib_18_m_axi_gmem_WREADY;
	output wire fib_18_m_axi_gmem_WVALID;
	output wire [63:0] fib_18_m_axi_gmem_WDATA;
	output wire [7:0] fib_18_m_axi_gmem_WSTRB;
	output wire fib_18_m_axi_gmem_WLAST;
	output wire fib_18_m_axi_gmem_WUSER;
	output wire fib_18_m_axi_gmem_BREADY;
	input fib_18_m_axi_gmem_BVALID;
	input fib_18_m_axi_gmem_BID;
	input [1:0] fib_18_m_axi_gmem_BRESP;
	input fib_18_m_axi_gmem_BUSER;
	output wire fib_18_s_axi_control_ARREADY;
	input fib_18_s_axi_control_ARVALID;
	input [4:0] fib_18_s_axi_control_ARADDR;
	input fib_18_s_axi_control_RREADY;
	output wire fib_18_s_axi_control_RVALID;
	output wire [31:0] fib_18_s_axi_control_RDATA;
	output wire [1:0] fib_18_s_axi_control_RRESP;
	output wire fib_18_s_axi_control_AWREADY;
	input fib_18_s_axi_control_AWVALID;
	input [4:0] fib_18_s_axi_control_AWADDR;
	output wire fib_18_s_axi_control_WREADY;
	input fib_18_s_axi_control_WVALID;
	input [31:0] fib_18_s_axi_control_WDATA;
	input [3:0] fib_18_s_axi_control_WSTRB;
	input fib_18_s_axi_control_BREADY;
	output wire fib_18_s_axi_control_BVALID;
	output wire [1:0] fib_18_s_axi_control_BRESP;
	input fib_19_m_axi_gmem_ARREADY;
	output wire fib_19_m_axi_gmem_ARVALID;
	output wire fib_19_m_axi_gmem_ARID;
	output wire [63:0] fib_19_m_axi_gmem_ARADDR;
	output wire [7:0] fib_19_m_axi_gmem_ARLEN;
	output wire [2:0] fib_19_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_19_m_axi_gmem_ARBURST;
	output wire fib_19_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_19_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_19_m_axi_gmem_ARPROT;
	output wire [3:0] fib_19_m_axi_gmem_ARQOS;
	output wire [3:0] fib_19_m_axi_gmem_ARREGION;
	output wire fib_19_m_axi_gmem_ARUSER;
	output wire fib_19_m_axi_gmem_RREADY;
	input fib_19_m_axi_gmem_RVALID;
	input fib_19_m_axi_gmem_RID;
	input [63:0] fib_19_m_axi_gmem_RDATA;
	input [1:0] fib_19_m_axi_gmem_RRESP;
	input fib_19_m_axi_gmem_RLAST;
	input fib_19_m_axi_gmem_RUSER;
	input fib_19_m_axi_gmem_AWREADY;
	output wire fib_19_m_axi_gmem_AWVALID;
	output wire fib_19_m_axi_gmem_AWID;
	output wire [63:0] fib_19_m_axi_gmem_AWADDR;
	output wire [7:0] fib_19_m_axi_gmem_AWLEN;
	output wire [2:0] fib_19_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_19_m_axi_gmem_AWBURST;
	output wire fib_19_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_19_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_19_m_axi_gmem_AWPROT;
	output wire [3:0] fib_19_m_axi_gmem_AWQOS;
	output wire [3:0] fib_19_m_axi_gmem_AWREGION;
	output wire fib_19_m_axi_gmem_AWUSER;
	input fib_19_m_axi_gmem_WREADY;
	output wire fib_19_m_axi_gmem_WVALID;
	output wire [63:0] fib_19_m_axi_gmem_WDATA;
	output wire [7:0] fib_19_m_axi_gmem_WSTRB;
	output wire fib_19_m_axi_gmem_WLAST;
	output wire fib_19_m_axi_gmem_WUSER;
	output wire fib_19_m_axi_gmem_BREADY;
	input fib_19_m_axi_gmem_BVALID;
	input fib_19_m_axi_gmem_BID;
	input [1:0] fib_19_m_axi_gmem_BRESP;
	input fib_19_m_axi_gmem_BUSER;
	output wire fib_19_s_axi_control_ARREADY;
	input fib_19_s_axi_control_ARVALID;
	input [4:0] fib_19_s_axi_control_ARADDR;
	input fib_19_s_axi_control_RREADY;
	output wire fib_19_s_axi_control_RVALID;
	output wire [31:0] fib_19_s_axi_control_RDATA;
	output wire [1:0] fib_19_s_axi_control_RRESP;
	output wire fib_19_s_axi_control_AWREADY;
	input fib_19_s_axi_control_AWVALID;
	input [4:0] fib_19_s_axi_control_AWADDR;
	output wire fib_19_s_axi_control_WREADY;
	input fib_19_s_axi_control_WVALID;
	input [31:0] fib_19_s_axi_control_WDATA;
	input [3:0] fib_19_s_axi_control_WSTRB;
	input fib_19_s_axi_control_BREADY;
	output wire fib_19_s_axi_control_BVALID;
	output wire [1:0] fib_19_s_axi_control_BRESP;
	input fib_20_m_axi_gmem_ARREADY;
	output wire fib_20_m_axi_gmem_ARVALID;
	output wire fib_20_m_axi_gmem_ARID;
	output wire [63:0] fib_20_m_axi_gmem_ARADDR;
	output wire [7:0] fib_20_m_axi_gmem_ARLEN;
	output wire [2:0] fib_20_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_20_m_axi_gmem_ARBURST;
	output wire fib_20_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_20_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_20_m_axi_gmem_ARPROT;
	output wire [3:0] fib_20_m_axi_gmem_ARQOS;
	output wire [3:0] fib_20_m_axi_gmem_ARREGION;
	output wire fib_20_m_axi_gmem_ARUSER;
	output wire fib_20_m_axi_gmem_RREADY;
	input fib_20_m_axi_gmem_RVALID;
	input fib_20_m_axi_gmem_RID;
	input [63:0] fib_20_m_axi_gmem_RDATA;
	input [1:0] fib_20_m_axi_gmem_RRESP;
	input fib_20_m_axi_gmem_RLAST;
	input fib_20_m_axi_gmem_RUSER;
	input fib_20_m_axi_gmem_AWREADY;
	output wire fib_20_m_axi_gmem_AWVALID;
	output wire fib_20_m_axi_gmem_AWID;
	output wire [63:0] fib_20_m_axi_gmem_AWADDR;
	output wire [7:0] fib_20_m_axi_gmem_AWLEN;
	output wire [2:0] fib_20_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_20_m_axi_gmem_AWBURST;
	output wire fib_20_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_20_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_20_m_axi_gmem_AWPROT;
	output wire [3:0] fib_20_m_axi_gmem_AWQOS;
	output wire [3:0] fib_20_m_axi_gmem_AWREGION;
	output wire fib_20_m_axi_gmem_AWUSER;
	input fib_20_m_axi_gmem_WREADY;
	output wire fib_20_m_axi_gmem_WVALID;
	output wire [63:0] fib_20_m_axi_gmem_WDATA;
	output wire [7:0] fib_20_m_axi_gmem_WSTRB;
	output wire fib_20_m_axi_gmem_WLAST;
	output wire fib_20_m_axi_gmem_WUSER;
	output wire fib_20_m_axi_gmem_BREADY;
	input fib_20_m_axi_gmem_BVALID;
	input fib_20_m_axi_gmem_BID;
	input [1:0] fib_20_m_axi_gmem_BRESP;
	input fib_20_m_axi_gmem_BUSER;
	output wire fib_20_s_axi_control_ARREADY;
	input fib_20_s_axi_control_ARVALID;
	input [4:0] fib_20_s_axi_control_ARADDR;
	input fib_20_s_axi_control_RREADY;
	output wire fib_20_s_axi_control_RVALID;
	output wire [31:0] fib_20_s_axi_control_RDATA;
	output wire [1:0] fib_20_s_axi_control_RRESP;
	output wire fib_20_s_axi_control_AWREADY;
	input fib_20_s_axi_control_AWVALID;
	input [4:0] fib_20_s_axi_control_AWADDR;
	output wire fib_20_s_axi_control_WREADY;
	input fib_20_s_axi_control_WVALID;
	input [31:0] fib_20_s_axi_control_WDATA;
	input [3:0] fib_20_s_axi_control_WSTRB;
	input fib_20_s_axi_control_BREADY;
	output wire fib_20_s_axi_control_BVALID;
	output wire [1:0] fib_20_s_axi_control_BRESP;
	input fib_21_m_axi_gmem_ARREADY;
	output wire fib_21_m_axi_gmem_ARVALID;
	output wire fib_21_m_axi_gmem_ARID;
	output wire [63:0] fib_21_m_axi_gmem_ARADDR;
	output wire [7:0] fib_21_m_axi_gmem_ARLEN;
	output wire [2:0] fib_21_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_21_m_axi_gmem_ARBURST;
	output wire fib_21_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_21_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_21_m_axi_gmem_ARPROT;
	output wire [3:0] fib_21_m_axi_gmem_ARQOS;
	output wire [3:0] fib_21_m_axi_gmem_ARREGION;
	output wire fib_21_m_axi_gmem_ARUSER;
	output wire fib_21_m_axi_gmem_RREADY;
	input fib_21_m_axi_gmem_RVALID;
	input fib_21_m_axi_gmem_RID;
	input [63:0] fib_21_m_axi_gmem_RDATA;
	input [1:0] fib_21_m_axi_gmem_RRESP;
	input fib_21_m_axi_gmem_RLAST;
	input fib_21_m_axi_gmem_RUSER;
	input fib_21_m_axi_gmem_AWREADY;
	output wire fib_21_m_axi_gmem_AWVALID;
	output wire fib_21_m_axi_gmem_AWID;
	output wire [63:0] fib_21_m_axi_gmem_AWADDR;
	output wire [7:0] fib_21_m_axi_gmem_AWLEN;
	output wire [2:0] fib_21_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_21_m_axi_gmem_AWBURST;
	output wire fib_21_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_21_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_21_m_axi_gmem_AWPROT;
	output wire [3:0] fib_21_m_axi_gmem_AWQOS;
	output wire [3:0] fib_21_m_axi_gmem_AWREGION;
	output wire fib_21_m_axi_gmem_AWUSER;
	input fib_21_m_axi_gmem_WREADY;
	output wire fib_21_m_axi_gmem_WVALID;
	output wire [63:0] fib_21_m_axi_gmem_WDATA;
	output wire [7:0] fib_21_m_axi_gmem_WSTRB;
	output wire fib_21_m_axi_gmem_WLAST;
	output wire fib_21_m_axi_gmem_WUSER;
	output wire fib_21_m_axi_gmem_BREADY;
	input fib_21_m_axi_gmem_BVALID;
	input fib_21_m_axi_gmem_BID;
	input [1:0] fib_21_m_axi_gmem_BRESP;
	input fib_21_m_axi_gmem_BUSER;
	output wire fib_21_s_axi_control_ARREADY;
	input fib_21_s_axi_control_ARVALID;
	input [4:0] fib_21_s_axi_control_ARADDR;
	input fib_21_s_axi_control_RREADY;
	output wire fib_21_s_axi_control_RVALID;
	output wire [31:0] fib_21_s_axi_control_RDATA;
	output wire [1:0] fib_21_s_axi_control_RRESP;
	output wire fib_21_s_axi_control_AWREADY;
	input fib_21_s_axi_control_AWVALID;
	input [4:0] fib_21_s_axi_control_AWADDR;
	output wire fib_21_s_axi_control_WREADY;
	input fib_21_s_axi_control_WVALID;
	input [31:0] fib_21_s_axi_control_WDATA;
	input [3:0] fib_21_s_axi_control_WSTRB;
	input fib_21_s_axi_control_BREADY;
	output wire fib_21_s_axi_control_BVALID;
	output wire [1:0] fib_21_s_axi_control_BRESP;
	input fib_22_m_axi_gmem_ARREADY;
	output wire fib_22_m_axi_gmem_ARVALID;
	output wire fib_22_m_axi_gmem_ARID;
	output wire [63:0] fib_22_m_axi_gmem_ARADDR;
	output wire [7:0] fib_22_m_axi_gmem_ARLEN;
	output wire [2:0] fib_22_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_22_m_axi_gmem_ARBURST;
	output wire fib_22_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_22_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_22_m_axi_gmem_ARPROT;
	output wire [3:0] fib_22_m_axi_gmem_ARQOS;
	output wire [3:0] fib_22_m_axi_gmem_ARREGION;
	output wire fib_22_m_axi_gmem_ARUSER;
	output wire fib_22_m_axi_gmem_RREADY;
	input fib_22_m_axi_gmem_RVALID;
	input fib_22_m_axi_gmem_RID;
	input [63:0] fib_22_m_axi_gmem_RDATA;
	input [1:0] fib_22_m_axi_gmem_RRESP;
	input fib_22_m_axi_gmem_RLAST;
	input fib_22_m_axi_gmem_RUSER;
	input fib_22_m_axi_gmem_AWREADY;
	output wire fib_22_m_axi_gmem_AWVALID;
	output wire fib_22_m_axi_gmem_AWID;
	output wire [63:0] fib_22_m_axi_gmem_AWADDR;
	output wire [7:0] fib_22_m_axi_gmem_AWLEN;
	output wire [2:0] fib_22_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_22_m_axi_gmem_AWBURST;
	output wire fib_22_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_22_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_22_m_axi_gmem_AWPROT;
	output wire [3:0] fib_22_m_axi_gmem_AWQOS;
	output wire [3:0] fib_22_m_axi_gmem_AWREGION;
	output wire fib_22_m_axi_gmem_AWUSER;
	input fib_22_m_axi_gmem_WREADY;
	output wire fib_22_m_axi_gmem_WVALID;
	output wire [63:0] fib_22_m_axi_gmem_WDATA;
	output wire [7:0] fib_22_m_axi_gmem_WSTRB;
	output wire fib_22_m_axi_gmem_WLAST;
	output wire fib_22_m_axi_gmem_WUSER;
	output wire fib_22_m_axi_gmem_BREADY;
	input fib_22_m_axi_gmem_BVALID;
	input fib_22_m_axi_gmem_BID;
	input [1:0] fib_22_m_axi_gmem_BRESP;
	input fib_22_m_axi_gmem_BUSER;
	output wire fib_22_s_axi_control_ARREADY;
	input fib_22_s_axi_control_ARVALID;
	input [4:0] fib_22_s_axi_control_ARADDR;
	input fib_22_s_axi_control_RREADY;
	output wire fib_22_s_axi_control_RVALID;
	output wire [31:0] fib_22_s_axi_control_RDATA;
	output wire [1:0] fib_22_s_axi_control_RRESP;
	output wire fib_22_s_axi_control_AWREADY;
	input fib_22_s_axi_control_AWVALID;
	input [4:0] fib_22_s_axi_control_AWADDR;
	output wire fib_22_s_axi_control_WREADY;
	input fib_22_s_axi_control_WVALID;
	input [31:0] fib_22_s_axi_control_WDATA;
	input [3:0] fib_22_s_axi_control_WSTRB;
	input fib_22_s_axi_control_BREADY;
	output wire fib_22_s_axi_control_BVALID;
	output wire [1:0] fib_22_s_axi_control_BRESP;
	input fib_23_m_axi_gmem_ARREADY;
	output wire fib_23_m_axi_gmem_ARVALID;
	output wire fib_23_m_axi_gmem_ARID;
	output wire [63:0] fib_23_m_axi_gmem_ARADDR;
	output wire [7:0] fib_23_m_axi_gmem_ARLEN;
	output wire [2:0] fib_23_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_23_m_axi_gmem_ARBURST;
	output wire fib_23_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_23_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_23_m_axi_gmem_ARPROT;
	output wire [3:0] fib_23_m_axi_gmem_ARQOS;
	output wire [3:0] fib_23_m_axi_gmem_ARREGION;
	output wire fib_23_m_axi_gmem_ARUSER;
	output wire fib_23_m_axi_gmem_RREADY;
	input fib_23_m_axi_gmem_RVALID;
	input fib_23_m_axi_gmem_RID;
	input [63:0] fib_23_m_axi_gmem_RDATA;
	input [1:0] fib_23_m_axi_gmem_RRESP;
	input fib_23_m_axi_gmem_RLAST;
	input fib_23_m_axi_gmem_RUSER;
	input fib_23_m_axi_gmem_AWREADY;
	output wire fib_23_m_axi_gmem_AWVALID;
	output wire fib_23_m_axi_gmem_AWID;
	output wire [63:0] fib_23_m_axi_gmem_AWADDR;
	output wire [7:0] fib_23_m_axi_gmem_AWLEN;
	output wire [2:0] fib_23_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_23_m_axi_gmem_AWBURST;
	output wire fib_23_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_23_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_23_m_axi_gmem_AWPROT;
	output wire [3:0] fib_23_m_axi_gmem_AWQOS;
	output wire [3:0] fib_23_m_axi_gmem_AWREGION;
	output wire fib_23_m_axi_gmem_AWUSER;
	input fib_23_m_axi_gmem_WREADY;
	output wire fib_23_m_axi_gmem_WVALID;
	output wire [63:0] fib_23_m_axi_gmem_WDATA;
	output wire [7:0] fib_23_m_axi_gmem_WSTRB;
	output wire fib_23_m_axi_gmem_WLAST;
	output wire fib_23_m_axi_gmem_WUSER;
	output wire fib_23_m_axi_gmem_BREADY;
	input fib_23_m_axi_gmem_BVALID;
	input fib_23_m_axi_gmem_BID;
	input [1:0] fib_23_m_axi_gmem_BRESP;
	input fib_23_m_axi_gmem_BUSER;
	output wire fib_23_s_axi_control_ARREADY;
	input fib_23_s_axi_control_ARVALID;
	input [4:0] fib_23_s_axi_control_ARADDR;
	input fib_23_s_axi_control_RREADY;
	output wire fib_23_s_axi_control_RVALID;
	output wire [31:0] fib_23_s_axi_control_RDATA;
	output wire [1:0] fib_23_s_axi_control_RRESP;
	output wire fib_23_s_axi_control_AWREADY;
	input fib_23_s_axi_control_AWVALID;
	input [4:0] fib_23_s_axi_control_AWADDR;
	output wire fib_23_s_axi_control_WREADY;
	input fib_23_s_axi_control_WVALID;
	input [31:0] fib_23_s_axi_control_WDATA;
	input [3:0] fib_23_s_axi_control_WSTRB;
	input fib_23_s_axi_control_BREADY;
	output wire fib_23_s_axi_control_BVALID;
	output wire [1:0] fib_23_s_axi_control_BRESP;
	input fib_24_m_axi_gmem_ARREADY;
	output wire fib_24_m_axi_gmem_ARVALID;
	output wire fib_24_m_axi_gmem_ARID;
	output wire [63:0] fib_24_m_axi_gmem_ARADDR;
	output wire [7:0] fib_24_m_axi_gmem_ARLEN;
	output wire [2:0] fib_24_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_24_m_axi_gmem_ARBURST;
	output wire fib_24_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_24_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_24_m_axi_gmem_ARPROT;
	output wire [3:0] fib_24_m_axi_gmem_ARQOS;
	output wire [3:0] fib_24_m_axi_gmem_ARREGION;
	output wire fib_24_m_axi_gmem_ARUSER;
	output wire fib_24_m_axi_gmem_RREADY;
	input fib_24_m_axi_gmem_RVALID;
	input fib_24_m_axi_gmem_RID;
	input [63:0] fib_24_m_axi_gmem_RDATA;
	input [1:0] fib_24_m_axi_gmem_RRESP;
	input fib_24_m_axi_gmem_RLAST;
	input fib_24_m_axi_gmem_RUSER;
	input fib_24_m_axi_gmem_AWREADY;
	output wire fib_24_m_axi_gmem_AWVALID;
	output wire fib_24_m_axi_gmem_AWID;
	output wire [63:0] fib_24_m_axi_gmem_AWADDR;
	output wire [7:0] fib_24_m_axi_gmem_AWLEN;
	output wire [2:0] fib_24_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_24_m_axi_gmem_AWBURST;
	output wire fib_24_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_24_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_24_m_axi_gmem_AWPROT;
	output wire [3:0] fib_24_m_axi_gmem_AWQOS;
	output wire [3:0] fib_24_m_axi_gmem_AWREGION;
	output wire fib_24_m_axi_gmem_AWUSER;
	input fib_24_m_axi_gmem_WREADY;
	output wire fib_24_m_axi_gmem_WVALID;
	output wire [63:0] fib_24_m_axi_gmem_WDATA;
	output wire [7:0] fib_24_m_axi_gmem_WSTRB;
	output wire fib_24_m_axi_gmem_WLAST;
	output wire fib_24_m_axi_gmem_WUSER;
	output wire fib_24_m_axi_gmem_BREADY;
	input fib_24_m_axi_gmem_BVALID;
	input fib_24_m_axi_gmem_BID;
	input [1:0] fib_24_m_axi_gmem_BRESP;
	input fib_24_m_axi_gmem_BUSER;
	output wire fib_24_s_axi_control_ARREADY;
	input fib_24_s_axi_control_ARVALID;
	input [4:0] fib_24_s_axi_control_ARADDR;
	input fib_24_s_axi_control_RREADY;
	output wire fib_24_s_axi_control_RVALID;
	output wire [31:0] fib_24_s_axi_control_RDATA;
	output wire [1:0] fib_24_s_axi_control_RRESP;
	output wire fib_24_s_axi_control_AWREADY;
	input fib_24_s_axi_control_AWVALID;
	input [4:0] fib_24_s_axi_control_AWADDR;
	output wire fib_24_s_axi_control_WREADY;
	input fib_24_s_axi_control_WVALID;
	input [31:0] fib_24_s_axi_control_WDATA;
	input [3:0] fib_24_s_axi_control_WSTRB;
	input fib_24_s_axi_control_BREADY;
	output wire fib_24_s_axi_control_BVALID;
	output wire [1:0] fib_24_s_axi_control_BRESP;
	input fib_25_m_axi_gmem_ARREADY;
	output wire fib_25_m_axi_gmem_ARVALID;
	output wire fib_25_m_axi_gmem_ARID;
	output wire [63:0] fib_25_m_axi_gmem_ARADDR;
	output wire [7:0] fib_25_m_axi_gmem_ARLEN;
	output wire [2:0] fib_25_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_25_m_axi_gmem_ARBURST;
	output wire fib_25_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_25_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_25_m_axi_gmem_ARPROT;
	output wire [3:0] fib_25_m_axi_gmem_ARQOS;
	output wire [3:0] fib_25_m_axi_gmem_ARREGION;
	output wire fib_25_m_axi_gmem_ARUSER;
	output wire fib_25_m_axi_gmem_RREADY;
	input fib_25_m_axi_gmem_RVALID;
	input fib_25_m_axi_gmem_RID;
	input [63:0] fib_25_m_axi_gmem_RDATA;
	input [1:0] fib_25_m_axi_gmem_RRESP;
	input fib_25_m_axi_gmem_RLAST;
	input fib_25_m_axi_gmem_RUSER;
	input fib_25_m_axi_gmem_AWREADY;
	output wire fib_25_m_axi_gmem_AWVALID;
	output wire fib_25_m_axi_gmem_AWID;
	output wire [63:0] fib_25_m_axi_gmem_AWADDR;
	output wire [7:0] fib_25_m_axi_gmem_AWLEN;
	output wire [2:0] fib_25_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_25_m_axi_gmem_AWBURST;
	output wire fib_25_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_25_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_25_m_axi_gmem_AWPROT;
	output wire [3:0] fib_25_m_axi_gmem_AWQOS;
	output wire [3:0] fib_25_m_axi_gmem_AWREGION;
	output wire fib_25_m_axi_gmem_AWUSER;
	input fib_25_m_axi_gmem_WREADY;
	output wire fib_25_m_axi_gmem_WVALID;
	output wire [63:0] fib_25_m_axi_gmem_WDATA;
	output wire [7:0] fib_25_m_axi_gmem_WSTRB;
	output wire fib_25_m_axi_gmem_WLAST;
	output wire fib_25_m_axi_gmem_WUSER;
	output wire fib_25_m_axi_gmem_BREADY;
	input fib_25_m_axi_gmem_BVALID;
	input fib_25_m_axi_gmem_BID;
	input [1:0] fib_25_m_axi_gmem_BRESP;
	input fib_25_m_axi_gmem_BUSER;
	output wire fib_25_s_axi_control_ARREADY;
	input fib_25_s_axi_control_ARVALID;
	input [4:0] fib_25_s_axi_control_ARADDR;
	input fib_25_s_axi_control_RREADY;
	output wire fib_25_s_axi_control_RVALID;
	output wire [31:0] fib_25_s_axi_control_RDATA;
	output wire [1:0] fib_25_s_axi_control_RRESP;
	output wire fib_25_s_axi_control_AWREADY;
	input fib_25_s_axi_control_AWVALID;
	input [4:0] fib_25_s_axi_control_AWADDR;
	output wire fib_25_s_axi_control_WREADY;
	input fib_25_s_axi_control_WVALID;
	input [31:0] fib_25_s_axi_control_WDATA;
	input [3:0] fib_25_s_axi_control_WSTRB;
	input fib_25_s_axi_control_BREADY;
	output wire fib_25_s_axi_control_BVALID;
	output wire [1:0] fib_25_s_axi_control_BRESP;
	input fib_26_m_axi_gmem_ARREADY;
	output wire fib_26_m_axi_gmem_ARVALID;
	output wire fib_26_m_axi_gmem_ARID;
	output wire [63:0] fib_26_m_axi_gmem_ARADDR;
	output wire [7:0] fib_26_m_axi_gmem_ARLEN;
	output wire [2:0] fib_26_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_26_m_axi_gmem_ARBURST;
	output wire fib_26_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_26_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_26_m_axi_gmem_ARPROT;
	output wire [3:0] fib_26_m_axi_gmem_ARQOS;
	output wire [3:0] fib_26_m_axi_gmem_ARREGION;
	output wire fib_26_m_axi_gmem_ARUSER;
	output wire fib_26_m_axi_gmem_RREADY;
	input fib_26_m_axi_gmem_RVALID;
	input fib_26_m_axi_gmem_RID;
	input [63:0] fib_26_m_axi_gmem_RDATA;
	input [1:0] fib_26_m_axi_gmem_RRESP;
	input fib_26_m_axi_gmem_RLAST;
	input fib_26_m_axi_gmem_RUSER;
	input fib_26_m_axi_gmem_AWREADY;
	output wire fib_26_m_axi_gmem_AWVALID;
	output wire fib_26_m_axi_gmem_AWID;
	output wire [63:0] fib_26_m_axi_gmem_AWADDR;
	output wire [7:0] fib_26_m_axi_gmem_AWLEN;
	output wire [2:0] fib_26_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_26_m_axi_gmem_AWBURST;
	output wire fib_26_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_26_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_26_m_axi_gmem_AWPROT;
	output wire [3:0] fib_26_m_axi_gmem_AWQOS;
	output wire [3:0] fib_26_m_axi_gmem_AWREGION;
	output wire fib_26_m_axi_gmem_AWUSER;
	input fib_26_m_axi_gmem_WREADY;
	output wire fib_26_m_axi_gmem_WVALID;
	output wire [63:0] fib_26_m_axi_gmem_WDATA;
	output wire [7:0] fib_26_m_axi_gmem_WSTRB;
	output wire fib_26_m_axi_gmem_WLAST;
	output wire fib_26_m_axi_gmem_WUSER;
	output wire fib_26_m_axi_gmem_BREADY;
	input fib_26_m_axi_gmem_BVALID;
	input fib_26_m_axi_gmem_BID;
	input [1:0] fib_26_m_axi_gmem_BRESP;
	input fib_26_m_axi_gmem_BUSER;
	output wire fib_26_s_axi_control_ARREADY;
	input fib_26_s_axi_control_ARVALID;
	input [4:0] fib_26_s_axi_control_ARADDR;
	input fib_26_s_axi_control_RREADY;
	output wire fib_26_s_axi_control_RVALID;
	output wire [31:0] fib_26_s_axi_control_RDATA;
	output wire [1:0] fib_26_s_axi_control_RRESP;
	output wire fib_26_s_axi_control_AWREADY;
	input fib_26_s_axi_control_AWVALID;
	input [4:0] fib_26_s_axi_control_AWADDR;
	output wire fib_26_s_axi_control_WREADY;
	input fib_26_s_axi_control_WVALID;
	input [31:0] fib_26_s_axi_control_WDATA;
	input [3:0] fib_26_s_axi_control_WSTRB;
	input fib_26_s_axi_control_BREADY;
	output wire fib_26_s_axi_control_BVALID;
	output wire [1:0] fib_26_s_axi_control_BRESP;
	input fib_27_m_axi_gmem_ARREADY;
	output wire fib_27_m_axi_gmem_ARVALID;
	output wire fib_27_m_axi_gmem_ARID;
	output wire [63:0] fib_27_m_axi_gmem_ARADDR;
	output wire [7:0] fib_27_m_axi_gmem_ARLEN;
	output wire [2:0] fib_27_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_27_m_axi_gmem_ARBURST;
	output wire fib_27_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_27_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_27_m_axi_gmem_ARPROT;
	output wire [3:0] fib_27_m_axi_gmem_ARQOS;
	output wire [3:0] fib_27_m_axi_gmem_ARREGION;
	output wire fib_27_m_axi_gmem_ARUSER;
	output wire fib_27_m_axi_gmem_RREADY;
	input fib_27_m_axi_gmem_RVALID;
	input fib_27_m_axi_gmem_RID;
	input [63:0] fib_27_m_axi_gmem_RDATA;
	input [1:0] fib_27_m_axi_gmem_RRESP;
	input fib_27_m_axi_gmem_RLAST;
	input fib_27_m_axi_gmem_RUSER;
	input fib_27_m_axi_gmem_AWREADY;
	output wire fib_27_m_axi_gmem_AWVALID;
	output wire fib_27_m_axi_gmem_AWID;
	output wire [63:0] fib_27_m_axi_gmem_AWADDR;
	output wire [7:0] fib_27_m_axi_gmem_AWLEN;
	output wire [2:0] fib_27_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_27_m_axi_gmem_AWBURST;
	output wire fib_27_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_27_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_27_m_axi_gmem_AWPROT;
	output wire [3:0] fib_27_m_axi_gmem_AWQOS;
	output wire [3:0] fib_27_m_axi_gmem_AWREGION;
	output wire fib_27_m_axi_gmem_AWUSER;
	input fib_27_m_axi_gmem_WREADY;
	output wire fib_27_m_axi_gmem_WVALID;
	output wire [63:0] fib_27_m_axi_gmem_WDATA;
	output wire [7:0] fib_27_m_axi_gmem_WSTRB;
	output wire fib_27_m_axi_gmem_WLAST;
	output wire fib_27_m_axi_gmem_WUSER;
	output wire fib_27_m_axi_gmem_BREADY;
	input fib_27_m_axi_gmem_BVALID;
	input fib_27_m_axi_gmem_BID;
	input [1:0] fib_27_m_axi_gmem_BRESP;
	input fib_27_m_axi_gmem_BUSER;
	output wire fib_27_s_axi_control_ARREADY;
	input fib_27_s_axi_control_ARVALID;
	input [4:0] fib_27_s_axi_control_ARADDR;
	input fib_27_s_axi_control_RREADY;
	output wire fib_27_s_axi_control_RVALID;
	output wire [31:0] fib_27_s_axi_control_RDATA;
	output wire [1:0] fib_27_s_axi_control_RRESP;
	output wire fib_27_s_axi_control_AWREADY;
	input fib_27_s_axi_control_AWVALID;
	input [4:0] fib_27_s_axi_control_AWADDR;
	output wire fib_27_s_axi_control_WREADY;
	input fib_27_s_axi_control_WVALID;
	input [31:0] fib_27_s_axi_control_WDATA;
	input [3:0] fib_27_s_axi_control_WSTRB;
	input fib_27_s_axi_control_BREADY;
	output wire fib_27_s_axi_control_BVALID;
	output wire [1:0] fib_27_s_axi_control_BRESP;
	input fib_28_m_axi_gmem_ARREADY;
	output wire fib_28_m_axi_gmem_ARVALID;
	output wire fib_28_m_axi_gmem_ARID;
	output wire [63:0] fib_28_m_axi_gmem_ARADDR;
	output wire [7:0] fib_28_m_axi_gmem_ARLEN;
	output wire [2:0] fib_28_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_28_m_axi_gmem_ARBURST;
	output wire fib_28_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_28_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_28_m_axi_gmem_ARPROT;
	output wire [3:0] fib_28_m_axi_gmem_ARQOS;
	output wire [3:0] fib_28_m_axi_gmem_ARREGION;
	output wire fib_28_m_axi_gmem_ARUSER;
	output wire fib_28_m_axi_gmem_RREADY;
	input fib_28_m_axi_gmem_RVALID;
	input fib_28_m_axi_gmem_RID;
	input [63:0] fib_28_m_axi_gmem_RDATA;
	input [1:0] fib_28_m_axi_gmem_RRESP;
	input fib_28_m_axi_gmem_RLAST;
	input fib_28_m_axi_gmem_RUSER;
	input fib_28_m_axi_gmem_AWREADY;
	output wire fib_28_m_axi_gmem_AWVALID;
	output wire fib_28_m_axi_gmem_AWID;
	output wire [63:0] fib_28_m_axi_gmem_AWADDR;
	output wire [7:0] fib_28_m_axi_gmem_AWLEN;
	output wire [2:0] fib_28_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_28_m_axi_gmem_AWBURST;
	output wire fib_28_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_28_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_28_m_axi_gmem_AWPROT;
	output wire [3:0] fib_28_m_axi_gmem_AWQOS;
	output wire [3:0] fib_28_m_axi_gmem_AWREGION;
	output wire fib_28_m_axi_gmem_AWUSER;
	input fib_28_m_axi_gmem_WREADY;
	output wire fib_28_m_axi_gmem_WVALID;
	output wire [63:0] fib_28_m_axi_gmem_WDATA;
	output wire [7:0] fib_28_m_axi_gmem_WSTRB;
	output wire fib_28_m_axi_gmem_WLAST;
	output wire fib_28_m_axi_gmem_WUSER;
	output wire fib_28_m_axi_gmem_BREADY;
	input fib_28_m_axi_gmem_BVALID;
	input fib_28_m_axi_gmem_BID;
	input [1:0] fib_28_m_axi_gmem_BRESP;
	input fib_28_m_axi_gmem_BUSER;
	output wire fib_28_s_axi_control_ARREADY;
	input fib_28_s_axi_control_ARVALID;
	input [4:0] fib_28_s_axi_control_ARADDR;
	input fib_28_s_axi_control_RREADY;
	output wire fib_28_s_axi_control_RVALID;
	output wire [31:0] fib_28_s_axi_control_RDATA;
	output wire [1:0] fib_28_s_axi_control_RRESP;
	output wire fib_28_s_axi_control_AWREADY;
	input fib_28_s_axi_control_AWVALID;
	input [4:0] fib_28_s_axi_control_AWADDR;
	output wire fib_28_s_axi_control_WREADY;
	input fib_28_s_axi_control_WVALID;
	input [31:0] fib_28_s_axi_control_WDATA;
	input [3:0] fib_28_s_axi_control_WSTRB;
	input fib_28_s_axi_control_BREADY;
	output wire fib_28_s_axi_control_BVALID;
	output wire [1:0] fib_28_s_axi_control_BRESP;
	input fib_29_m_axi_gmem_ARREADY;
	output wire fib_29_m_axi_gmem_ARVALID;
	output wire fib_29_m_axi_gmem_ARID;
	output wire [63:0] fib_29_m_axi_gmem_ARADDR;
	output wire [7:0] fib_29_m_axi_gmem_ARLEN;
	output wire [2:0] fib_29_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_29_m_axi_gmem_ARBURST;
	output wire fib_29_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_29_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_29_m_axi_gmem_ARPROT;
	output wire [3:0] fib_29_m_axi_gmem_ARQOS;
	output wire [3:0] fib_29_m_axi_gmem_ARREGION;
	output wire fib_29_m_axi_gmem_ARUSER;
	output wire fib_29_m_axi_gmem_RREADY;
	input fib_29_m_axi_gmem_RVALID;
	input fib_29_m_axi_gmem_RID;
	input [63:0] fib_29_m_axi_gmem_RDATA;
	input [1:0] fib_29_m_axi_gmem_RRESP;
	input fib_29_m_axi_gmem_RLAST;
	input fib_29_m_axi_gmem_RUSER;
	input fib_29_m_axi_gmem_AWREADY;
	output wire fib_29_m_axi_gmem_AWVALID;
	output wire fib_29_m_axi_gmem_AWID;
	output wire [63:0] fib_29_m_axi_gmem_AWADDR;
	output wire [7:0] fib_29_m_axi_gmem_AWLEN;
	output wire [2:0] fib_29_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_29_m_axi_gmem_AWBURST;
	output wire fib_29_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_29_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_29_m_axi_gmem_AWPROT;
	output wire [3:0] fib_29_m_axi_gmem_AWQOS;
	output wire [3:0] fib_29_m_axi_gmem_AWREGION;
	output wire fib_29_m_axi_gmem_AWUSER;
	input fib_29_m_axi_gmem_WREADY;
	output wire fib_29_m_axi_gmem_WVALID;
	output wire [63:0] fib_29_m_axi_gmem_WDATA;
	output wire [7:0] fib_29_m_axi_gmem_WSTRB;
	output wire fib_29_m_axi_gmem_WLAST;
	output wire fib_29_m_axi_gmem_WUSER;
	output wire fib_29_m_axi_gmem_BREADY;
	input fib_29_m_axi_gmem_BVALID;
	input fib_29_m_axi_gmem_BID;
	input [1:0] fib_29_m_axi_gmem_BRESP;
	input fib_29_m_axi_gmem_BUSER;
	output wire fib_29_s_axi_control_ARREADY;
	input fib_29_s_axi_control_ARVALID;
	input [4:0] fib_29_s_axi_control_ARADDR;
	input fib_29_s_axi_control_RREADY;
	output wire fib_29_s_axi_control_RVALID;
	output wire [31:0] fib_29_s_axi_control_RDATA;
	output wire [1:0] fib_29_s_axi_control_RRESP;
	output wire fib_29_s_axi_control_AWREADY;
	input fib_29_s_axi_control_AWVALID;
	input [4:0] fib_29_s_axi_control_AWADDR;
	output wire fib_29_s_axi_control_WREADY;
	input fib_29_s_axi_control_WVALID;
	input [31:0] fib_29_s_axi_control_WDATA;
	input [3:0] fib_29_s_axi_control_WSTRB;
	input fib_29_s_axi_control_BREADY;
	output wire fib_29_s_axi_control_BVALID;
	output wire [1:0] fib_29_s_axi_control_BRESP;
	input fib_30_m_axi_gmem_ARREADY;
	output wire fib_30_m_axi_gmem_ARVALID;
	output wire fib_30_m_axi_gmem_ARID;
	output wire [63:0] fib_30_m_axi_gmem_ARADDR;
	output wire [7:0] fib_30_m_axi_gmem_ARLEN;
	output wire [2:0] fib_30_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_30_m_axi_gmem_ARBURST;
	output wire fib_30_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_30_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_30_m_axi_gmem_ARPROT;
	output wire [3:0] fib_30_m_axi_gmem_ARQOS;
	output wire [3:0] fib_30_m_axi_gmem_ARREGION;
	output wire fib_30_m_axi_gmem_ARUSER;
	output wire fib_30_m_axi_gmem_RREADY;
	input fib_30_m_axi_gmem_RVALID;
	input fib_30_m_axi_gmem_RID;
	input [63:0] fib_30_m_axi_gmem_RDATA;
	input [1:0] fib_30_m_axi_gmem_RRESP;
	input fib_30_m_axi_gmem_RLAST;
	input fib_30_m_axi_gmem_RUSER;
	input fib_30_m_axi_gmem_AWREADY;
	output wire fib_30_m_axi_gmem_AWVALID;
	output wire fib_30_m_axi_gmem_AWID;
	output wire [63:0] fib_30_m_axi_gmem_AWADDR;
	output wire [7:0] fib_30_m_axi_gmem_AWLEN;
	output wire [2:0] fib_30_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_30_m_axi_gmem_AWBURST;
	output wire fib_30_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_30_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_30_m_axi_gmem_AWPROT;
	output wire [3:0] fib_30_m_axi_gmem_AWQOS;
	output wire [3:0] fib_30_m_axi_gmem_AWREGION;
	output wire fib_30_m_axi_gmem_AWUSER;
	input fib_30_m_axi_gmem_WREADY;
	output wire fib_30_m_axi_gmem_WVALID;
	output wire [63:0] fib_30_m_axi_gmem_WDATA;
	output wire [7:0] fib_30_m_axi_gmem_WSTRB;
	output wire fib_30_m_axi_gmem_WLAST;
	output wire fib_30_m_axi_gmem_WUSER;
	output wire fib_30_m_axi_gmem_BREADY;
	input fib_30_m_axi_gmem_BVALID;
	input fib_30_m_axi_gmem_BID;
	input [1:0] fib_30_m_axi_gmem_BRESP;
	input fib_30_m_axi_gmem_BUSER;
	output wire fib_30_s_axi_control_ARREADY;
	input fib_30_s_axi_control_ARVALID;
	input [4:0] fib_30_s_axi_control_ARADDR;
	input fib_30_s_axi_control_RREADY;
	output wire fib_30_s_axi_control_RVALID;
	output wire [31:0] fib_30_s_axi_control_RDATA;
	output wire [1:0] fib_30_s_axi_control_RRESP;
	output wire fib_30_s_axi_control_AWREADY;
	input fib_30_s_axi_control_AWVALID;
	input [4:0] fib_30_s_axi_control_AWADDR;
	output wire fib_30_s_axi_control_WREADY;
	input fib_30_s_axi_control_WVALID;
	input [31:0] fib_30_s_axi_control_WDATA;
	input [3:0] fib_30_s_axi_control_WSTRB;
	input fib_30_s_axi_control_BREADY;
	output wire fib_30_s_axi_control_BVALID;
	output wire [1:0] fib_30_s_axi_control_BRESP;
	input fib_31_m_axi_gmem_ARREADY;
	output wire fib_31_m_axi_gmem_ARVALID;
	output wire fib_31_m_axi_gmem_ARID;
	output wire [63:0] fib_31_m_axi_gmem_ARADDR;
	output wire [7:0] fib_31_m_axi_gmem_ARLEN;
	output wire [2:0] fib_31_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_31_m_axi_gmem_ARBURST;
	output wire fib_31_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_31_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_31_m_axi_gmem_ARPROT;
	output wire [3:0] fib_31_m_axi_gmem_ARQOS;
	output wire [3:0] fib_31_m_axi_gmem_ARREGION;
	output wire fib_31_m_axi_gmem_ARUSER;
	output wire fib_31_m_axi_gmem_RREADY;
	input fib_31_m_axi_gmem_RVALID;
	input fib_31_m_axi_gmem_RID;
	input [63:0] fib_31_m_axi_gmem_RDATA;
	input [1:0] fib_31_m_axi_gmem_RRESP;
	input fib_31_m_axi_gmem_RLAST;
	input fib_31_m_axi_gmem_RUSER;
	input fib_31_m_axi_gmem_AWREADY;
	output wire fib_31_m_axi_gmem_AWVALID;
	output wire fib_31_m_axi_gmem_AWID;
	output wire [63:0] fib_31_m_axi_gmem_AWADDR;
	output wire [7:0] fib_31_m_axi_gmem_AWLEN;
	output wire [2:0] fib_31_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_31_m_axi_gmem_AWBURST;
	output wire fib_31_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_31_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_31_m_axi_gmem_AWPROT;
	output wire [3:0] fib_31_m_axi_gmem_AWQOS;
	output wire [3:0] fib_31_m_axi_gmem_AWREGION;
	output wire fib_31_m_axi_gmem_AWUSER;
	input fib_31_m_axi_gmem_WREADY;
	output wire fib_31_m_axi_gmem_WVALID;
	output wire [63:0] fib_31_m_axi_gmem_WDATA;
	output wire [7:0] fib_31_m_axi_gmem_WSTRB;
	output wire fib_31_m_axi_gmem_WLAST;
	output wire fib_31_m_axi_gmem_WUSER;
	output wire fib_31_m_axi_gmem_BREADY;
	input fib_31_m_axi_gmem_BVALID;
	input fib_31_m_axi_gmem_BID;
	input [1:0] fib_31_m_axi_gmem_BRESP;
	input fib_31_m_axi_gmem_BUSER;
	output wire fib_31_s_axi_control_ARREADY;
	input fib_31_s_axi_control_ARVALID;
	input [4:0] fib_31_s_axi_control_ARADDR;
	input fib_31_s_axi_control_RREADY;
	output wire fib_31_s_axi_control_RVALID;
	output wire [31:0] fib_31_s_axi_control_RDATA;
	output wire [1:0] fib_31_s_axi_control_RRESP;
	output wire fib_31_s_axi_control_AWREADY;
	input fib_31_s_axi_control_AWVALID;
	input [4:0] fib_31_s_axi_control_AWADDR;
	output wire fib_31_s_axi_control_WREADY;
	input fib_31_s_axi_control_WVALID;
	input [31:0] fib_31_s_axi_control_WDATA;
	input [3:0] fib_31_s_axi_control_WSTRB;
	input fib_31_s_axi_control_BREADY;
	output wire fib_31_s_axi_control_BVALID;
	output wire [1:0] fib_31_s_axi_control_BRESP;
	input fib_32_m_axi_gmem_ARREADY;
	output wire fib_32_m_axi_gmem_ARVALID;
	output wire fib_32_m_axi_gmem_ARID;
	output wire [63:0] fib_32_m_axi_gmem_ARADDR;
	output wire [7:0] fib_32_m_axi_gmem_ARLEN;
	output wire [2:0] fib_32_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_32_m_axi_gmem_ARBURST;
	output wire fib_32_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_32_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_32_m_axi_gmem_ARPROT;
	output wire [3:0] fib_32_m_axi_gmem_ARQOS;
	output wire [3:0] fib_32_m_axi_gmem_ARREGION;
	output wire fib_32_m_axi_gmem_ARUSER;
	output wire fib_32_m_axi_gmem_RREADY;
	input fib_32_m_axi_gmem_RVALID;
	input fib_32_m_axi_gmem_RID;
	input [63:0] fib_32_m_axi_gmem_RDATA;
	input [1:0] fib_32_m_axi_gmem_RRESP;
	input fib_32_m_axi_gmem_RLAST;
	input fib_32_m_axi_gmem_RUSER;
	input fib_32_m_axi_gmem_AWREADY;
	output wire fib_32_m_axi_gmem_AWVALID;
	output wire fib_32_m_axi_gmem_AWID;
	output wire [63:0] fib_32_m_axi_gmem_AWADDR;
	output wire [7:0] fib_32_m_axi_gmem_AWLEN;
	output wire [2:0] fib_32_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_32_m_axi_gmem_AWBURST;
	output wire fib_32_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_32_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_32_m_axi_gmem_AWPROT;
	output wire [3:0] fib_32_m_axi_gmem_AWQOS;
	output wire [3:0] fib_32_m_axi_gmem_AWREGION;
	output wire fib_32_m_axi_gmem_AWUSER;
	input fib_32_m_axi_gmem_WREADY;
	output wire fib_32_m_axi_gmem_WVALID;
	output wire [63:0] fib_32_m_axi_gmem_WDATA;
	output wire [7:0] fib_32_m_axi_gmem_WSTRB;
	output wire fib_32_m_axi_gmem_WLAST;
	output wire fib_32_m_axi_gmem_WUSER;
	output wire fib_32_m_axi_gmem_BREADY;
	input fib_32_m_axi_gmem_BVALID;
	input fib_32_m_axi_gmem_BID;
	input [1:0] fib_32_m_axi_gmem_BRESP;
	input fib_32_m_axi_gmem_BUSER;
	output wire fib_32_s_axi_control_ARREADY;
	input fib_32_s_axi_control_ARVALID;
	input [4:0] fib_32_s_axi_control_ARADDR;
	input fib_32_s_axi_control_RREADY;
	output wire fib_32_s_axi_control_RVALID;
	output wire [31:0] fib_32_s_axi_control_RDATA;
	output wire [1:0] fib_32_s_axi_control_RRESP;
	output wire fib_32_s_axi_control_AWREADY;
	input fib_32_s_axi_control_AWVALID;
	input [4:0] fib_32_s_axi_control_AWADDR;
	output wire fib_32_s_axi_control_WREADY;
	input fib_32_s_axi_control_WVALID;
	input [31:0] fib_32_s_axi_control_WDATA;
	input [3:0] fib_32_s_axi_control_WSTRB;
	input fib_32_s_axi_control_BREADY;
	output wire fib_32_s_axi_control_BVALID;
	output wire [1:0] fib_32_s_axi_control_BRESP;
	input fib_33_m_axi_gmem_ARREADY;
	output wire fib_33_m_axi_gmem_ARVALID;
	output wire fib_33_m_axi_gmem_ARID;
	output wire [63:0] fib_33_m_axi_gmem_ARADDR;
	output wire [7:0] fib_33_m_axi_gmem_ARLEN;
	output wire [2:0] fib_33_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_33_m_axi_gmem_ARBURST;
	output wire fib_33_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_33_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_33_m_axi_gmem_ARPROT;
	output wire [3:0] fib_33_m_axi_gmem_ARQOS;
	output wire [3:0] fib_33_m_axi_gmem_ARREGION;
	output wire fib_33_m_axi_gmem_ARUSER;
	output wire fib_33_m_axi_gmem_RREADY;
	input fib_33_m_axi_gmem_RVALID;
	input fib_33_m_axi_gmem_RID;
	input [63:0] fib_33_m_axi_gmem_RDATA;
	input [1:0] fib_33_m_axi_gmem_RRESP;
	input fib_33_m_axi_gmem_RLAST;
	input fib_33_m_axi_gmem_RUSER;
	input fib_33_m_axi_gmem_AWREADY;
	output wire fib_33_m_axi_gmem_AWVALID;
	output wire fib_33_m_axi_gmem_AWID;
	output wire [63:0] fib_33_m_axi_gmem_AWADDR;
	output wire [7:0] fib_33_m_axi_gmem_AWLEN;
	output wire [2:0] fib_33_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_33_m_axi_gmem_AWBURST;
	output wire fib_33_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_33_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_33_m_axi_gmem_AWPROT;
	output wire [3:0] fib_33_m_axi_gmem_AWQOS;
	output wire [3:0] fib_33_m_axi_gmem_AWREGION;
	output wire fib_33_m_axi_gmem_AWUSER;
	input fib_33_m_axi_gmem_WREADY;
	output wire fib_33_m_axi_gmem_WVALID;
	output wire [63:0] fib_33_m_axi_gmem_WDATA;
	output wire [7:0] fib_33_m_axi_gmem_WSTRB;
	output wire fib_33_m_axi_gmem_WLAST;
	output wire fib_33_m_axi_gmem_WUSER;
	output wire fib_33_m_axi_gmem_BREADY;
	input fib_33_m_axi_gmem_BVALID;
	input fib_33_m_axi_gmem_BID;
	input [1:0] fib_33_m_axi_gmem_BRESP;
	input fib_33_m_axi_gmem_BUSER;
	output wire fib_33_s_axi_control_ARREADY;
	input fib_33_s_axi_control_ARVALID;
	input [4:0] fib_33_s_axi_control_ARADDR;
	input fib_33_s_axi_control_RREADY;
	output wire fib_33_s_axi_control_RVALID;
	output wire [31:0] fib_33_s_axi_control_RDATA;
	output wire [1:0] fib_33_s_axi_control_RRESP;
	output wire fib_33_s_axi_control_AWREADY;
	input fib_33_s_axi_control_AWVALID;
	input [4:0] fib_33_s_axi_control_AWADDR;
	output wire fib_33_s_axi_control_WREADY;
	input fib_33_s_axi_control_WVALID;
	input [31:0] fib_33_s_axi_control_WDATA;
	input [3:0] fib_33_s_axi_control_WSTRB;
	input fib_33_s_axi_control_BREADY;
	output wire fib_33_s_axi_control_BVALID;
	output wire [1:0] fib_33_s_axi_control_BRESP;
	input fib_34_m_axi_gmem_ARREADY;
	output wire fib_34_m_axi_gmem_ARVALID;
	output wire fib_34_m_axi_gmem_ARID;
	output wire [63:0] fib_34_m_axi_gmem_ARADDR;
	output wire [7:0] fib_34_m_axi_gmem_ARLEN;
	output wire [2:0] fib_34_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_34_m_axi_gmem_ARBURST;
	output wire fib_34_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_34_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_34_m_axi_gmem_ARPROT;
	output wire [3:0] fib_34_m_axi_gmem_ARQOS;
	output wire [3:0] fib_34_m_axi_gmem_ARREGION;
	output wire fib_34_m_axi_gmem_ARUSER;
	output wire fib_34_m_axi_gmem_RREADY;
	input fib_34_m_axi_gmem_RVALID;
	input fib_34_m_axi_gmem_RID;
	input [63:0] fib_34_m_axi_gmem_RDATA;
	input [1:0] fib_34_m_axi_gmem_RRESP;
	input fib_34_m_axi_gmem_RLAST;
	input fib_34_m_axi_gmem_RUSER;
	input fib_34_m_axi_gmem_AWREADY;
	output wire fib_34_m_axi_gmem_AWVALID;
	output wire fib_34_m_axi_gmem_AWID;
	output wire [63:0] fib_34_m_axi_gmem_AWADDR;
	output wire [7:0] fib_34_m_axi_gmem_AWLEN;
	output wire [2:0] fib_34_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_34_m_axi_gmem_AWBURST;
	output wire fib_34_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_34_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_34_m_axi_gmem_AWPROT;
	output wire [3:0] fib_34_m_axi_gmem_AWQOS;
	output wire [3:0] fib_34_m_axi_gmem_AWREGION;
	output wire fib_34_m_axi_gmem_AWUSER;
	input fib_34_m_axi_gmem_WREADY;
	output wire fib_34_m_axi_gmem_WVALID;
	output wire [63:0] fib_34_m_axi_gmem_WDATA;
	output wire [7:0] fib_34_m_axi_gmem_WSTRB;
	output wire fib_34_m_axi_gmem_WLAST;
	output wire fib_34_m_axi_gmem_WUSER;
	output wire fib_34_m_axi_gmem_BREADY;
	input fib_34_m_axi_gmem_BVALID;
	input fib_34_m_axi_gmem_BID;
	input [1:0] fib_34_m_axi_gmem_BRESP;
	input fib_34_m_axi_gmem_BUSER;
	output wire fib_34_s_axi_control_ARREADY;
	input fib_34_s_axi_control_ARVALID;
	input [4:0] fib_34_s_axi_control_ARADDR;
	input fib_34_s_axi_control_RREADY;
	output wire fib_34_s_axi_control_RVALID;
	output wire [31:0] fib_34_s_axi_control_RDATA;
	output wire [1:0] fib_34_s_axi_control_RRESP;
	output wire fib_34_s_axi_control_AWREADY;
	input fib_34_s_axi_control_AWVALID;
	input [4:0] fib_34_s_axi_control_AWADDR;
	output wire fib_34_s_axi_control_WREADY;
	input fib_34_s_axi_control_WVALID;
	input [31:0] fib_34_s_axi_control_WDATA;
	input [3:0] fib_34_s_axi_control_WSTRB;
	input fib_34_s_axi_control_BREADY;
	output wire fib_34_s_axi_control_BVALID;
	output wire [1:0] fib_34_s_axi_control_BRESP;
	input fib_35_m_axi_gmem_ARREADY;
	output wire fib_35_m_axi_gmem_ARVALID;
	output wire fib_35_m_axi_gmem_ARID;
	output wire [63:0] fib_35_m_axi_gmem_ARADDR;
	output wire [7:0] fib_35_m_axi_gmem_ARLEN;
	output wire [2:0] fib_35_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_35_m_axi_gmem_ARBURST;
	output wire fib_35_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_35_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_35_m_axi_gmem_ARPROT;
	output wire [3:0] fib_35_m_axi_gmem_ARQOS;
	output wire [3:0] fib_35_m_axi_gmem_ARREGION;
	output wire fib_35_m_axi_gmem_ARUSER;
	output wire fib_35_m_axi_gmem_RREADY;
	input fib_35_m_axi_gmem_RVALID;
	input fib_35_m_axi_gmem_RID;
	input [63:0] fib_35_m_axi_gmem_RDATA;
	input [1:0] fib_35_m_axi_gmem_RRESP;
	input fib_35_m_axi_gmem_RLAST;
	input fib_35_m_axi_gmem_RUSER;
	input fib_35_m_axi_gmem_AWREADY;
	output wire fib_35_m_axi_gmem_AWVALID;
	output wire fib_35_m_axi_gmem_AWID;
	output wire [63:0] fib_35_m_axi_gmem_AWADDR;
	output wire [7:0] fib_35_m_axi_gmem_AWLEN;
	output wire [2:0] fib_35_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_35_m_axi_gmem_AWBURST;
	output wire fib_35_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_35_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_35_m_axi_gmem_AWPROT;
	output wire [3:0] fib_35_m_axi_gmem_AWQOS;
	output wire [3:0] fib_35_m_axi_gmem_AWREGION;
	output wire fib_35_m_axi_gmem_AWUSER;
	input fib_35_m_axi_gmem_WREADY;
	output wire fib_35_m_axi_gmem_WVALID;
	output wire [63:0] fib_35_m_axi_gmem_WDATA;
	output wire [7:0] fib_35_m_axi_gmem_WSTRB;
	output wire fib_35_m_axi_gmem_WLAST;
	output wire fib_35_m_axi_gmem_WUSER;
	output wire fib_35_m_axi_gmem_BREADY;
	input fib_35_m_axi_gmem_BVALID;
	input fib_35_m_axi_gmem_BID;
	input [1:0] fib_35_m_axi_gmem_BRESP;
	input fib_35_m_axi_gmem_BUSER;
	output wire fib_35_s_axi_control_ARREADY;
	input fib_35_s_axi_control_ARVALID;
	input [4:0] fib_35_s_axi_control_ARADDR;
	input fib_35_s_axi_control_RREADY;
	output wire fib_35_s_axi_control_RVALID;
	output wire [31:0] fib_35_s_axi_control_RDATA;
	output wire [1:0] fib_35_s_axi_control_RRESP;
	output wire fib_35_s_axi_control_AWREADY;
	input fib_35_s_axi_control_AWVALID;
	input [4:0] fib_35_s_axi_control_AWADDR;
	output wire fib_35_s_axi_control_WREADY;
	input fib_35_s_axi_control_WVALID;
	input [31:0] fib_35_s_axi_control_WDATA;
	input [3:0] fib_35_s_axi_control_WSTRB;
	input fib_35_s_axi_control_BREADY;
	output wire fib_35_s_axi_control_BVALID;
	output wire [1:0] fib_35_s_axi_control_BRESP;
	input fib_36_m_axi_gmem_ARREADY;
	output wire fib_36_m_axi_gmem_ARVALID;
	output wire fib_36_m_axi_gmem_ARID;
	output wire [63:0] fib_36_m_axi_gmem_ARADDR;
	output wire [7:0] fib_36_m_axi_gmem_ARLEN;
	output wire [2:0] fib_36_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_36_m_axi_gmem_ARBURST;
	output wire fib_36_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_36_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_36_m_axi_gmem_ARPROT;
	output wire [3:0] fib_36_m_axi_gmem_ARQOS;
	output wire [3:0] fib_36_m_axi_gmem_ARREGION;
	output wire fib_36_m_axi_gmem_ARUSER;
	output wire fib_36_m_axi_gmem_RREADY;
	input fib_36_m_axi_gmem_RVALID;
	input fib_36_m_axi_gmem_RID;
	input [63:0] fib_36_m_axi_gmem_RDATA;
	input [1:0] fib_36_m_axi_gmem_RRESP;
	input fib_36_m_axi_gmem_RLAST;
	input fib_36_m_axi_gmem_RUSER;
	input fib_36_m_axi_gmem_AWREADY;
	output wire fib_36_m_axi_gmem_AWVALID;
	output wire fib_36_m_axi_gmem_AWID;
	output wire [63:0] fib_36_m_axi_gmem_AWADDR;
	output wire [7:0] fib_36_m_axi_gmem_AWLEN;
	output wire [2:0] fib_36_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_36_m_axi_gmem_AWBURST;
	output wire fib_36_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_36_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_36_m_axi_gmem_AWPROT;
	output wire [3:0] fib_36_m_axi_gmem_AWQOS;
	output wire [3:0] fib_36_m_axi_gmem_AWREGION;
	output wire fib_36_m_axi_gmem_AWUSER;
	input fib_36_m_axi_gmem_WREADY;
	output wire fib_36_m_axi_gmem_WVALID;
	output wire [63:0] fib_36_m_axi_gmem_WDATA;
	output wire [7:0] fib_36_m_axi_gmem_WSTRB;
	output wire fib_36_m_axi_gmem_WLAST;
	output wire fib_36_m_axi_gmem_WUSER;
	output wire fib_36_m_axi_gmem_BREADY;
	input fib_36_m_axi_gmem_BVALID;
	input fib_36_m_axi_gmem_BID;
	input [1:0] fib_36_m_axi_gmem_BRESP;
	input fib_36_m_axi_gmem_BUSER;
	output wire fib_36_s_axi_control_ARREADY;
	input fib_36_s_axi_control_ARVALID;
	input [4:0] fib_36_s_axi_control_ARADDR;
	input fib_36_s_axi_control_RREADY;
	output wire fib_36_s_axi_control_RVALID;
	output wire [31:0] fib_36_s_axi_control_RDATA;
	output wire [1:0] fib_36_s_axi_control_RRESP;
	output wire fib_36_s_axi_control_AWREADY;
	input fib_36_s_axi_control_AWVALID;
	input [4:0] fib_36_s_axi_control_AWADDR;
	output wire fib_36_s_axi_control_WREADY;
	input fib_36_s_axi_control_WVALID;
	input [31:0] fib_36_s_axi_control_WDATA;
	input [3:0] fib_36_s_axi_control_WSTRB;
	input fib_36_s_axi_control_BREADY;
	output wire fib_36_s_axi_control_BVALID;
	output wire [1:0] fib_36_s_axi_control_BRESP;
	input fib_37_m_axi_gmem_ARREADY;
	output wire fib_37_m_axi_gmem_ARVALID;
	output wire fib_37_m_axi_gmem_ARID;
	output wire [63:0] fib_37_m_axi_gmem_ARADDR;
	output wire [7:0] fib_37_m_axi_gmem_ARLEN;
	output wire [2:0] fib_37_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_37_m_axi_gmem_ARBURST;
	output wire fib_37_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_37_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_37_m_axi_gmem_ARPROT;
	output wire [3:0] fib_37_m_axi_gmem_ARQOS;
	output wire [3:0] fib_37_m_axi_gmem_ARREGION;
	output wire fib_37_m_axi_gmem_ARUSER;
	output wire fib_37_m_axi_gmem_RREADY;
	input fib_37_m_axi_gmem_RVALID;
	input fib_37_m_axi_gmem_RID;
	input [63:0] fib_37_m_axi_gmem_RDATA;
	input [1:0] fib_37_m_axi_gmem_RRESP;
	input fib_37_m_axi_gmem_RLAST;
	input fib_37_m_axi_gmem_RUSER;
	input fib_37_m_axi_gmem_AWREADY;
	output wire fib_37_m_axi_gmem_AWVALID;
	output wire fib_37_m_axi_gmem_AWID;
	output wire [63:0] fib_37_m_axi_gmem_AWADDR;
	output wire [7:0] fib_37_m_axi_gmem_AWLEN;
	output wire [2:0] fib_37_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_37_m_axi_gmem_AWBURST;
	output wire fib_37_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_37_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_37_m_axi_gmem_AWPROT;
	output wire [3:0] fib_37_m_axi_gmem_AWQOS;
	output wire [3:0] fib_37_m_axi_gmem_AWREGION;
	output wire fib_37_m_axi_gmem_AWUSER;
	input fib_37_m_axi_gmem_WREADY;
	output wire fib_37_m_axi_gmem_WVALID;
	output wire [63:0] fib_37_m_axi_gmem_WDATA;
	output wire [7:0] fib_37_m_axi_gmem_WSTRB;
	output wire fib_37_m_axi_gmem_WLAST;
	output wire fib_37_m_axi_gmem_WUSER;
	output wire fib_37_m_axi_gmem_BREADY;
	input fib_37_m_axi_gmem_BVALID;
	input fib_37_m_axi_gmem_BID;
	input [1:0] fib_37_m_axi_gmem_BRESP;
	input fib_37_m_axi_gmem_BUSER;
	output wire fib_37_s_axi_control_ARREADY;
	input fib_37_s_axi_control_ARVALID;
	input [4:0] fib_37_s_axi_control_ARADDR;
	input fib_37_s_axi_control_RREADY;
	output wire fib_37_s_axi_control_RVALID;
	output wire [31:0] fib_37_s_axi_control_RDATA;
	output wire [1:0] fib_37_s_axi_control_RRESP;
	output wire fib_37_s_axi_control_AWREADY;
	input fib_37_s_axi_control_AWVALID;
	input [4:0] fib_37_s_axi_control_AWADDR;
	output wire fib_37_s_axi_control_WREADY;
	input fib_37_s_axi_control_WVALID;
	input [31:0] fib_37_s_axi_control_WDATA;
	input [3:0] fib_37_s_axi_control_WSTRB;
	input fib_37_s_axi_control_BREADY;
	output wire fib_37_s_axi_control_BVALID;
	output wire [1:0] fib_37_s_axi_control_BRESP;
	input fib_38_m_axi_gmem_ARREADY;
	output wire fib_38_m_axi_gmem_ARVALID;
	output wire fib_38_m_axi_gmem_ARID;
	output wire [63:0] fib_38_m_axi_gmem_ARADDR;
	output wire [7:0] fib_38_m_axi_gmem_ARLEN;
	output wire [2:0] fib_38_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_38_m_axi_gmem_ARBURST;
	output wire fib_38_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_38_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_38_m_axi_gmem_ARPROT;
	output wire [3:0] fib_38_m_axi_gmem_ARQOS;
	output wire [3:0] fib_38_m_axi_gmem_ARREGION;
	output wire fib_38_m_axi_gmem_ARUSER;
	output wire fib_38_m_axi_gmem_RREADY;
	input fib_38_m_axi_gmem_RVALID;
	input fib_38_m_axi_gmem_RID;
	input [63:0] fib_38_m_axi_gmem_RDATA;
	input [1:0] fib_38_m_axi_gmem_RRESP;
	input fib_38_m_axi_gmem_RLAST;
	input fib_38_m_axi_gmem_RUSER;
	input fib_38_m_axi_gmem_AWREADY;
	output wire fib_38_m_axi_gmem_AWVALID;
	output wire fib_38_m_axi_gmem_AWID;
	output wire [63:0] fib_38_m_axi_gmem_AWADDR;
	output wire [7:0] fib_38_m_axi_gmem_AWLEN;
	output wire [2:0] fib_38_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_38_m_axi_gmem_AWBURST;
	output wire fib_38_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_38_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_38_m_axi_gmem_AWPROT;
	output wire [3:0] fib_38_m_axi_gmem_AWQOS;
	output wire [3:0] fib_38_m_axi_gmem_AWREGION;
	output wire fib_38_m_axi_gmem_AWUSER;
	input fib_38_m_axi_gmem_WREADY;
	output wire fib_38_m_axi_gmem_WVALID;
	output wire [63:0] fib_38_m_axi_gmem_WDATA;
	output wire [7:0] fib_38_m_axi_gmem_WSTRB;
	output wire fib_38_m_axi_gmem_WLAST;
	output wire fib_38_m_axi_gmem_WUSER;
	output wire fib_38_m_axi_gmem_BREADY;
	input fib_38_m_axi_gmem_BVALID;
	input fib_38_m_axi_gmem_BID;
	input [1:0] fib_38_m_axi_gmem_BRESP;
	input fib_38_m_axi_gmem_BUSER;
	output wire fib_38_s_axi_control_ARREADY;
	input fib_38_s_axi_control_ARVALID;
	input [4:0] fib_38_s_axi_control_ARADDR;
	input fib_38_s_axi_control_RREADY;
	output wire fib_38_s_axi_control_RVALID;
	output wire [31:0] fib_38_s_axi_control_RDATA;
	output wire [1:0] fib_38_s_axi_control_RRESP;
	output wire fib_38_s_axi_control_AWREADY;
	input fib_38_s_axi_control_AWVALID;
	input [4:0] fib_38_s_axi_control_AWADDR;
	output wire fib_38_s_axi_control_WREADY;
	input fib_38_s_axi_control_WVALID;
	input [31:0] fib_38_s_axi_control_WDATA;
	input [3:0] fib_38_s_axi_control_WSTRB;
	input fib_38_s_axi_control_BREADY;
	output wire fib_38_s_axi_control_BVALID;
	output wire [1:0] fib_38_s_axi_control_BRESP;
	input fib_39_m_axi_gmem_ARREADY;
	output wire fib_39_m_axi_gmem_ARVALID;
	output wire fib_39_m_axi_gmem_ARID;
	output wire [63:0] fib_39_m_axi_gmem_ARADDR;
	output wire [7:0] fib_39_m_axi_gmem_ARLEN;
	output wire [2:0] fib_39_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_39_m_axi_gmem_ARBURST;
	output wire fib_39_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_39_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_39_m_axi_gmem_ARPROT;
	output wire [3:0] fib_39_m_axi_gmem_ARQOS;
	output wire [3:0] fib_39_m_axi_gmem_ARREGION;
	output wire fib_39_m_axi_gmem_ARUSER;
	output wire fib_39_m_axi_gmem_RREADY;
	input fib_39_m_axi_gmem_RVALID;
	input fib_39_m_axi_gmem_RID;
	input [63:0] fib_39_m_axi_gmem_RDATA;
	input [1:0] fib_39_m_axi_gmem_RRESP;
	input fib_39_m_axi_gmem_RLAST;
	input fib_39_m_axi_gmem_RUSER;
	input fib_39_m_axi_gmem_AWREADY;
	output wire fib_39_m_axi_gmem_AWVALID;
	output wire fib_39_m_axi_gmem_AWID;
	output wire [63:0] fib_39_m_axi_gmem_AWADDR;
	output wire [7:0] fib_39_m_axi_gmem_AWLEN;
	output wire [2:0] fib_39_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_39_m_axi_gmem_AWBURST;
	output wire fib_39_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_39_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_39_m_axi_gmem_AWPROT;
	output wire [3:0] fib_39_m_axi_gmem_AWQOS;
	output wire [3:0] fib_39_m_axi_gmem_AWREGION;
	output wire fib_39_m_axi_gmem_AWUSER;
	input fib_39_m_axi_gmem_WREADY;
	output wire fib_39_m_axi_gmem_WVALID;
	output wire [63:0] fib_39_m_axi_gmem_WDATA;
	output wire [7:0] fib_39_m_axi_gmem_WSTRB;
	output wire fib_39_m_axi_gmem_WLAST;
	output wire fib_39_m_axi_gmem_WUSER;
	output wire fib_39_m_axi_gmem_BREADY;
	input fib_39_m_axi_gmem_BVALID;
	input fib_39_m_axi_gmem_BID;
	input [1:0] fib_39_m_axi_gmem_BRESP;
	input fib_39_m_axi_gmem_BUSER;
	output wire fib_39_s_axi_control_ARREADY;
	input fib_39_s_axi_control_ARVALID;
	input [4:0] fib_39_s_axi_control_ARADDR;
	input fib_39_s_axi_control_RREADY;
	output wire fib_39_s_axi_control_RVALID;
	output wire [31:0] fib_39_s_axi_control_RDATA;
	output wire [1:0] fib_39_s_axi_control_RRESP;
	output wire fib_39_s_axi_control_AWREADY;
	input fib_39_s_axi_control_AWVALID;
	input [4:0] fib_39_s_axi_control_AWADDR;
	output wire fib_39_s_axi_control_WREADY;
	input fib_39_s_axi_control_WVALID;
	input [31:0] fib_39_s_axi_control_WDATA;
	input [3:0] fib_39_s_axi_control_WSTRB;
	input fib_39_s_axi_control_BREADY;
	output wire fib_39_s_axi_control_BVALID;
	output wire [1:0] fib_39_s_axi_control_BRESP;
	input fib_40_m_axi_gmem_ARREADY;
	output wire fib_40_m_axi_gmem_ARVALID;
	output wire fib_40_m_axi_gmem_ARID;
	output wire [63:0] fib_40_m_axi_gmem_ARADDR;
	output wire [7:0] fib_40_m_axi_gmem_ARLEN;
	output wire [2:0] fib_40_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_40_m_axi_gmem_ARBURST;
	output wire fib_40_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_40_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_40_m_axi_gmem_ARPROT;
	output wire [3:0] fib_40_m_axi_gmem_ARQOS;
	output wire [3:0] fib_40_m_axi_gmem_ARREGION;
	output wire fib_40_m_axi_gmem_ARUSER;
	output wire fib_40_m_axi_gmem_RREADY;
	input fib_40_m_axi_gmem_RVALID;
	input fib_40_m_axi_gmem_RID;
	input [63:0] fib_40_m_axi_gmem_RDATA;
	input [1:0] fib_40_m_axi_gmem_RRESP;
	input fib_40_m_axi_gmem_RLAST;
	input fib_40_m_axi_gmem_RUSER;
	input fib_40_m_axi_gmem_AWREADY;
	output wire fib_40_m_axi_gmem_AWVALID;
	output wire fib_40_m_axi_gmem_AWID;
	output wire [63:0] fib_40_m_axi_gmem_AWADDR;
	output wire [7:0] fib_40_m_axi_gmem_AWLEN;
	output wire [2:0] fib_40_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_40_m_axi_gmem_AWBURST;
	output wire fib_40_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_40_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_40_m_axi_gmem_AWPROT;
	output wire [3:0] fib_40_m_axi_gmem_AWQOS;
	output wire [3:0] fib_40_m_axi_gmem_AWREGION;
	output wire fib_40_m_axi_gmem_AWUSER;
	input fib_40_m_axi_gmem_WREADY;
	output wire fib_40_m_axi_gmem_WVALID;
	output wire [63:0] fib_40_m_axi_gmem_WDATA;
	output wire [7:0] fib_40_m_axi_gmem_WSTRB;
	output wire fib_40_m_axi_gmem_WLAST;
	output wire fib_40_m_axi_gmem_WUSER;
	output wire fib_40_m_axi_gmem_BREADY;
	input fib_40_m_axi_gmem_BVALID;
	input fib_40_m_axi_gmem_BID;
	input [1:0] fib_40_m_axi_gmem_BRESP;
	input fib_40_m_axi_gmem_BUSER;
	output wire fib_40_s_axi_control_ARREADY;
	input fib_40_s_axi_control_ARVALID;
	input [4:0] fib_40_s_axi_control_ARADDR;
	input fib_40_s_axi_control_RREADY;
	output wire fib_40_s_axi_control_RVALID;
	output wire [31:0] fib_40_s_axi_control_RDATA;
	output wire [1:0] fib_40_s_axi_control_RRESP;
	output wire fib_40_s_axi_control_AWREADY;
	input fib_40_s_axi_control_AWVALID;
	input [4:0] fib_40_s_axi_control_AWADDR;
	output wire fib_40_s_axi_control_WREADY;
	input fib_40_s_axi_control_WVALID;
	input [31:0] fib_40_s_axi_control_WDATA;
	input [3:0] fib_40_s_axi_control_WSTRB;
	input fib_40_s_axi_control_BREADY;
	output wire fib_40_s_axi_control_BVALID;
	output wire [1:0] fib_40_s_axi_control_BRESP;
	input fib_41_m_axi_gmem_ARREADY;
	output wire fib_41_m_axi_gmem_ARVALID;
	output wire fib_41_m_axi_gmem_ARID;
	output wire [63:0] fib_41_m_axi_gmem_ARADDR;
	output wire [7:0] fib_41_m_axi_gmem_ARLEN;
	output wire [2:0] fib_41_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_41_m_axi_gmem_ARBURST;
	output wire fib_41_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_41_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_41_m_axi_gmem_ARPROT;
	output wire [3:0] fib_41_m_axi_gmem_ARQOS;
	output wire [3:0] fib_41_m_axi_gmem_ARREGION;
	output wire fib_41_m_axi_gmem_ARUSER;
	output wire fib_41_m_axi_gmem_RREADY;
	input fib_41_m_axi_gmem_RVALID;
	input fib_41_m_axi_gmem_RID;
	input [63:0] fib_41_m_axi_gmem_RDATA;
	input [1:0] fib_41_m_axi_gmem_RRESP;
	input fib_41_m_axi_gmem_RLAST;
	input fib_41_m_axi_gmem_RUSER;
	input fib_41_m_axi_gmem_AWREADY;
	output wire fib_41_m_axi_gmem_AWVALID;
	output wire fib_41_m_axi_gmem_AWID;
	output wire [63:0] fib_41_m_axi_gmem_AWADDR;
	output wire [7:0] fib_41_m_axi_gmem_AWLEN;
	output wire [2:0] fib_41_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_41_m_axi_gmem_AWBURST;
	output wire fib_41_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_41_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_41_m_axi_gmem_AWPROT;
	output wire [3:0] fib_41_m_axi_gmem_AWQOS;
	output wire [3:0] fib_41_m_axi_gmem_AWREGION;
	output wire fib_41_m_axi_gmem_AWUSER;
	input fib_41_m_axi_gmem_WREADY;
	output wire fib_41_m_axi_gmem_WVALID;
	output wire [63:0] fib_41_m_axi_gmem_WDATA;
	output wire [7:0] fib_41_m_axi_gmem_WSTRB;
	output wire fib_41_m_axi_gmem_WLAST;
	output wire fib_41_m_axi_gmem_WUSER;
	output wire fib_41_m_axi_gmem_BREADY;
	input fib_41_m_axi_gmem_BVALID;
	input fib_41_m_axi_gmem_BID;
	input [1:0] fib_41_m_axi_gmem_BRESP;
	input fib_41_m_axi_gmem_BUSER;
	output wire fib_41_s_axi_control_ARREADY;
	input fib_41_s_axi_control_ARVALID;
	input [4:0] fib_41_s_axi_control_ARADDR;
	input fib_41_s_axi_control_RREADY;
	output wire fib_41_s_axi_control_RVALID;
	output wire [31:0] fib_41_s_axi_control_RDATA;
	output wire [1:0] fib_41_s_axi_control_RRESP;
	output wire fib_41_s_axi_control_AWREADY;
	input fib_41_s_axi_control_AWVALID;
	input [4:0] fib_41_s_axi_control_AWADDR;
	output wire fib_41_s_axi_control_WREADY;
	input fib_41_s_axi_control_WVALID;
	input [31:0] fib_41_s_axi_control_WDATA;
	input [3:0] fib_41_s_axi_control_WSTRB;
	input fib_41_s_axi_control_BREADY;
	output wire fib_41_s_axi_control_BVALID;
	output wire [1:0] fib_41_s_axi_control_BRESP;
	input fib_42_m_axi_gmem_ARREADY;
	output wire fib_42_m_axi_gmem_ARVALID;
	output wire fib_42_m_axi_gmem_ARID;
	output wire [63:0] fib_42_m_axi_gmem_ARADDR;
	output wire [7:0] fib_42_m_axi_gmem_ARLEN;
	output wire [2:0] fib_42_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_42_m_axi_gmem_ARBURST;
	output wire fib_42_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_42_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_42_m_axi_gmem_ARPROT;
	output wire [3:0] fib_42_m_axi_gmem_ARQOS;
	output wire [3:0] fib_42_m_axi_gmem_ARREGION;
	output wire fib_42_m_axi_gmem_ARUSER;
	output wire fib_42_m_axi_gmem_RREADY;
	input fib_42_m_axi_gmem_RVALID;
	input fib_42_m_axi_gmem_RID;
	input [63:0] fib_42_m_axi_gmem_RDATA;
	input [1:0] fib_42_m_axi_gmem_RRESP;
	input fib_42_m_axi_gmem_RLAST;
	input fib_42_m_axi_gmem_RUSER;
	input fib_42_m_axi_gmem_AWREADY;
	output wire fib_42_m_axi_gmem_AWVALID;
	output wire fib_42_m_axi_gmem_AWID;
	output wire [63:0] fib_42_m_axi_gmem_AWADDR;
	output wire [7:0] fib_42_m_axi_gmem_AWLEN;
	output wire [2:0] fib_42_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_42_m_axi_gmem_AWBURST;
	output wire fib_42_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_42_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_42_m_axi_gmem_AWPROT;
	output wire [3:0] fib_42_m_axi_gmem_AWQOS;
	output wire [3:0] fib_42_m_axi_gmem_AWREGION;
	output wire fib_42_m_axi_gmem_AWUSER;
	input fib_42_m_axi_gmem_WREADY;
	output wire fib_42_m_axi_gmem_WVALID;
	output wire [63:0] fib_42_m_axi_gmem_WDATA;
	output wire [7:0] fib_42_m_axi_gmem_WSTRB;
	output wire fib_42_m_axi_gmem_WLAST;
	output wire fib_42_m_axi_gmem_WUSER;
	output wire fib_42_m_axi_gmem_BREADY;
	input fib_42_m_axi_gmem_BVALID;
	input fib_42_m_axi_gmem_BID;
	input [1:0] fib_42_m_axi_gmem_BRESP;
	input fib_42_m_axi_gmem_BUSER;
	output wire fib_42_s_axi_control_ARREADY;
	input fib_42_s_axi_control_ARVALID;
	input [4:0] fib_42_s_axi_control_ARADDR;
	input fib_42_s_axi_control_RREADY;
	output wire fib_42_s_axi_control_RVALID;
	output wire [31:0] fib_42_s_axi_control_RDATA;
	output wire [1:0] fib_42_s_axi_control_RRESP;
	output wire fib_42_s_axi_control_AWREADY;
	input fib_42_s_axi_control_AWVALID;
	input [4:0] fib_42_s_axi_control_AWADDR;
	output wire fib_42_s_axi_control_WREADY;
	input fib_42_s_axi_control_WVALID;
	input [31:0] fib_42_s_axi_control_WDATA;
	input [3:0] fib_42_s_axi_control_WSTRB;
	input fib_42_s_axi_control_BREADY;
	output wire fib_42_s_axi_control_BVALID;
	output wire [1:0] fib_42_s_axi_control_BRESP;
	input fib_43_m_axi_gmem_ARREADY;
	output wire fib_43_m_axi_gmem_ARVALID;
	output wire fib_43_m_axi_gmem_ARID;
	output wire [63:0] fib_43_m_axi_gmem_ARADDR;
	output wire [7:0] fib_43_m_axi_gmem_ARLEN;
	output wire [2:0] fib_43_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_43_m_axi_gmem_ARBURST;
	output wire fib_43_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_43_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_43_m_axi_gmem_ARPROT;
	output wire [3:0] fib_43_m_axi_gmem_ARQOS;
	output wire [3:0] fib_43_m_axi_gmem_ARREGION;
	output wire fib_43_m_axi_gmem_ARUSER;
	output wire fib_43_m_axi_gmem_RREADY;
	input fib_43_m_axi_gmem_RVALID;
	input fib_43_m_axi_gmem_RID;
	input [63:0] fib_43_m_axi_gmem_RDATA;
	input [1:0] fib_43_m_axi_gmem_RRESP;
	input fib_43_m_axi_gmem_RLAST;
	input fib_43_m_axi_gmem_RUSER;
	input fib_43_m_axi_gmem_AWREADY;
	output wire fib_43_m_axi_gmem_AWVALID;
	output wire fib_43_m_axi_gmem_AWID;
	output wire [63:0] fib_43_m_axi_gmem_AWADDR;
	output wire [7:0] fib_43_m_axi_gmem_AWLEN;
	output wire [2:0] fib_43_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_43_m_axi_gmem_AWBURST;
	output wire fib_43_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_43_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_43_m_axi_gmem_AWPROT;
	output wire [3:0] fib_43_m_axi_gmem_AWQOS;
	output wire [3:0] fib_43_m_axi_gmem_AWREGION;
	output wire fib_43_m_axi_gmem_AWUSER;
	input fib_43_m_axi_gmem_WREADY;
	output wire fib_43_m_axi_gmem_WVALID;
	output wire [63:0] fib_43_m_axi_gmem_WDATA;
	output wire [7:0] fib_43_m_axi_gmem_WSTRB;
	output wire fib_43_m_axi_gmem_WLAST;
	output wire fib_43_m_axi_gmem_WUSER;
	output wire fib_43_m_axi_gmem_BREADY;
	input fib_43_m_axi_gmem_BVALID;
	input fib_43_m_axi_gmem_BID;
	input [1:0] fib_43_m_axi_gmem_BRESP;
	input fib_43_m_axi_gmem_BUSER;
	output wire fib_43_s_axi_control_ARREADY;
	input fib_43_s_axi_control_ARVALID;
	input [4:0] fib_43_s_axi_control_ARADDR;
	input fib_43_s_axi_control_RREADY;
	output wire fib_43_s_axi_control_RVALID;
	output wire [31:0] fib_43_s_axi_control_RDATA;
	output wire [1:0] fib_43_s_axi_control_RRESP;
	output wire fib_43_s_axi_control_AWREADY;
	input fib_43_s_axi_control_AWVALID;
	input [4:0] fib_43_s_axi_control_AWADDR;
	output wire fib_43_s_axi_control_WREADY;
	input fib_43_s_axi_control_WVALID;
	input [31:0] fib_43_s_axi_control_WDATA;
	input [3:0] fib_43_s_axi_control_WSTRB;
	input fib_43_s_axi_control_BREADY;
	output wire fib_43_s_axi_control_BVALID;
	output wire [1:0] fib_43_s_axi_control_BRESP;
	input fib_44_m_axi_gmem_ARREADY;
	output wire fib_44_m_axi_gmem_ARVALID;
	output wire fib_44_m_axi_gmem_ARID;
	output wire [63:0] fib_44_m_axi_gmem_ARADDR;
	output wire [7:0] fib_44_m_axi_gmem_ARLEN;
	output wire [2:0] fib_44_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_44_m_axi_gmem_ARBURST;
	output wire fib_44_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_44_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_44_m_axi_gmem_ARPROT;
	output wire [3:0] fib_44_m_axi_gmem_ARQOS;
	output wire [3:0] fib_44_m_axi_gmem_ARREGION;
	output wire fib_44_m_axi_gmem_ARUSER;
	output wire fib_44_m_axi_gmem_RREADY;
	input fib_44_m_axi_gmem_RVALID;
	input fib_44_m_axi_gmem_RID;
	input [63:0] fib_44_m_axi_gmem_RDATA;
	input [1:0] fib_44_m_axi_gmem_RRESP;
	input fib_44_m_axi_gmem_RLAST;
	input fib_44_m_axi_gmem_RUSER;
	input fib_44_m_axi_gmem_AWREADY;
	output wire fib_44_m_axi_gmem_AWVALID;
	output wire fib_44_m_axi_gmem_AWID;
	output wire [63:0] fib_44_m_axi_gmem_AWADDR;
	output wire [7:0] fib_44_m_axi_gmem_AWLEN;
	output wire [2:0] fib_44_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_44_m_axi_gmem_AWBURST;
	output wire fib_44_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_44_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_44_m_axi_gmem_AWPROT;
	output wire [3:0] fib_44_m_axi_gmem_AWQOS;
	output wire [3:0] fib_44_m_axi_gmem_AWREGION;
	output wire fib_44_m_axi_gmem_AWUSER;
	input fib_44_m_axi_gmem_WREADY;
	output wire fib_44_m_axi_gmem_WVALID;
	output wire [63:0] fib_44_m_axi_gmem_WDATA;
	output wire [7:0] fib_44_m_axi_gmem_WSTRB;
	output wire fib_44_m_axi_gmem_WLAST;
	output wire fib_44_m_axi_gmem_WUSER;
	output wire fib_44_m_axi_gmem_BREADY;
	input fib_44_m_axi_gmem_BVALID;
	input fib_44_m_axi_gmem_BID;
	input [1:0] fib_44_m_axi_gmem_BRESP;
	input fib_44_m_axi_gmem_BUSER;
	output wire fib_44_s_axi_control_ARREADY;
	input fib_44_s_axi_control_ARVALID;
	input [4:0] fib_44_s_axi_control_ARADDR;
	input fib_44_s_axi_control_RREADY;
	output wire fib_44_s_axi_control_RVALID;
	output wire [31:0] fib_44_s_axi_control_RDATA;
	output wire [1:0] fib_44_s_axi_control_RRESP;
	output wire fib_44_s_axi_control_AWREADY;
	input fib_44_s_axi_control_AWVALID;
	input [4:0] fib_44_s_axi_control_AWADDR;
	output wire fib_44_s_axi_control_WREADY;
	input fib_44_s_axi_control_WVALID;
	input [31:0] fib_44_s_axi_control_WDATA;
	input [3:0] fib_44_s_axi_control_WSTRB;
	input fib_44_s_axi_control_BREADY;
	output wire fib_44_s_axi_control_BVALID;
	output wire [1:0] fib_44_s_axi_control_BRESP;
	input fib_45_m_axi_gmem_ARREADY;
	output wire fib_45_m_axi_gmem_ARVALID;
	output wire fib_45_m_axi_gmem_ARID;
	output wire [63:0] fib_45_m_axi_gmem_ARADDR;
	output wire [7:0] fib_45_m_axi_gmem_ARLEN;
	output wire [2:0] fib_45_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_45_m_axi_gmem_ARBURST;
	output wire fib_45_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_45_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_45_m_axi_gmem_ARPROT;
	output wire [3:0] fib_45_m_axi_gmem_ARQOS;
	output wire [3:0] fib_45_m_axi_gmem_ARREGION;
	output wire fib_45_m_axi_gmem_ARUSER;
	output wire fib_45_m_axi_gmem_RREADY;
	input fib_45_m_axi_gmem_RVALID;
	input fib_45_m_axi_gmem_RID;
	input [63:0] fib_45_m_axi_gmem_RDATA;
	input [1:0] fib_45_m_axi_gmem_RRESP;
	input fib_45_m_axi_gmem_RLAST;
	input fib_45_m_axi_gmem_RUSER;
	input fib_45_m_axi_gmem_AWREADY;
	output wire fib_45_m_axi_gmem_AWVALID;
	output wire fib_45_m_axi_gmem_AWID;
	output wire [63:0] fib_45_m_axi_gmem_AWADDR;
	output wire [7:0] fib_45_m_axi_gmem_AWLEN;
	output wire [2:0] fib_45_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_45_m_axi_gmem_AWBURST;
	output wire fib_45_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_45_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_45_m_axi_gmem_AWPROT;
	output wire [3:0] fib_45_m_axi_gmem_AWQOS;
	output wire [3:0] fib_45_m_axi_gmem_AWREGION;
	output wire fib_45_m_axi_gmem_AWUSER;
	input fib_45_m_axi_gmem_WREADY;
	output wire fib_45_m_axi_gmem_WVALID;
	output wire [63:0] fib_45_m_axi_gmem_WDATA;
	output wire [7:0] fib_45_m_axi_gmem_WSTRB;
	output wire fib_45_m_axi_gmem_WLAST;
	output wire fib_45_m_axi_gmem_WUSER;
	output wire fib_45_m_axi_gmem_BREADY;
	input fib_45_m_axi_gmem_BVALID;
	input fib_45_m_axi_gmem_BID;
	input [1:0] fib_45_m_axi_gmem_BRESP;
	input fib_45_m_axi_gmem_BUSER;
	output wire fib_45_s_axi_control_ARREADY;
	input fib_45_s_axi_control_ARVALID;
	input [4:0] fib_45_s_axi_control_ARADDR;
	input fib_45_s_axi_control_RREADY;
	output wire fib_45_s_axi_control_RVALID;
	output wire [31:0] fib_45_s_axi_control_RDATA;
	output wire [1:0] fib_45_s_axi_control_RRESP;
	output wire fib_45_s_axi_control_AWREADY;
	input fib_45_s_axi_control_AWVALID;
	input [4:0] fib_45_s_axi_control_AWADDR;
	output wire fib_45_s_axi_control_WREADY;
	input fib_45_s_axi_control_WVALID;
	input [31:0] fib_45_s_axi_control_WDATA;
	input [3:0] fib_45_s_axi_control_WSTRB;
	input fib_45_s_axi_control_BREADY;
	output wire fib_45_s_axi_control_BVALID;
	output wire [1:0] fib_45_s_axi_control_BRESP;
	input fib_46_m_axi_gmem_ARREADY;
	output wire fib_46_m_axi_gmem_ARVALID;
	output wire fib_46_m_axi_gmem_ARID;
	output wire [63:0] fib_46_m_axi_gmem_ARADDR;
	output wire [7:0] fib_46_m_axi_gmem_ARLEN;
	output wire [2:0] fib_46_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_46_m_axi_gmem_ARBURST;
	output wire fib_46_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_46_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_46_m_axi_gmem_ARPROT;
	output wire [3:0] fib_46_m_axi_gmem_ARQOS;
	output wire [3:0] fib_46_m_axi_gmem_ARREGION;
	output wire fib_46_m_axi_gmem_ARUSER;
	output wire fib_46_m_axi_gmem_RREADY;
	input fib_46_m_axi_gmem_RVALID;
	input fib_46_m_axi_gmem_RID;
	input [63:0] fib_46_m_axi_gmem_RDATA;
	input [1:0] fib_46_m_axi_gmem_RRESP;
	input fib_46_m_axi_gmem_RLAST;
	input fib_46_m_axi_gmem_RUSER;
	input fib_46_m_axi_gmem_AWREADY;
	output wire fib_46_m_axi_gmem_AWVALID;
	output wire fib_46_m_axi_gmem_AWID;
	output wire [63:0] fib_46_m_axi_gmem_AWADDR;
	output wire [7:0] fib_46_m_axi_gmem_AWLEN;
	output wire [2:0] fib_46_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_46_m_axi_gmem_AWBURST;
	output wire fib_46_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_46_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_46_m_axi_gmem_AWPROT;
	output wire [3:0] fib_46_m_axi_gmem_AWQOS;
	output wire [3:0] fib_46_m_axi_gmem_AWREGION;
	output wire fib_46_m_axi_gmem_AWUSER;
	input fib_46_m_axi_gmem_WREADY;
	output wire fib_46_m_axi_gmem_WVALID;
	output wire [63:0] fib_46_m_axi_gmem_WDATA;
	output wire [7:0] fib_46_m_axi_gmem_WSTRB;
	output wire fib_46_m_axi_gmem_WLAST;
	output wire fib_46_m_axi_gmem_WUSER;
	output wire fib_46_m_axi_gmem_BREADY;
	input fib_46_m_axi_gmem_BVALID;
	input fib_46_m_axi_gmem_BID;
	input [1:0] fib_46_m_axi_gmem_BRESP;
	input fib_46_m_axi_gmem_BUSER;
	output wire fib_46_s_axi_control_ARREADY;
	input fib_46_s_axi_control_ARVALID;
	input [4:0] fib_46_s_axi_control_ARADDR;
	input fib_46_s_axi_control_RREADY;
	output wire fib_46_s_axi_control_RVALID;
	output wire [31:0] fib_46_s_axi_control_RDATA;
	output wire [1:0] fib_46_s_axi_control_RRESP;
	output wire fib_46_s_axi_control_AWREADY;
	input fib_46_s_axi_control_AWVALID;
	input [4:0] fib_46_s_axi_control_AWADDR;
	output wire fib_46_s_axi_control_WREADY;
	input fib_46_s_axi_control_WVALID;
	input [31:0] fib_46_s_axi_control_WDATA;
	input [3:0] fib_46_s_axi_control_WSTRB;
	input fib_46_s_axi_control_BREADY;
	output wire fib_46_s_axi_control_BVALID;
	output wire [1:0] fib_46_s_axi_control_BRESP;
	input fib_47_m_axi_gmem_ARREADY;
	output wire fib_47_m_axi_gmem_ARVALID;
	output wire fib_47_m_axi_gmem_ARID;
	output wire [63:0] fib_47_m_axi_gmem_ARADDR;
	output wire [7:0] fib_47_m_axi_gmem_ARLEN;
	output wire [2:0] fib_47_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_47_m_axi_gmem_ARBURST;
	output wire fib_47_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_47_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_47_m_axi_gmem_ARPROT;
	output wire [3:0] fib_47_m_axi_gmem_ARQOS;
	output wire [3:0] fib_47_m_axi_gmem_ARREGION;
	output wire fib_47_m_axi_gmem_ARUSER;
	output wire fib_47_m_axi_gmem_RREADY;
	input fib_47_m_axi_gmem_RVALID;
	input fib_47_m_axi_gmem_RID;
	input [63:0] fib_47_m_axi_gmem_RDATA;
	input [1:0] fib_47_m_axi_gmem_RRESP;
	input fib_47_m_axi_gmem_RLAST;
	input fib_47_m_axi_gmem_RUSER;
	input fib_47_m_axi_gmem_AWREADY;
	output wire fib_47_m_axi_gmem_AWVALID;
	output wire fib_47_m_axi_gmem_AWID;
	output wire [63:0] fib_47_m_axi_gmem_AWADDR;
	output wire [7:0] fib_47_m_axi_gmem_AWLEN;
	output wire [2:0] fib_47_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_47_m_axi_gmem_AWBURST;
	output wire fib_47_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_47_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_47_m_axi_gmem_AWPROT;
	output wire [3:0] fib_47_m_axi_gmem_AWQOS;
	output wire [3:0] fib_47_m_axi_gmem_AWREGION;
	output wire fib_47_m_axi_gmem_AWUSER;
	input fib_47_m_axi_gmem_WREADY;
	output wire fib_47_m_axi_gmem_WVALID;
	output wire [63:0] fib_47_m_axi_gmem_WDATA;
	output wire [7:0] fib_47_m_axi_gmem_WSTRB;
	output wire fib_47_m_axi_gmem_WLAST;
	output wire fib_47_m_axi_gmem_WUSER;
	output wire fib_47_m_axi_gmem_BREADY;
	input fib_47_m_axi_gmem_BVALID;
	input fib_47_m_axi_gmem_BID;
	input [1:0] fib_47_m_axi_gmem_BRESP;
	input fib_47_m_axi_gmem_BUSER;
	output wire fib_47_s_axi_control_ARREADY;
	input fib_47_s_axi_control_ARVALID;
	input [4:0] fib_47_s_axi_control_ARADDR;
	input fib_47_s_axi_control_RREADY;
	output wire fib_47_s_axi_control_RVALID;
	output wire [31:0] fib_47_s_axi_control_RDATA;
	output wire [1:0] fib_47_s_axi_control_RRESP;
	output wire fib_47_s_axi_control_AWREADY;
	input fib_47_s_axi_control_AWVALID;
	input [4:0] fib_47_s_axi_control_AWADDR;
	output wire fib_47_s_axi_control_WREADY;
	input fib_47_s_axi_control_WVALID;
	input [31:0] fib_47_s_axi_control_WDATA;
	input [3:0] fib_47_s_axi_control_WSTRB;
	input fib_47_s_axi_control_BREADY;
	output wire fib_47_s_axi_control_BVALID;
	output wire [1:0] fib_47_s_axi_control_BRESP;
	input fib_48_m_axi_gmem_ARREADY;
	output wire fib_48_m_axi_gmem_ARVALID;
	output wire fib_48_m_axi_gmem_ARID;
	output wire [63:0] fib_48_m_axi_gmem_ARADDR;
	output wire [7:0] fib_48_m_axi_gmem_ARLEN;
	output wire [2:0] fib_48_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_48_m_axi_gmem_ARBURST;
	output wire fib_48_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_48_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_48_m_axi_gmem_ARPROT;
	output wire [3:0] fib_48_m_axi_gmem_ARQOS;
	output wire [3:0] fib_48_m_axi_gmem_ARREGION;
	output wire fib_48_m_axi_gmem_ARUSER;
	output wire fib_48_m_axi_gmem_RREADY;
	input fib_48_m_axi_gmem_RVALID;
	input fib_48_m_axi_gmem_RID;
	input [63:0] fib_48_m_axi_gmem_RDATA;
	input [1:0] fib_48_m_axi_gmem_RRESP;
	input fib_48_m_axi_gmem_RLAST;
	input fib_48_m_axi_gmem_RUSER;
	input fib_48_m_axi_gmem_AWREADY;
	output wire fib_48_m_axi_gmem_AWVALID;
	output wire fib_48_m_axi_gmem_AWID;
	output wire [63:0] fib_48_m_axi_gmem_AWADDR;
	output wire [7:0] fib_48_m_axi_gmem_AWLEN;
	output wire [2:0] fib_48_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_48_m_axi_gmem_AWBURST;
	output wire fib_48_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_48_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_48_m_axi_gmem_AWPROT;
	output wire [3:0] fib_48_m_axi_gmem_AWQOS;
	output wire [3:0] fib_48_m_axi_gmem_AWREGION;
	output wire fib_48_m_axi_gmem_AWUSER;
	input fib_48_m_axi_gmem_WREADY;
	output wire fib_48_m_axi_gmem_WVALID;
	output wire [63:0] fib_48_m_axi_gmem_WDATA;
	output wire [7:0] fib_48_m_axi_gmem_WSTRB;
	output wire fib_48_m_axi_gmem_WLAST;
	output wire fib_48_m_axi_gmem_WUSER;
	output wire fib_48_m_axi_gmem_BREADY;
	input fib_48_m_axi_gmem_BVALID;
	input fib_48_m_axi_gmem_BID;
	input [1:0] fib_48_m_axi_gmem_BRESP;
	input fib_48_m_axi_gmem_BUSER;
	output wire fib_48_s_axi_control_ARREADY;
	input fib_48_s_axi_control_ARVALID;
	input [4:0] fib_48_s_axi_control_ARADDR;
	input fib_48_s_axi_control_RREADY;
	output wire fib_48_s_axi_control_RVALID;
	output wire [31:0] fib_48_s_axi_control_RDATA;
	output wire [1:0] fib_48_s_axi_control_RRESP;
	output wire fib_48_s_axi_control_AWREADY;
	input fib_48_s_axi_control_AWVALID;
	input [4:0] fib_48_s_axi_control_AWADDR;
	output wire fib_48_s_axi_control_WREADY;
	input fib_48_s_axi_control_WVALID;
	input [31:0] fib_48_s_axi_control_WDATA;
	input [3:0] fib_48_s_axi_control_WSTRB;
	input fib_48_s_axi_control_BREADY;
	output wire fib_48_s_axi_control_BVALID;
	output wire [1:0] fib_48_s_axi_control_BRESP;
	input fib_49_m_axi_gmem_ARREADY;
	output wire fib_49_m_axi_gmem_ARVALID;
	output wire fib_49_m_axi_gmem_ARID;
	output wire [63:0] fib_49_m_axi_gmem_ARADDR;
	output wire [7:0] fib_49_m_axi_gmem_ARLEN;
	output wire [2:0] fib_49_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_49_m_axi_gmem_ARBURST;
	output wire fib_49_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_49_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_49_m_axi_gmem_ARPROT;
	output wire [3:0] fib_49_m_axi_gmem_ARQOS;
	output wire [3:0] fib_49_m_axi_gmem_ARREGION;
	output wire fib_49_m_axi_gmem_ARUSER;
	output wire fib_49_m_axi_gmem_RREADY;
	input fib_49_m_axi_gmem_RVALID;
	input fib_49_m_axi_gmem_RID;
	input [63:0] fib_49_m_axi_gmem_RDATA;
	input [1:0] fib_49_m_axi_gmem_RRESP;
	input fib_49_m_axi_gmem_RLAST;
	input fib_49_m_axi_gmem_RUSER;
	input fib_49_m_axi_gmem_AWREADY;
	output wire fib_49_m_axi_gmem_AWVALID;
	output wire fib_49_m_axi_gmem_AWID;
	output wire [63:0] fib_49_m_axi_gmem_AWADDR;
	output wire [7:0] fib_49_m_axi_gmem_AWLEN;
	output wire [2:0] fib_49_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_49_m_axi_gmem_AWBURST;
	output wire fib_49_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_49_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_49_m_axi_gmem_AWPROT;
	output wire [3:0] fib_49_m_axi_gmem_AWQOS;
	output wire [3:0] fib_49_m_axi_gmem_AWREGION;
	output wire fib_49_m_axi_gmem_AWUSER;
	input fib_49_m_axi_gmem_WREADY;
	output wire fib_49_m_axi_gmem_WVALID;
	output wire [63:0] fib_49_m_axi_gmem_WDATA;
	output wire [7:0] fib_49_m_axi_gmem_WSTRB;
	output wire fib_49_m_axi_gmem_WLAST;
	output wire fib_49_m_axi_gmem_WUSER;
	output wire fib_49_m_axi_gmem_BREADY;
	input fib_49_m_axi_gmem_BVALID;
	input fib_49_m_axi_gmem_BID;
	input [1:0] fib_49_m_axi_gmem_BRESP;
	input fib_49_m_axi_gmem_BUSER;
	output wire fib_49_s_axi_control_ARREADY;
	input fib_49_s_axi_control_ARVALID;
	input [4:0] fib_49_s_axi_control_ARADDR;
	input fib_49_s_axi_control_RREADY;
	output wire fib_49_s_axi_control_RVALID;
	output wire [31:0] fib_49_s_axi_control_RDATA;
	output wire [1:0] fib_49_s_axi_control_RRESP;
	output wire fib_49_s_axi_control_AWREADY;
	input fib_49_s_axi_control_AWVALID;
	input [4:0] fib_49_s_axi_control_AWADDR;
	output wire fib_49_s_axi_control_WREADY;
	input fib_49_s_axi_control_WVALID;
	input [31:0] fib_49_s_axi_control_WDATA;
	input [3:0] fib_49_s_axi_control_WSTRB;
	input fib_49_s_axi_control_BREADY;
	output wire fib_49_s_axi_control_BVALID;
	output wire [1:0] fib_49_s_axi_control_BRESP;
	input fib_50_m_axi_gmem_ARREADY;
	output wire fib_50_m_axi_gmem_ARVALID;
	output wire fib_50_m_axi_gmem_ARID;
	output wire [63:0] fib_50_m_axi_gmem_ARADDR;
	output wire [7:0] fib_50_m_axi_gmem_ARLEN;
	output wire [2:0] fib_50_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_50_m_axi_gmem_ARBURST;
	output wire fib_50_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_50_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_50_m_axi_gmem_ARPROT;
	output wire [3:0] fib_50_m_axi_gmem_ARQOS;
	output wire [3:0] fib_50_m_axi_gmem_ARREGION;
	output wire fib_50_m_axi_gmem_ARUSER;
	output wire fib_50_m_axi_gmem_RREADY;
	input fib_50_m_axi_gmem_RVALID;
	input fib_50_m_axi_gmem_RID;
	input [63:0] fib_50_m_axi_gmem_RDATA;
	input [1:0] fib_50_m_axi_gmem_RRESP;
	input fib_50_m_axi_gmem_RLAST;
	input fib_50_m_axi_gmem_RUSER;
	input fib_50_m_axi_gmem_AWREADY;
	output wire fib_50_m_axi_gmem_AWVALID;
	output wire fib_50_m_axi_gmem_AWID;
	output wire [63:0] fib_50_m_axi_gmem_AWADDR;
	output wire [7:0] fib_50_m_axi_gmem_AWLEN;
	output wire [2:0] fib_50_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_50_m_axi_gmem_AWBURST;
	output wire fib_50_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_50_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_50_m_axi_gmem_AWPROT;
	output wire [3:0] fib_50_m_axi_gmem_AWQOS;
	output wire [3:0] fib_50_m_axi_gmem_AWREGION;
	output wire fib_50_m_axi_gmem_AWUSER;
	input fib_50_m_axi_gmem_WREADY;
	output wire fib_50_m_axi_gmem_WVALID;
	output wire [63:0] fib_50_m_axi_gmem_WDATA;
	output wire [7:0] fib_50_m_axi_gmem_WSTRB;
	output wire fib_50_m_axi_gmem_WLAST;
	output wire fib_50_m_axi_gmem_WUSER;
	output wire fib_50_m_axi_gmem_BREADY;
	input fib_50_m_axi_gmem_BVALID;
	input fib_50_m_axi_gmem_BID;
	input [1:0] fib_50_m_axi_gmem_BRESP;
	input fib_50_m_axi_gmem_BUSER;
	output wire fib_50_s_axi_control_ARREADY;
	input fib_50_s_axi_control_ARVALID;
	input [4:0] fib_50_s_axi_control_ARADDR;
	input fib_50_s_axi_control_RREADY;
	output wire fib_50_s_axi_control_RVALID;
	output wire [31:0] fib_50_s_axi_control_RDATA;
	output wire [1:0] fib_50_s_axi_control_RRESP;
	output wire fib_50_s_axi_control_AWREADY;
	input fib_50_s_axi_control_AWVALID;
	input [4:0] fib_50_s_axi_control_AWADDR;
	output wire fib_50_s_axi_control_WREADY;
	input fib_50_s_axi_control_WVALID;
	input [31:0] fib_50_s_axi_control_WDATA;
	input [3:0] fib_50_s_axi_control_WSTRB;
	input fib_50_s_axi_control_BREADY;
	output wire fib_50_s_axi_control_BVALID;
	output wire [1:0] fib_50_s_axi_control_BRESP;
	input fib_51_m_axi_gmem_ARREADY;
	output wire fib_51_m_axi_gmem_ARVALID;
	output wire fib_51_m_axi_gmem_ARID;
	output wire [63:0] fib_51_m_axi_gmem_ARADDR;
	output wire [7:0] fib_51_m_axi_gmem_ARLEN;
	output wire [2:0] fib_51_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_51_m_axi_gmem_ARBURST;
	output wire fib_51_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_51_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_51_m_axi_gmem_ARPROT;
	output wire [3:0] fib_51_m_axi_gmem_ARQOS;
	output wire [3:0] fib_51_m_axi_gmem_ARREGION;
	output wire fib_51_m_axi_gmem_ARUSER;
	output wire fib_51_m_axi_gmem_RREADY;
	input fib_51_m_axi_gmem_RVALID;
	input fib_51_m_axi_gmem_RID;
	input [63:0] fib_51_m_axi_gmem_RDATA;
	input [1:0] fib_51_m_axi_gmem_RRESP;
	input fib_51_m_axi_gmem_RLAST;
	input fib_51_m_axi_gmem_RUSER;
	input fib_51_m_axi_gmem_AWREADY;
	output wire fib_51_m_axi_gmem_AWVALID;
	output wire fib_51_m_axi_gmem_AWID;
	output wire [63:0] fib_51_m_axi_gmem_AWADDR;
	output wire [7:0] fib_51_m_axi_gmem_AWLEN;
	output wire [2:0] fib_51_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_51_m_axi_gmem_AWBURST;
	output wire fib_51_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_51_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_51_m_axi_gmem_AWPROT;
	output wire [3:0] fib_51_m_axi_gmem_AWQOS;
	output wire [3:0] fib_51_m_axi_gmem_AWREGION;
	output wire fib_51_m_axi_gmem_AWUSER;
	input fib_51_m_axi_gmem_WREADY;
	output wire fib_51_m_axi_gmem_WVALID;
	output wire [63:0] fib_51_m_axi_gmem_WDATA;
	output wire [7:0] fib_51_m_axi_gmem_WSTRB;
	output wire fib_51_m_axi_gmem_WLAST;
	output wire fib_51_m_axi_gmem_WUSER;
	output wire fib_51_m_axi_gmem_BREADY;
	input fib_51_m_axi_gmem_BVALID;
	input fib_51_m_axi_gmem_BID;
	input [1:0] fib_51_m_axi_gmem_BRESP;
	input fib_51_m_axi_gmem_BUSER;
	output wire fib_51_s_axi_control_ARREADY;
	input fib_51_s_axi_control_ARVALID;
	input [4:0] fib_51_s_axi_control_ARADDR;
	input fib_51_s_axi_control_RREADY;
	output wire fib_51_s_axi_control_RVALID;
	output wire [31:0] fib_51_s_axi_control_RDATA;
	output wire [1:0] fib_51_s_axi_control_RRESP;
	output wire fib_51_s_axi_control_AWREADY;
	input fib_51_s_axi_control_AWVALID;
	input [4:0] fib_51_s_axi_control_AWADDR;
	output wire fib_51_s_axi_control_WREADY;
	input fib_51_s_axi_control_WVALID;
	input [31:0] fib_51_s_axi_control_WDATA;
	input [3:0] fib_51_s_axi_control_WSTRB;
	input fib_51_s_axi_control_BREADY;
	output wire fib_51_s_axi_control_BVALID;
	output wire [1:0] fib_51_s_axi_control_BRESP;
	input fib_52_m_axi_gmem_ARREADY;
	output wire fib_52_m_axi_gmem_ARVALID;
	output wire fib_52_m_axi_gmem_ARID;
	output wire [63:0] fib_52_m_axi_gmem_ARADDR;
	output wire [7:0] fib_52_m_axi_gmem_ARLEN;
	output wire [2:0] fib_52_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_52_m_axi_gmem_ARBURST;
	output wire fib_52_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_52_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_52_m_axi_gmem_ARPROT;
	output wire [3:0] fib_52_m_axi_gmem_ARQOS;
	output wire [3:0] fib_52_m_axi_gmem_ARREGION;
	output wire fib_52_m_axi_gmem_ARUSER;
	output wire fib_52_m_axi_gmem_RREADY;
	input fib_52_m_axi_gmem_RVALID;
	input fib_52_m_axi_gmem_RID;
	input [63:0] fib_52_m_axi_gmem_RDATA;
	input [1:0] fib_52_m_axi_gmem_RRESP;
	input fib_52_m_axi_gmem_RLAST;
	input fib_52_m_axi_gmem_RUSER;
	input fib_52_m_axi_gmem_AWREADY;
	output wire fib_52_m_axi_gmem_AWVALID;
	output wire fib_52_m_axi_gmem_AWID;
	output wire [63:0] fib_52_m_axi_gmem_AWADDR;
	output wire [7:0] fib_52_m_axi_gmem_AWLEN;
	output wire [2:0] fib_52_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_52_m_axi_gmem_AWBURST;
	output wire fib_52_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_52_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_52_m_axi_gmem_AWPROT;
	output wire [3:0] fib_52_m_axi_gmem_AWQOS;
	output wire [3:0] fib_52_m_axi_gmem_AWREGION;
	output wire fib_52_m_axi_gmem_AWUSER;
	input fib_52_m_axi_gmem_WREADY;
	output wire fib_52_m_axi_gmem_WVALID;
	output wire [63:0] fib_52_m_axi_gmem_WDATA;
	output wire [7:0] fib_52_m_axi_gmem_WSTRB;
	output wire fib_52_m_axi_gmem_WLAST;
	output wire fib_52_m_axi_gmem_WUSER;
	output wire fib_52_m_axi_gmem_BREADY;
	input fib_52_m_axi_gmem_BVALID;
	input fib_52_m_axi_gmem_BID;
	input [1:0] fib_52_m_axi_gmem_BRESP;
	input fib_52_m_axi_gmem_BUSER;
	output wire fib_52_s_axi_control_ARREADY;
	input fib_52_s_axi_control_ARVALID;
	input [4:0] fib_52_s_axi_control_ARADDR;
	input fib_52_s_axi_control_RREADY;
	output wire fib_52_s_axi_control_RVALID;
	output wire [31:0] fib_52_s_axi_control_RDATA;
	output wire [1:0] fib_52_s_axi_control_RRESP;
	output wire fib_52_s_axi_control_AWREADY;
	input fib_52_s_axi_control_AWVALID;
	input [4:0] fib_52_s_axi_control_AWADDR;
	output wire fib_52_s_axi_control_WREADY;
	input fib_52_s_axi_control_WVALID;
	input [31:0] fib_52_s_axi_control_WDATA;
	input [3:0] fib_52_s_axi_control_WSTRB;
	input fib_52_s_axi_control_BREADY;
	output wire fib_52_s_axi_control_BVALID;
	output wire [1:0] fib_52_s_axi_control_BRESP;
	input fib_53_m_axi_gmem_ARREADY;
	output wire fib_53_m_axi_gmem_ARVALID;
	output wire fib_53_m_axi_gmem_ARID;
	output wire [63:0] fib_53_m_axi_gmem_ARADDR;
	output wire [7:0] fib_53_m_axi_gmem_ARLEN;
	output wire [2:0] fib_53_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_53_m_axi_gmem_ARBURST;
	output wire fib_53_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_53_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_53_m_axi_gmem_ARPROT;
	output wire [3:0] fib_53_m_axi_gmem_ARQOS;
	output wire [3:0] fib_53_m_axi_gmem_ARREGION;
	output wire fib_53_m_axi_gmem_ARUSER;
	output wire fib_53_m_axi_gmem_RREADY;
	input fib_53_m_axi_gmem_RVALID;
	input fib_53_m_axi_gmem_RID;
	input [63:0] fib_53_m_axi_gmem_RDATA;
	input [1:0] fib_53_m_axi_gmem_RRESP;
	input fib_53_m_axi_gmem_RLAST;
	input fib_53_m_axi_gmem_RUSER;
	input fib_53_m_axi_gmem_AWREADY;
	output wire fib_53_m_axi_gmem_AWVALID;
	output wire fib_53_m_axi_gmem_AWID;
	output wire [63:0] fib_53_m_axi_gmem_AWADDR;
	output wire [7:0] fib_53_m_axi_gmem_AWLEN;
	output wire [2:0] fib_53_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_53_m_axi_gmem_AWBURST;
	output wire fib_53_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_53_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_53_m_axi_gmem_AWPROT;
	output wire [3:0] fib_53_m_axi_gmem_AWQOS;
	output wire [3:0] fib_53_m_axi_gmem_AWREGION;
	output wire fib_53_m_axi_gmem_AWUSER;
	input fib_53_m_axi_gmem_WREADY;
	output wire fib_53_m_axi_gmem_WVALID;
	output wire [63:0] fib_53_m_axi_gmem_WDATA;
	output wire [7:0] fib_53_m_axi_gmem_WSTRB;
	output wire fib_53_m_axi_gmem_WLAST;
	output wire fib_53_m_axi_gmem_WUSER;
	output wire fib_53_m_axi_gmem_BREADY;
	input fib_53_m_axi_gmem_BVALID;
	input fib_53_m_axi_gmem_BID;
	input [1:0] fib_53_m_axi_gmem_BRESP;
	input fib_53_m_axi_gmem_BUSER;
	output wire fib_53_s_axi_control_ARREADY;
	input fib_53_s_axi_control_ARVALID;
	input [4:0] fib_53_s_axi_control_ARADDR;
	input fib_53_s_axi_control_RREADY;
	output wire fib_53_s_axi_control_RVALID;
	output wire [31:0] fib_53_s_axi_control_RDATA;
	output wire [1:0] fib_53_s_axi_control_RRESP;
	output wire fib_53_s_axi_control_AWREADY;
	input fib_53_s_axi_control_AWVALID;
	input [4:0] fib_53_s_axi_control_AWADDR;
	output wire fib_53_s_axi_control_WREADY;
	input fib_53_s_axi_control_WVALID;
	input [31:0] fib_53_s_axi_control_WDATA;
	input [3:0] fib_53_s_axi_control_WSTRB;
	input fib_53_s_axi_control_BREADY;
	output wire fib_53_s_axi_control_BVALID;
	output wire [1:0] fib_53_s_axi_control_BRESP;
	input fib_54_m_axi_gmem_ARREADY;
	output wire fib_54_m_axi_gmem_ARVALID;
	output wire fib_54_m_axi_gmem_ARID;
	output wire [63:0] fib_54_m_axi_gmem_ARADDR;
	output wire [7:0] fib_54_m_axi_gmem_ARLEN;
	output wire [2:0] fib_54_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_54_m_axi_gmem_ARBURST;
	output wire fib_54_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_54_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_54_m_axi_gmem_ARPROT;
	output wire [3:0] fib_54_m_axi_gmem_ARQOS;
	output wire [3:0] fib_54_m_axi_gmem_ARREGION;
	output wire fib_54_m_axi_gmem_ARUSER;
	output wire fib_54_m_axi_gmem_RREADY;
	input fib_54_m_axi_gmem_RVALID;
	input fib_54_m_axi_gmem_RID;
	input [63:0] fib_54_m_axi_gmem_RDATA;
	input [1:0] fib_54_m_axi_gmem_RRESP;
	input fib_54_m_axi_gmem_RLAST;
	input fib_54_m_axi_gmem_RUSER;
	input fib_54_m_axi_gmem_AWREADY;
	output wire fib_54_m_axi_gmem_AWVALID;
	output wire fib_54_m_axi_gmem_AWID;
	output wire [63:0] fib_54_m_axi_gmem_AWADDR;
	output wire [7:0] fib_54_m_axi_gmem_AWLEN;
	output wire [2:0] fib_54_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_54_m_axi_gmem_AWBURST;
	output wire fib_54_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_54_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_54_m_axi_gmem_AWPROT;
	output wire [3:0] fib_54_m_axi_gmem_AWQOS;
	output wire [3:0] fib_54_m_axi_gmem_AWREGION;
	output wire fib_54_m_axi_gmem_AWUSER;
	input fib_54_m_axi_gmem_WREADY;
	output wire fib_54_m_axi_gmem_WVALID;
	output wire [63:0] fib_54_m_axi_gmem_WDATA;
	output wire [7:0] fib_54_m_axi_gmem_WSTRB;
	output wire fib_54_m_axi_gmem_WLAST;
	output wire fib_54_m_axi_gmem_WUSER;
	output wire fib_54_m_axi_gmem_BREADY;
	input fib_54_m_axi_gmem_BVALID;
	input fib_54_m_axi_gmem_BID;
	input [1:0] fib_54_m_axi_gmem_BRESP;
	input fib_54_m_axi_gmem_BUSER;
	output wire fib_54_s_axi_control_ARREADY;
	input fib_54_s_axi_control_ARVALID;
	input [4:0] fib_54_s_axi_control_ARADDR;
	input fib_54_s_axi_control_RREADY;
	output wire fib_54_s_axi_control_RVALID;
	output wire [31:0] fib_54_s_axi_control_RDATA;
	output wire [1:0] fib_54_s_axi_control_RRESP;
	output wire fib_54_s_axi_control_AWREADY;
	input fib_54_s_axi_control_AWVALID;
	input [4:0] fib_54_s_axi_control_AWADDR;
	output wire fib_54_s_axi_control_WREADY;
	input fib_54_s_axi_control_WVALID;
	input [31:0] fib_54_s_axi_control_WDATA;
	input [3:0] fib_54_s_axi_control_WSTRB;
	input fib_54_s_axi_control_BREADY;
	output wire fib_54_s_axi_control_BVALID;
	output wire [1:0] fib_54_s_axi_control_BRESP;
	input fib_55_m_axi_gmem_ARREADY;
	output wire fib_55_m_axi_gmem_ARVALID;
	output wire fib_55_m_axi_gmem_ARID;
	output wire [63:0] fib_55_m_axi_gmem_ARADDR;
	output wire [7:0] fib_55_m_axi_gmem_ARLEN;
	output wire [2:0] fib_55_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_55_m_axi_gmem_ARBURST;
	output wire fib_55_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_55_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_55_m_axi_gmem_ARPROT;
	output wire [3:0] fib_55_m_axi_gmem_ARQOS;
	output wire [3:0] fib_55_m_axi_gmem_ARREGION;
	output wire fib_55_m_axi_gmem_ARUSER;
	output wire fib_55_m_axi_gmem_RREADY;
	input fib_55_m_axi_gmem_RVALID;
	input fib_55_m_axi_gmem_RID;
	input [63:0] fib_55_m_axi_gmem_RDATA;
	input [1:0] fib_55_m_axi_gmem_RRESP;
	input fib_55_m_axi_gmem_RLAST;
	input fib_55_m_axi_gmem_RUSER;
	input fib_55_m_axi_gmem_AWREADY;
	output wire fib_55_m_axi_gmem_AWVALID;
	output wire fib_55_m_axi_gmem_AWID;
	output wire [63:0] fib_55_m_axi_gmem_AWADDR;
	output wire [7:0] fib_55_m_axi_gmem_AWLEN;
	output wire [2:0] fib_55_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_55_m_axi_gmem_AWBURST;
	output wire fib_55_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_55_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_55_m_axi_gmem_AWPROT;
	output wire [3:0] fib_55_m_axi_gmem_AWQOS;
	output wire [3:0] fib_55_m_axi_gmem_AWREGION;
	output wire fib_55_m_axi_gmem_AWUSER;
	input fib_55_m_axi_gmem_WREADY;
	output wire fib_55_m_axi_gmem_WVALID;
	output wire [63:0] fib_55_m_axi_gmem_WDATA;
	output wire [7:0] fib_55_m_axi_gmem_WSTRB;
	output wire fib_55_m_axi_gmem_WLAST;
	output wire fib_55_m_axi_gmem_WUSER;
	output wire fib_55_m_axi_gmem_BREADY;
	input fib_55_m_axi_gmem_BVALID;
	input fib_55_m_axi_gmem_BID;
	input [1:0] fib_55_m_axi_gmem_BRESP;
	input fib_55_m_axi_gmem_BUSER;
	output wire fib_55_s_axi_control_ARREADY;
	input fib_55_s_axi_control_ARVALID;
	input [4:0] fib_55_s_axi_control_ARADDR;
	input fib_55_s_axi_control_RREADY;
	output wire fib_55_s_axi_control_RVALID;
	output wire [31:0] fib_55_s_axi_control_RDATA;
	output wire [1:0] fib_55_s_axi_control_RRESP;
	output wire fib_55_s_axi_control_AWREADY;
	input fib_55_s_axi_control_AWVALID;
	input [4:0] fib_55_s_axi_control_AWADDR;
	output wire fib_55_s_axi_control_WREADY;
	input fib_55_s_axi_control_WVALID;
	input [31:0] fib_55_s_axi_control_WDATA;
	input [3:0] fib_55_s_axi_control_WSTRB;
	input fib_55_s_axi_control_BREADY;
	output wire fib_55_s_axi_control_BVALID;
	output wire [1:0] fib_55_s_axi_control_BRESP;
	input fib_56_m_axi_gmem_ARREADY;
	output wire fib_56_m_axi_gmem_ARVALID;
	output wire fib_56_m_axi_gmem_ARID;
	output wire [63:0] fib_56_m_axi_gmem_ARADDR;
	output wire [7:0] fib_56_m_axi_gmem_ARLEN;
	output wire [2:0] fib_56_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_56_m_axi_gmem_ARBURST;
	output wire fib_56_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_56_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_56_m_axi_gmem_ARPROT;
	output wire [3:0] fib_56_m_axi_gmem_ARQOS;
	output wire [3:0] fib_56_m_axi_gmem_ARREGION;
	output wire fib_56_m_axi_gmem_ARUSER;
	output wire fib_56_m_axi_gmem_RREADY;
	input fib_56_m_axi_gmem_RVALID;
	input fib_56_m_axi_gmem_RID;
	input [63:0] fib_56_m_axi_gmem_RDATA;
	input [1:0] fib_56_m_axi_gmem_RRESP;
	input fib_56_m_axi_gmem_RLAST;
	input fib_56_m_axi_gmem_RUSER;
	input fib_56_m_axi_gmem_AWREADY;
	output wire fib_56_m_axi_gmem_AWVALID;
	output wire fib_56_m_axi_gmem_AWID;
	output wire [63:0] fib_56_m_axi_gmem_AWADDR;
	output wire [7:0] fib_56_m_axi_gmem_AWLEN;
	output wire [2:0] fib_56_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_56_m_axi_gmem_AWBURST;
	output wire fib_56_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_56_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_56_m_axi_gmem_AWPROT;
	output wire [3:0] fib_56_m_axi_gmem_AWQOS;
	output wire [3:0] fib_56_m_axi_gmem_AWREGION;
	output wire fib_56_m_axi_gmem_AWUSER;
	input fib_56_m_axi_gmem_WREADY;
	output wire fib_56_m_axi_gmem_WVALID;
	output wire [63:0] fib_56_m_axi_gmem_WDATA;
	output wire [7:0] fib_56_m_axi_gmem_WSTRB;
	output wire fib_56_m_axi_gmem_WLAST;
	output wire fib_56_m_axi_gmem_WUSER;
	output wire fib_56_m_axi_gmem_BREADY;
	input fib_56_m_axi_gmem_BVALID;
	input fib_56_m_axi_gmem_BID;
	input [1:0] fib_56_m_axi_gmem_BRESP;
	input fib_56_m_axi_gmem_BUSER;
	output wire fib_56_s_axi_control_ARREADY;
	input fib_56_s_axi_control_ARVALID;
	input [4:0] fib_56_s_axi_control_ARADDR;
	input fib_56_s_axi_control_RREADY;
	output wire fib_56_s_axi_control_RVALID;
	output wire [31:0] fib_56_s_axi_control_RDATA;
	output wire [1:0] fib_56_s_axi_control_RRESP;
	output wire fib_56_s_axi_control_AWREADY;
	input fib_56_s_axi_control_AWVALID;
	input [4:0] fib_56_s_axi_control_AWADDR;
	output wire fib_56_s_axi_control_WREADY;
	input fib_56_s_axi_control_WVALID;
	input [31:0] fib_56_s_axi_control_WDATA;
	input [3:0] fib_56_s_axi_control_WSTRB;
	input fib_56_s_axi_control_BREADY;
	output wire fib_56_s_axi_control_BVALID;
	output wire [1:0] fib_56_s_axi_control_BRESP;
	input fib_57_m_axi_gmem_ARREADY;
	output wire fib_57_m_axi_gmem_ARVALID;
	output wire fib_57_m_axi_gmem_ARID;
	output wire [63:0] fib_57_m_axi_gmem_ARADDR;
	output wire [7:0] fib_57_m_axi_gmem_ARLEN;
	output wire [2:0] fib_57_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_57_m_axi_gmem_ARBURST;
	output wire fib_57_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_57_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_57_m_axi_gmem_ARPROT;
	output wire [3:0] fib_57_m_axi_gmem_ARQOS;
	output wire [3:0] fib_57_m_axi_gmem_ARREGION;
	output wire fib_57_m_axi_gmem_ARUSER;
	output wire fib_57_m_axi_gmem_RREADY;
	input fib_57_m_axi_gmem_RVALID;
	input fib_57_m_axi_gmem_RID;
	input [63:0] fib_57_m_axi_gmem_RDATA;
	input [1:0] fib_57_m_axi_gmem_RRESP;
	input fib_57_m_axi_gmem_RLAST;
	input fib_57_m_axi_gmem_RUSER;
	input fib_57_m_axi_gmem_AWREADY;
	output wire fib_57_m_axi_gmem_AWVALID;
	output wire fib_57_m_axi_gmem_AWID;
	output wire [63:0] fib_57_m_axi_gmem_AWADDR;
	output wire [7:0] fib_57_m_axi_gmem_AWLEN;
	output wire [2:0] fib_57_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_57_m_axi_gmem_AWBURST;
	output wire fib_57_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_57_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_57_m_axi_gmem_AWPROT;
	output wire [3:0] fib_57_m_axi_gmem_AWQOS;
	output wire [3:0] fib_57_m_axi_gmem_AWREGION;
	output wire fib_57_m_axi_gmem_AWUSER;
	input fib_57_m_axi_gmem_WREADY;
	output wire fib_57_m_axi_gmem_WVALID;
	output wire [63:0] fib_57_m_axi_gmem_WDATA;
	output wire [7:0] fib_57_m_axi_gmem_WSTRB;
	output wire fib_57_m_axi_gmem_WLAST;
	output wire fib_57_m_axi_gmem_WUSER;
	output wire fib_57_m_axi_gmem_BREADY;
	input fib_57_m_axi_gmem_BVALID;
	input fib_57_m_axi_gmem_BID;
	input [1:0] fib_57_m_axi_gmem_BRESP;
	input fib_57_m_axi_gmem_BUSER;
	output wire fib_57_s_axi_control_ARREADY;
	input fib_57_s_axi_control_ARVALID;
	input [4:0] fib_57_s_axi_control_ARADDR;
	input fib_57_s_axi_control_RREADY;
	output wire fib_57_s_axi_control_RVALID;
	output wire [31:0] fib_57_s_axi_control_RDATA;
	output wire [1:0] fib_57_s_axi_control_RRESP;
	output wire fib_57_s_axi_control_AWREADY;
	input fib_57_s_axi_control_AWVALID;
	input [4:0] fib_57_s_axi_control_AWADDR;
	output wire fib_57_s_axi_control_WREADY;
	input fib_57_s_axi_control_WVALID;
	input [31:0] fib_57_s_axi_control_WDATA;
	input [3:0] fib_57_s_axi_control_WSTRB;
	input fib_57_s_axi_control_BREADY;
	output wire fib_57_s_axi_control_BVALID;
	output wire [1:0] fib_57_s_axi_control_BRESP;
	input fib_58_m_axi_gmem_ARREADY;
	output wire fib_58_m_axi_gmem_ARVALID;
	output wire fib_58_m_axi_gmem_ARID;
	output wire [63:0] fib_58_m_axi_gmem_ARADDR;
	output wire [7:0] fib_58_m_axi_gmem_ARLEN;
	output wire [2:0] fib_58_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_58_m_axi_gmem_ARBURST;
	output wire fib_58_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_58_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_58_m_axi_gmem_ARPROT;
	output wire [3:0] fib_58_m_axi_gmem_ARQOS;
	output wire [3:0] fib_58_m_axi_gmem_ARREGION;
	output wire fib_58_m_axi_gmem_ARUSER;
	output wire fib_58_m_axi_gmem_RREADY;
	input fib_58_m_axi_gmem_RVALID;
	input fib_58_m_axi_gmem_RID;
	input [63:0] fib_58_m_axi_gmem_RDATA;
	input [1:0] fib_58_m_axi_gmem_RRESP;
	input fib_58_m_axi_gmem_RLAST;
	input fib_58_m_axi_gmem_RUSER;
	input fib_58_m_axi_gmem_AWREADY;
	output wire fib_58_m_axi_gmem_AWVALID;
	output wire fib_58_m_axi_gmem_AWID;
	output wire [63:0] fib_58_m_axi_gmem_AWADDR;
	output wire [7:0] fib_58_m_axi_gmem_AWLEN;
	output wire [2:0] fib_58_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_58_m_axi_gmem_AWBURST;
	output wire fib_58_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_58_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_58_m_axi_gmem_AWPROT;
	output wire [3:0] fib_58_m_axi_gmem_AWQOS;
	output wire [3:0] fib_58_m_axi_gmem_AWREGION;
	output wire fib_58_m_axi_gmem_AWUSER;
	input fib_58_m_axi_gmem_WREADY;
	output wire fib_58_m_axi_gmem_WVALID;
	output wire [63:0] fib_58_m_axi_gmem_WDATA;
	output wire [7:0] fib_58_m_axi_gmem_WSTRB;
	output wire fib_58_m_axi_gmem_WLAST;
	output wire fib_58_m_axi_gmem_WUSER;
	output wire fib_58_m_axi_gmem_BREADY;
	input fib_58_m_axi_gmem_BVALID;
	input fib_58_m_axi_gmem_BID;
	input [1:0] fib_58_m_axi_gmem_BRESP;
	input fib_58_m_axi_gmem_BUSER;
	output wire fib_58_s_axi_control_ARREADY;
	input fib_58_s_axi_control_ARVALID;
	input [4:0] fib_58_s_axi_control_ARADDR;
	input fib_58_s_axi_control_RREADY;
	output wire fib_58_s_axi_control_RVALID;
	output wire [31:0] fib_58_s_axi_control_RDATA;
	output wire [1:0] fib_58_s_axi_control_RRESP;
	output wire fib_58_s_axi_control_AWREADY;
	input fib_58_s_axi_control_AWVALID;
	input [4:0] fib_58_s_axi_control_AWADDR;
	output wire fib_58_s_axi_control_WREADY;
	input fib_58_s_axi_control_WVALID;
	input [31:0] fib_58_s_axi_control_WDATA;
	input [3:0] fib_58_s_axi_control_WSTRB;
	input fib_58_s_axi_control_BREADY;
	output wire fib_58_s_axi_control_BVALID;
	output wire [1:0] fib_58_s_axi_control_BRESP;
	input fib_59_m_axi_gmem_ARREADY;
	output wire fib_59_m_axi_gmem_ARVALID;
	output wire fib_59_m_axi_gmem_ARID;
	output wire [63:0] fib_59_m_axi_gmem_ARADDR;
	output wire [7:0] fib_59_m_axi_gmem_ARLEN;
	output wire [2:0] fib_59_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_59_m_axi_gmem_ARBURST;
	output wire fib_59_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_59_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_59_m_axi_gmem_ARPROT;
	output wire [3:0] fib_59_m_axi_gmem_ARQOS;
	output wire [3:0] fib_59_m_axi_gmem_ARREGION;
	output wire fib_59_m_axi_gmem_ARUSER;
	output wire fib_59_m_axi_gmem_RREADY;
	input fib_59_m_axi_gmem_RVALID;
	input fib_59_m_axi_gmem_RID;
	input [63:0] fib_59_m_axi_gmem_RDATA;
	input [1:0] fib_59_m_axi_gmem_RRESP;
	input fib_59_m_axi_gmem_RLAST;
	input fib_59_m_axi_gmem_RUSER;
	input fib_59_m_axi_gmem_AWREADY;
	output wire fib_59_m_axi_gmem_AWVALID;
	output wire fib_59_m_axi_gmem_AWID;
	output wire [63:0] fib_59_m_axi_gmem_AWADDR;
	output wire [7:0] fib_59_m_axi_gmem_AWLEN;
	output wire [2:0] fib_59_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_59_m_axi_gmem_AWBURST;
	output wire fib_59_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_59_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_59_m_axi_gmem_AWPROT;
	output wire [3:0] fib_59_m_axi_gmem_AWQOS;
	output wire [3:0] fib_59_m_axi_gmem_AWREGION;
	output wire fib_59_m_axi_gmem_AWUSER;
	input fib_59_m_axi_gmem_WREADY;
	output wire fib_59_m_axi_gmem_WVALID;
	output wire [63:0] fib_59_m_axi_gmem_WDATA;
	output wire [7:0] fib_59_m_axi_gmem_WSTRB;
	output wire fib_59_m_axi_gmem_WLAST;
	output wire fib_59_m_axi_gmem_WUSER;
	output wire fib_59_m_axi_gmem_BREADY;
	input fib_59_m_axi_gmem_BVALID;
	input fib_59_m_axi_gmem_BID;
	input [1:0] fib_59_m_axi_gmem_BRESP;
	input fib_59_m_axi_gmem_BUSER;
	output wire fib_59_s_axi_control_ARREADY;
	input fib_59_s_axi_control_ARVALID;
	input [4:0] fib_59_s_axi_control_ARADDR;
	input fib_59_s_axi_control_RREADY;
	output wire fib_59_s_axi_control_RVALID;
	output wire [31:0] fib_59_s_axi_control_RDATA;
	output wire [1:0] fib_59_s_axi_control_RRESP;
	output wire fib_59_s_axi_control_AWREADY;
	input fib_59_s_axi_control_AWVALID;
	input [4:0] fib_59_s_axi_control_AWADDR;
	output wire fib_59_s_axi_control_WREADY;
	input fib_59_s_axi_control_WVALID;
	input [31:0] fib_59_s_axi_control_WDATA;
	input [3:0] fib_59_s_axi_control_WSTRB;
	input fib_59_s_axi_control_BREADY;
	output wire fib_59_s_axi_control_BVALID;
	output wire [1:0] fib_59_s_axi_control_BRESP;
	input fib_60_m_axi_gmem_ARREADY;
	output wire fib_60_m_axi_gmem_ARVALID;
	output wire fib_60_m_axi_gmem_ARID;
	output wire [63:0] fib_60_m_axi_gmem_ARADDR;
	output wire [7:0] fib_60_m_axi_gmem_ARLEN;
	output wire [2:0] fib_60_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_60_m_axi_gmem_ARBURST;
	output wire fib_60_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_60_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_60_m_axi_gmem_ARPROT;
	output wire [3:0] fib_60_m_axi_gmem_ARQOS;
	output wire [3:0] fib_60_m_axi_gmem_ARREGION;
	output wire fib_60_m_axi_gmem_ARUSER;
	output wire fib_60_m_axi_gmem_RREADY;
	input fib_60_m_axi_gmem_RVALID;
	input fib_60_m_axi_gmem_RID;
	input [63:0] fib_60_m_axi_gmem_RDATA;
	input [1:0] fib_60_m_axi_gmem_RRESP;
	input fib_60_m_axi_gmem_RLAST;
	input fib_60_m_axi_gmem_RUSER;
	input fib_60_m_axi_gmem_AWREADY;
	output wire fib_60_m_axi_gmem_AWVALID;
	output wire fib_60_m_axi_gmem_AWID;
	output wire [63:0] fib_60_m_axi_gmem_AWADDR;
	output wire [7:0] fib_60_m_axi_gmem_AWLEN;
	output wire [2:0] fib_60_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_60_m_axi_gmem_AWBURST;
	output wire fib_60_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_60_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_60_m_axi_gmem_AWPROT;
	output wire [3:0] fib_60_m_axi_gmem_AWQOS;
	output wire [3:0] fib_60_m_axi_gmem_AWREGION;
	output wire fib_60_m_axi_gmem_AWUSER;
	input fib_60_m_axi_gmem_WREADY;
	output wire fib_60_m_axi_gmem_WVALID;
	output wire [63:0] fib_60_m_axi_gmem_WDATA;
	output wire [7:0] fib_60_m_axi_gmem_WSTRB;
	output wire fib_60_m_axi_gmem_WLAST;
	output wire fib_60_m_axi_gmem_WUSER;
	output wire fib_60_m_axi_gmem_BREADY;
	input fib_60_m_axi_gmem_BVALID;
	input fib_60_m_axi_gmem_BID;
	input [1:0] fib_60_m_axi_gmem_BRESP;
	input fib_60_m_axi_gmem_BUSER;
	output wire fib_60_s_axi_control_ARREADY;
	input fib_60_s_axi_control_ARVALID;
	input [4:0] fib_60_s_axi_control_ARADDR;
	input fib_60_s_axi_control_RREADY;
	output wire fib_60_s_axi_control_RVALID;
	output wire [31:0] fib_60_s_axi_control_RDATA;
	output wire [1:0] fib_60_s_axi_control_RRESP;
	output wire fib_60_s_axi_control_AWREADY;
	input fib_60_s_axi_control_AWVALID;
	input [4:0] fib_60_s_axi_control_AWADDR;
	output wire fib_60_s_axi_control_WREADY;
	input fib_60_s_axi_control_WVALID;
	input [31:0] fib_60_s_axi_control_WDATA;
	input [3:0] fib_60_s_axi_control_WSTRB;
	input fib_60_s_axi_control_BREADY;
	output wire fib_60_s_axi_control_BVALID;
	output wire [1:0] fib_60_s_axi_control_BRESP;
	input fib_61_m_axi_gmem_ARREADY;
	output wire fib_61_m_axi_gmem_ARVALID;
	output wire fib_61_m_axi_gmem_ARID;
	output wire [63:0] fib_61_m_axi_gmem_ARADDR;
	output wire [7:0] fib_61_m_axi_gmem_ARLEN;
	output wire [2:0] fib_61_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_61_m_axi_gmem_ARBURST;
	output wire fib_61_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_61_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_61_m_axi_gmem_ARPROT;
	output wire [3:0] fib_61_m_axi_gmem_ARQOS;
	output wire [3:0] fib_61_m_axi_gmem_ARREGION;
	output wire fib_61_m_axi_gmem_ARUSER;
	output wire fib_61_m_axi_gmem_RREADY;
	input fib_61_m_axi_gmem_RVALID;
	input fib_61_m_axi_gmem_RID;
	input [63:0] fib_61_m_axi_gmem_RDATA;
	input [1:0] fib_61_m_axi_gmem_RRESP;
	input fib_61_m_axi_gmem_RLAST;
	input fib_61_m_axi_gmem_RUSER;
	input fib_61_m_axi_gmem_AWREADY;
	output wire fib_61_m_axi_gmem_AWVALID;
	output wire fib_61_m_axi_gmem_AWID;
	output wire [63:0] fib_61_m_axi_gmem_AWADDR;
	output wire [7:0] fib_61_m_axi_gmem_AWLEN;
	output wire [2:0] fib_61_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_61_m_axi_gmem_AWBURST;
	output wire fib_61_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_61_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_61_m_axi_gmem_AWPROT;
	output wire [3:0] fib_61_m_axi_gmem_AWQOS;
	output wire [3:0] fib_61_m_axi_gmem_AWREGION;
	output wire fib_61_m_axi_gmem_AWUSER;
	input fib_61_m_axi_gmem_WREADY;
	output wire fib_61_m_axi_gmem_WVALID;
	output wire [63:0] fib_61_m_axi_gmem_WDATA;
	output wire [7:0] fib_61_m_axi_gmem_WSTRB;
	output wire fib_61_m_axi_gmem_WLAST;
	output wire fib_61_m_axi_gmem_WUSER;
	output wire fib_61_m_axi_gmem_BREADY;
	input fib_61_m_axi_gmem_BVALID;
	input fib_61_m_axi_gmem_BID;
	input [1:0] fib_61_m_axi_gmem_BRESP;
	input fib_61_m_axi_gmem_BUSER;
	output wire fib_61_s_axi_control_ARREADY;
	input fib_61_s_axi_control_ARVALID;
	input [4:0] fib_61_s_axi_control_ARADDR;
	input fib_61_s_axi_control_RREADY;
	output wire fib_61_s_axi_control_RVALID;
	output wire [31:0] fib_61_s_axi_control_RDATA;
	output wire [1:0] fib_61_s_axi_control_RRESP;
	output wire fib_61_s_axi_control_AWREADY;
	input fib_61_s_axi_control_AWVALID;
	input [4:0] fib_61_s_axi_control_AWADDR;
	output wire fib_61_s_axi_control_WREADY;
	input fib_61_s_axi_control_WVALID;
	input [31:0] fib_61_s_axi_control_WDATA;
	input [3:0] fib_61_s_axi_control_WSTRB;
	input fib_61_s_axi_control_BREADY;
	output wire fib_61_s_axi_control_BVALID;
	output wire [1:0] fib_61_s_axi_control_BRESP;
	input fib_62_m_axi_gmem_ARREADY;
	output wire fib_62_m_axi_gmem_ARVALID;
	output wire fib_62_m_axi_gmem_ARID;
	output wire [63:0] fib_62_m_axi_gmem_ARADDR;
	output wire [7:0] fib_62_m_axi_gmem_ARLEN;
	output wire [2:0] fib_62_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_62_m_axi_gmem_ARBURST;
	output wire fib_62_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_62_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_62_m_axi_gmem_ARPROT;
	output wire [3:0] fib_62_m_axi_gmem_ARQOS;
	output wire [3:0] fib_62_m_axi_gmem_ARREGION;
	output wire fib_62_m_axi_gmem_ARUSER;
	output wire fib_62_m_axi_gmem_RREADY;
	input fib_62_m_axi_gmem_RVALID;
	input fib_62_m_axi_gmem_RID;
	input [63:0] fib_62_m_axi_gmem_RDATA;
	input [1:0] fib_62_m_axi_gmem_RRESP;
	input fib_62_m_axi_gmem_RLAST;
	input fib_62_m_axi_gmem_RUSER;
	input fib_62_m_axi_gmem_AWREADY;
	output wire fib_62_m_axi_gmem_AWVALID;
	output wire fib_62_m_axi_gmem_AWID;
	output wire [63:0] fib_62_m_axi_gmem_AWADDR;
	output wire [7:0] fib_62_m_axi_gmem_AWLEN;
	output wire [2:0] fib_62_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_62_m_axi_gmem_AWBURST;
	output wire fib_62_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_62_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_62_m_axi_gmem_AWPROT;
	output wire [3:0] fib_62_m_axi_gmem_AWQOS;
	output wire [3:0] fib_62_m_axi_gmem_AWREGION;
	output wire fib_62_m_axi_gmem_AWUSER;
	input fib_62_m_axi_gmem_WREADY;
	output wire fib_62_m_axi_gmem_WVALID;
	output wire [63:0] fib_62_m_axi_gmem_WDATA;
	output wire [7:0] fib_62_m_axi_gmem_WSTRB;
	output wire fib_62_m_axi_gmem_WLAST;
	output wire fib_62_m_axi_gmem_WUSER;
	output wire fib_62_m_axi_gmem_BREADY;
	input fib_62_m_axi_gmem_BVALID;
	input fib_62_m_axi_gmem_BID;
	input [1:0] fib_62_m_axi_gmem_BRESP;
	input fib_62_m_axi_gmem_BUSER;
	output wire fib_62_s_axi_control_ARREADY;
	input fib_62_s_axi_control_ARVALID;
	input [4:0] fib_62_s_axi_control_ARADDR;
	input fib_62_s_axi_control_RREADY;
	output wire fib_62_s_axi_control_RVALID;
	output wire [31:0] fib_62_s_axi_control_RDATA;
	output wire [1:0] fib_62_s_axi_control_RRESP;
	output wire fib_62_s_axi_control_AWREADY;
	input fib_62_s_axi_control_AWVALID;
	input [4:0] fib_62_s_axi_control_AWADDR;
	output wire fib_62_s_axi_control_WREADY;
	input fib_62_s_axi_control_WVALID;
	input [31:0] fib_62_s_axi_control_WDATA;
	input [3:0] fib_62_s_axi_control_WSTRB;
	input fib_62_s_axi_control_BREADY;
	output wire fib_62_s_axi_control_BVALID;
	output wire [1:0] fib_62_s_axi_control_BRESP;
	input fib_63_m_axi_gmem_ARREADY;
	output wire fib_63_m_axi_gmem_ARVALID;
	output wire fib_63_m_axi_gmem_ARID;
	output wire [63:0] fib_63_m_axi_gmem_ARADDR;
	output wire [7:0] fib_63_m_axi_gmem_ARLEN;
	output wire [2:0] fib_63_m_axi_gmem_ARSIZE;
	output wire [1:0] fib_63_m_axi_gmem_ARBURST;
	output wire fib_63_m_axi_gmem_ARLOCK;
	output wire [3:0] fib_63_m_axi_gmem_ARCACHE;
	output wire [2:0] fib_63_m_axi_gmem_ARPROT;
	output wire [3:0] fib_63_m_axi_gmem_ARQOS;
	output wire [3:0] fib_63_m_axi_gmem_ARREGION;
	output wire fib_63_m_axi_gmem_ARUSER;
	output wire fib_63_m_axi_gmem_RREADY;
	input fib_63_m_axi_gmem_RVALID;
	input fib_63_m_axi_gmem_RID;
	input [63:0] fib_63_m_axi_gmem_RDATA;
	input [1:0] fib_63_m_axi_gmem_RRESP;
	input fib_63_m_axi_gmem_RLAST;
	input fib_63_m_axi_gmem_RUSER;
	input fib_63_m_axi_gmem_AWREADY;
	output wire fib_63_m_axi_gmem_AWVALID;
	output wire fib_63_m_axi_gmem_AWID;
	output wire [63:0] fib_63_m_axi_gmem_AWADDR;
	output wire [7:0] fib_63_m_axi_gmem_AWLEN;
	output wire [2:0] fib_63_m_axi_gmem_AWSIZE;
	output wire [1:0] fib_63_m_axi_gmem_AWBURST;
	output wire fib_63_m_axi_gmem_AWLOCK;
	output wire [3:0] fib_63_m_axi_gmem_AWCACHE;
	output wire [2:0] fib_63_m_axi_gmem_AWPROT;
	output wire [3:0] fib_63_m_axi_gmem_AWQOS;
	output wire [3:0] fib_63_m_axi_gmem_AWREGION;
	output wire fib_63_m_axi_gmem_AWUSER;
	input fib_63_m_axi_gmem_WREADY;
	output wire fib_63_m_axi_gmem_WVALID;
	output wire [63:0] fib_63_m_axi_gmem_WDATA;
	output wire [7:0] fib_63_m_axi_gmem_WSTRB;
	output wire fib_63_m_axi_gmem_WLAST;
	output wire fib_63_m_axi_gmem_WUSER;
	output wire fib_63_m_axi_gmem_BREADY;
	input fib_63_m_axi_gmem_BVALID;
	input fib_63_m_axi_gmem_BID;
	input [1:0] fib_63_m_axi_gmem_BRESP;
	input fib_63_m_axi_gmem_BUSER;
	output wire fib_63_s_axi_control_ARREADY;
	input fib_63_s_axi_control_ARVALID;
	input [4:0] fib_63_s_axi_control_ARADDR;
	input fib_63_s_axi_control_RREADY;
	output wire fib_63_s_axi_control_RVALID;
	output wire [31:0] fib_63_s_axi_control_RDATA;
	output wire [1:0] fib_63_s_axi_control_RRESP;
	output wire fib_63_s_axi_control_AWREADY;
	input fib_63_s_axi_control_AWVALID;
	input [4:0] fib_63_s_axi_control_AWADDR;
	output wire fib_63_s_axi_control_WREADY;
	input fib_63_s_axi_control_WVALID;
	input [31:0] fib_63_s_axi_control_WDATA;
	input [3:0] fib_63_s_axi_control_WSTRB;
	input fib_63_s_axi_control_BREADY;
	output wire fib_63_s_axi_control_BVALID;
	output wire [1:0] fib_63_s_axi_control_BRESP;
	input fib_schedulerAXI_0_ARREADY;
	output wire fib_schedulerAXI_0_ARVALID;
	output wire [1:0] fib_schedulerAXI_0_ARID;
	output wire [63:0] fib_schedulerAXI_0_ARADDR;
	output wire [7:0] fib_schedulerAXI_0_ARLEN;
	output wire [2:0] fib_schedulerAXI_0_ARSIZE;
	output wire [1:0] fib_schedulerAXI_0_ARBURST;
	output wire fib_schedulerAXI_0_ARLOCK;
	output wire [3:0] fib_schedulerAXI_0_ARCACHE;
	output wire [2:0] fib_schedulerAXI_0_ARPROT;
	output wire [3:0] fib_schedulerAXI_0_ARQOS;
	output wire [3:0] fib_schedulerAXI_0_ARREGION;
	output wire fib_schedulerAXI_0_RREADY;
	input fib_schedulerAXI_0_RVALID;
	input [1:0] fib_schedulerAXI_0_RID;
	input [127:0] fib_schedulerAXI_0_RDATA;
	input [1:0] fib_schedulerAXI_0_RRESP;
	input fib_schedulerAXI_0_RLAST;
	input fib_schedulerAXI_0_AWREADY;
	output wire fib_schedulerAXI_0_AWVALID;
	output wire [1:0] fib_schedulerAXI_0_AWID;
	output wire [63:0] fib_schedulerAXI_0_AWADDR;
	output wire [7:0] fib_schedulerAXI_0_AWLEN;
	output wire [2:0] fib_schedulerAXI_0_AWSIZE;
	output wire [1:0] fib_schedulerAXI_0_AWBURST;
	output wire fib_schedulerAXI_0_AWLOCK;
	output wire [3:0] fib_schedulerAXI_0_AWCACHE;
	output wire [2:0] fib_schedulerAXI_0_AWPROT;
	output wire [3:0] fib_schedulerAXI_0_AWQOS;
	output wire [3:0] fib_schedulerAXI_0_AWREGION;
	input fib_schedulerAXI_0_WREADY;
	output wire fib_schedulerAXI_0_WVALID;
	output wire [127:0] fib_schedulerAXI_0_WDATA;
	output wire [15:0] fib_schedulerAXI_0_WSTRB;
	output wire fib_schedulerAXI_0_WLAST;
	output wire fib_schedulerAXI_0_BREADY;
	input fib_schedulerAXI_0_BVALID;
	input [1:0] fib_schedulerAXI_0_BID;
	input [1:0] fib_schedulerAXI_0_BRESP;
	input sum_0_m_axi_gmem_ARREADY;
	output wire sum_0_m_axi_gmem_ARVALID;
	output wire sum_0_m_axi_gmem_ARID;
	output wire [63:0] sum_0_m_axi_gmem_ARADDR;
	output wire [7:0] sum_0_m_axi_gmem_ARLEN;
	output wire [2:0] sum_0_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_0_m_axi_gmem_ARBURST;
	output wire sum_0_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_0_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_0_m_axi_gmem_ARPROT;
	output wire [3:0] sum_0_m_axi_gmem_ARQOS;
	output wire [3:0] sum_0_m_axi_gmem_ARREGION;
	output wire sum_0_m_axi_gmem_ARUSER;
	output wire sum_0_m_axi_gmem_RREADY;
	input sum_0_m_axi_gmem_RVALID;
	input sum_0_m_axi_gmem_RID;
	input [31:0] sum_0_m_axi_gmem_RDATA;
	input [1:0] sum_0_m_axi_gmem_RRESP;
	input sum_0_m_axi_gmem_RLAST;
	input sum_0_m_axi_gmem_RUSER;
	input sum_0_m_axi_gmem_AWREADY;
	output wire sum_0_m_axi_gmem_AWVALID;
	output wire sum_0_m_axi_gmem_AWID;
	output wire [63:0] sum_0_m_axi_gmem_AWADDR;
	output wire [7:0] sum_0_m_axi_gmem_AWLEN;
	output wire [2:0] sum_0_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_0_m_axi_gmem_AWBURST;
	output wire sum_0_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_0_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_0_m_axi_gmem_AWPROT;
	output wire [3:0] sum_0_m_axi_gmem_AWQOS;
	output wire [3:0] sum_0_m_axi_gmem_AWREGION;
	output wire sum_0_m_axi_gmem_AWUSER;
	input sum_0_m_axi_gmem_WREADY;
	output wire sum_0_m_axi_gmem_WVALID;
	output wire [31:0] sum_0_m_axi_gmem_WDATA;
	output wire [3:0] sum_0_m_axi_gmem_WSTRB;
	output wire sum_0_m_axi_gmem_WLAST;
	output wire sum_0_m_axi_gmem_WUSER;
	output wire sum_0_m_axi_gmem_BREADY;
	input sum_0_m_axi_gmem_BVALID;
	input sum_0_m_axi_gmem_BID;
	input [1:0] sum_0_m_axi_gmem_BRESP;
	input sum_0_m_axi_gmem_BUSER;
	output wire sum_0_s_axi_control_ARREADY;
	input sum_0_s_axi_control_ARVALID;
	input [4:0] sum_0_s_axi_control_ARADDR;
	input sum_0_s_axi_control_RREADY;
	output wire sum_0_s_axi_control_RVALID;
	output wire [31:0] sum_0_s_axi_control_RDATA;
	output wire [1:0] sum_0_s_axi_control_RRESP;
	output wire sum_0_s_axi_control_AWREADY;
	input sum_0_s_axi_control_AWVALID;
	input [4:0] sum_0_s_axi_control_AWADDR;
	output wire sum_0_s_axi_control_WREADY;
	input sum_0_s_axi_control_WVALID;
	input [31:0] sum_0_s_axi_control_WDATA;
	input [3:0] sum_0_s_axi_control_WSTRB;
	input sum_0_s_axi_control_BREADY;
	output wire sum_0_s_axi_control_BVALID;
	output wire [1:0] sum_0_s_axi_control_BRESP;
	input sum_1_m_axi_gmem_ARREADY;
	output wire sum_1_m_axi_gmem_ARVALID;
	output wire sum_1_m_axi_gmem_ARID;
	output wire [63:0] sum_1_m_axi_gmem_ARADDR;
	output wire [7:0] sum_1_m_axi_gmem_ARLEN;
	output wire [2:0] sum_1_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_1_m_axi_gmem_ARBURST;
	output wire sum_1_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_1_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_1_m_axi_gmem_ARPROT;
	output wire [3:0] sum_1_m_axi_gmem_ARQOS;
	output wire [3:0] sum_1_m_axi_gmem_ARREGION;
	output wire sum_1_m_axi_gmem_ARUSER;
	output wire sum_1_m_axi_gmem_RREADY;
	input sum_1_m_axi_gmem_RVALID;
	input sum_1_m_axi_gmem_RID;
	input [31:0] sum_1_m_axi_gmem_RDATA;
	input [1:0] sum_1_m_axi_gmem_RRESP;
	input sum_1_m_axi_gmem_RLAST;
	input sum_1_m_axi_gmem_RUSER;
	input sum_1_m_axi_gmem_AWREADY;
	output wire sum_1_m_axi_gmem_AWVALID;
	output wire sum_1_m_axi_gmem_AWID;
	output wire [63:0] sum_1_m_axi_gmem_AWADDR;
	output wire [7:0] sum_1_m_axi_gmem_AWLEN;
	output wire [2:0] sum_1_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_1_m_axi_gmem_AWBURST;
	output wire sum_1_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_1_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_1_m_axi_gmem_AWPROT;
	output wire [3:0] sum_1_m_axi_gmem_AWQOS;
	output wire [3:0] sum_1_m_axi_gmem_AWREGION;
	output wire sum_1_m_axi_gmem_AWUSER;
	input sum_1_m_axi_gmem_WREADY;
	output wire sum_1_m_axi_gmem_WVALID;
	output wire [31:0] sum_1_m_axi_gmem_WDATA;
	output wire [3:0] sum_1_m_axi_gmem_WSTRB;
	output wire sum_1_m_axi_gmem_WLAST;
	output wire sum_1_m_axi_gmem_WUSER;
	output wire sum_1_m_axi_gmem_BREADY;
	input sum_1_m_axi_gmem_BVALID;
	input sum_1_m_axi_gmem_BID;
	input [1:0] sum_1_m_axi_gmem_BRESP;
	input sum_1_m_axi_gmem_BUSER;
	output wire sum_1_s_axi_control_ARREADY;
	input sum_1_s_axi_control_ARVALID;
	input [4:0] sum_1_s_axi_control_ARADDR;
	input sum_1_s_axi_control_RREADY;
	output wire sum_1_s_axi_control_RVALID;
	output wire [31:0] sum_1_s_axi_control_RDATA;
	output wire [1:0] sum_1_s_axi_control_RRESP;
	output wire sum_1_s_axi_control_AWREADY;
	input sum_1_s_axi_control_AWVALID;
	input [4:0] sum_1_s_axi_control_AWADDR;
	output wire sum_1_s_axi_control_WREADY;
	input sum_1_s_axi_control_WVALID;
	input [31:0] sum_1_s_axi_control_WDATA;
	input [3:0] sum_1_s_axi_control_WSTRB;
	input sum_1_s_axi_control_BREADY;
	output wire sum_1_s_axi_control_BVALID;
	output wire [1:0] sum_1_s_axi_control_BRESP;
	input sum_2_m_axi_gmem_ARREADY;
	output wire sum_2_m_axi_gmem_ARVALID;
	output wire sum_2_m_axi_gmem_ARID;
	output wire [63:0] sum_2_m_axi_gmem_ARADDR;
	output wire [7:0] sum_2_m_axi_gmem_ARLEN;
	output wire [2:0] sum_2_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_2_m_axi_gmem_ARBURST;
	output wire sum_2_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_2_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_2_m_axi_gmem_ARPROT;
	output wire [3:0] sum_2_m_axi_gmem_ARQOS;
	output wire [3:0] sum_2_m_axi_gmem_ARREGION;
	output wire sum_2_m_axi_gmem_ARUSER;
	output wire sum_2_m_axi_gmem_RREADY;
	input sum_2_m_axi_gmem_RVALID;
	input sum_2_m_axi_gmem_RID;
	input [31:0] sum_2_m_axi_gmem_RDATA;
	input [1:0] sum_2_m_axi_gmem_RRESP;
	input sum_2_m_axi_gmem_RLAST;
	input sum_2_m_axi_gmem_RUSER;
	input sum_2_m_axi_gmem_AWREADY;
	output wire sum_2_m_axi_gmem_AWVALID;
	output wire sum_2_m_axi_gmem_AWID;
	output wire [63:0] sum_2_m_axi_gmem_AWADDR;
	output wire [7:0] sum_2_m_axi_gmem_AWLEN;
	output wire [2:0] sum_2_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_2_m_axi_gmem_AWBURST;
	output wire sum_2_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_2_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_2_m_axi_gmem_AWPROT;
	output wire [3:0] sum_2_m_axi_gmem_AWQOS;
	output wire [3:0] sum_2_m_axi_gmem_AWREGION;
	output wire sum_2_m_axi_gmem_AWUSER;
	input sum_2_m_axi_gmem_WREADY;
	output wire sum_2_m_axi_gmem_WVALID;
	output wire [31:0] sum_2_m_axi_gmem_WDATA;
	output wire [3:0] sum_2_m_axi_gmem_WSTRB;
	output wire sum_2_m_axi_gmem_WLAST;
	output wire sum_2_m_axi_gmem_WUSER;
	output wire sum_2_m_axi_gmem_BREADY;
	input sum_2_m_axi_gmem_BVALID;
	input sum_2_m_axi_gmem_BID;
	input [1:0] sum_2_m_axi_gmem_BRESP;
	input sum_2_m_axi_gmem_BUSER;
	output wire sum_2_s_axi_control_ARREADY;
	input sum_2_s_axi_control_ARVALID;
	input [4:0] sum_2_s_axi_control_ARADDR;
	input sum_2_s_axi_control_RREADY;
	output wire sum_2_s_axi_control_RVALID;
	output wire [31:0] sum_2_s_axi_control_RDATA;
	output wire [1:0] sum_2_s_axi_control_RRESP;
	output wire sum_2_s_axi_control_AWREADY;
	input sum_2_s_axi_control_AWVALID;
	input [4:0] sum_2_s_axi_control_AWADDR;
	output wire sum_2_s_axi_control_WREADY;
	input sum_2_s_axi_control_WVALID;
	input [31:0] sum_2_s_axi_control_WDATA;
	input [3:0] sum_2_s_axi_control_WSTRB;
	input sum_2_s_axi_control_BREADY;
	output wire sum_2_s_axi_control_BVALID;
	output wire [1:0] sum_2_s_axi_control_BRESP;
	input sum_3_m_axi_gmem_ARREADY;
	output wire sum_3_m_axi_gmem_ARVALID;
	output wire sum_3_m_axi_gmem_ARID;
	output wire [63:0] sum_3_m_axi_gmem_ARADDR;
	output wire [7:0] sum_3_m_axi_gmem_ARLEN;
	output wire [2:0] sum_3_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_3_m_axi_gmem_ARBURST;
	output wire sum_3_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_3_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_3_m_axi_gmem_ARPROT;
	output wire [3:0] sum_3_m_axi_gmem_ARQOS;
	output wire [3:0] sum_3_m_axi_gmem_ARREGION;
	output wire sum_3_m_axi_gmem_ARUSER;
	output wire sum_3_m_axi_gmem_RREADY;
	input sum_3_m_axi_gmem_RVALID;
	input sum_3_m_axi_gmem_RID;
	input [31:0] sum_3_m_axi_gmem_RDATA;
	input [1:0] sum_3_m_axi_gmem_RRESP;
	input sum_3_m_axi_gmem_RLAST;
	input sum_3_m_axi_gmem_RUSER;
	input sum_3_m_axi_gmem_AWREADY;
	output wire sum_3_m_axi_gmem_AWVALID;
	output wire sum_3_m_axi_gmem_AWID;
	output wire [63:0] sum_3_m_axi_gmem_AWADDR;
	output wire [7:0] sum_3_m_axi_gmem_AWLEN;
	output wire [2:0] sum_3_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_3_m_axi_gmem_AWBURST;
	output wire sum_3_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_3_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_3_m_axi_gmem_AWPROT;
	output wire [3:0] sum_3_m_axi_gmem_AWQOS;
	output wire [3:0] sum_3_m_axi_gmem_AWREGION;
	output wire sum_3_m_axi_gmem_AWUSER;
	input sum_3_m_axi_gmem_WREADY;
	output wire sum_3_m_axi_gmem_WVALID;
	output wire [31:0] sum_3_m_axi_gmem_WDATA;
	output wire [3:0] sum_3_m_axi_gmem_WSTRB;
	output wire sum_3_m_axi_gmem_WLAST;
	output wire sum_3_m_axi_gmem_WUSER;
	output wire sum_3_m_axi_gmem_BREADY;
	input sum_3_m_axi_gmem_BVALID;
	input sum_3_m_axi_gmem_BID;
	input [1:0] sum_3_m_axi_gmem_BRESP;
	input sum_3_m_axi_gmem_BUSER;
	output wire sum_3_s_axi_control_ARREADY;
	input sum_3_s_axi_control_ARVALID;
	input [4:0] sum_3_s_axi_control_ARADDR;
	input sum_3_s_axi_control_RREADY;
	output wire sum_3_s_axi_control_RVALID;
	output wire [31:0] sum_3_s_axi_control_RDATA;
	output wire [1:0] sum_3_s_axi_control_RRESP;
	output wire sum_3_s_axi_control_AWREADY;
	input sum_3_s_axi_control_AWVALID;
	input [4:0] sum_3_s_axi_control_AWADDR;
	output wire sum_3_s_axi_control_WREADY;
	input sum_3_s_axi_control_WVALID;
	input [31:0] sum_3_s_axi_control_WDATA;
	input [3:0] sum_3_s_axi_control_WSTRB;
	input sum_3_s_axi_control_BREADY;
	output wire sum_3_s_axi_control_BVALID;
	output wire [1:0] sum_3_s_axi_control_BRESP;
	input sum_4_m_axi_gmem_ARREADY;
	output wire sum_4_m_axi_gmem_ARVALID;
	output wire sum_4_m_axi_gmem_ARID;
	output wire [63:0] sum_4_m_axi_gmem_ARADDR;
	output wire [7:0] sum_4_m_axi_gmem_ARLEN;
	output wire [2:0] sum_4_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_4_m_axi_gmem_ARBURST;
	output wire sum_4_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_4_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_4_m_axi_gmem_ARPROT;
	output wire [3:0] sum_4_m_axi_gmem_ARQOS;
	output wire [3:0] sum_4_m_axi_gmem_ARREGION;
	output wire sum_4_m_axi_gmem_ARUSER;
	output wire sum_4_m_axi_gmem_RREADY;
	input sum_4_m_axi_gmem_RVALID;
	input sum_4_m_axi_gmem_RID;
	input [31:0] sum_4_m_axi_gmem_RDATA;
	input [1:0] sum_4_m_axi_gmem_RRESP;
	input sum_4_m_axi_gmem_RLAST;
	input sum_4_m_axi_gmem_RUSER;
	input sum_4_m_axi_gmem_AWREADY;
	output wire sum_4_m_axi_gmem_AWVALID;
	output wire sum_4_m_axi_gmem_AWID;
	output wire [63:0] sum_4_m_axi_gmem_AWADDR;
	output wire [7:0] sum_4_m_axi_gmem_AWLEN;
	output wire [2:0] sum_4_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_4_m_axi_gmem_AWBURST;
	output wire sum_4_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_4_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_4_m_axi_gmem_AWPROT;
	output wire [3:0] sum_4_m_axi_gmem_AWQOS;
	output wire [3:0] sum_4_m_axi_gmem_AWREGION;
	output wire sum_4_m_axi_gmem_AWUSER;
	input sum_4_m_axi_gmem_WREADY;
	output wire sum_4_m_axi_gmem_WVALID;
	output wire [31:0] sum_4_m_axi_gmem_WDATA;
	output wire [3:0] sum_4_m_axi_gmem_WSTRB;
	output wire sum_4_m_axi_gmem_WLAST;
	output wire sum_4_m_axi_gmem_WUSER;
	output wire sum_4_m_axi_gmem_BREADY;
	input sum_4_m_axi_gmem_BVALID;
	input sum_4_m_axi_gmem_BID;
	input [1:0] sum_4_m_axi_gmem_BRESP;
	input sum_4_m_axi_gmem_BUSER;
	output wire sum_4_s_axi_control_ARREADY;
	input sum_4_s_axi_control_ARVALID;
	input [4:0] sum_4_s_axi_control_ARADDR;
	input sum_4_s_axi_control_RREADY;
	output wire sum_4_s_axi_control_RVALID;
	output wire [31:0] sum_4_s_axi_control_RDATA;
	output wire [1:0] sum_4_s_axi_control_RRESP;
	output wire sum_4_s_axi_control_AWREADY;
	input sum_4_s_axi_control_AWVALID;
	input [4:0] sum_4_s_axi_control_AWADDR;
	output wire sum_4_s_axi_control_WREADY;
	input sum_4_s_axi_control_WVALID;
	input [31:0] sum_4_s_axi_control_WDATA;
	input [3:0] sum_4_s_axi_control_WSTRB;
	input sum_4_s_axi_control_BREADY;
	output wire sum_4_s_axi_control_BVALID;
	output wire [1:0] sum_4_s_axi_control_BRESP;
	input sum_5_m_axi_gmem_ARREADY;
	output wire sum_5_m_axi_gmem_ARVALID;
	output wire sum_5_m_axi_gmem_ARID;
	output wire [63:0] sum_5_m_axi_gmem_ARADDR;
	output wire [7:0] sum_5_m_axi_gmem_ARLEN;
	output wire [2:0] sum_5_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_5_m_axi_gmem_ARBURST;
	output wire sum_5_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_5_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_5_m_axi_gmem_ARPROT;
	output wire [3:0] sum_5_m_axi_gmem_ARQOS;
	output wire [3:0] sum_5_m_axi_gmem_ARREGION;
	output wire sum_5_m_axi_gmem_ARUSER;
	output wire sum_5_m_axi_gmem_RREADY;
	input sum_5_m_axi_gmem_RVALID;
	input sum_5_m_axi_gmem_RID;
	input [31:0] sum_5_m_axi_gmem_RDATA;
	input [1:0] sum_5_m_axi_gmem_RRESP;
	input sum_5_m_axi_gmem_RLAST;
	input sum_5_m_axi_gmem_RUSER;
	input sum_5_m_axi_gmem_AWREADY;
	output wire sum_5_m_axi_gmem_AWVALID;
	output wire sum_5_m_axi_gmem_AWID;
	output wire [63:0] sum_5_m_axi_gmem_AWADDR;
	output wire [7:0] sum_5_m_axi_gmem_AWLEN;
	output wire [2:0] sum_5_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_5_m_axi_gmem_AWBURST;
	output wire sum_5_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_5_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_5_m_axi_gmem_AWPROT;
	output wire [3:0] sum_5_m_axi_gmem_AWQOS;
	output wire [3:0] sum_5_m_axi_gmem_AWREGION;
	output wire sum_5_m_axi_gmem_AWUSER;
	input sum_5_m_axi_gmem_WREADY;
	output wire sum_5_m_axi_gmem_WVALID;
	output wire [31:0] sum_5_m_axi_gmem_WDATA;
	output wire [3:0] sum_5_m_axi_gmem_WSTRB;
	output wire sum_5_m_axi_gmem_WLAST;
	output wire sum_5_m_axi_gmem_WUSER;
	output wire sum_5_m_axi_gmem_BREADY;
	input sum_5_m_axi_gmem_BVALID;
	input sum_5_m_axi_gmem_BID;
	input [1:0] sum_5_m_axi_gmem_BRESP;
	input sum_5_m_axi_gmem_BUSER;
	output wire sum_5_s_axi_control_ARREADY;
	input sum_5_s_axi_control_ARVALID;
	input [4:0] sum_5_s_axi_control_ARADDR;
	input sum_5_s_axi_control_RREADY;
	output wire sum_5_s_axi_control_RVALID;
	output wire [31:0] sum_5_s_axi_control_RDATA;
	output wire [1:0] sum_5_s_axi_control_RRESP;
	output wire sum_5_s_axi_control_AWREADY;
	input sum_5_s_axi_control_AWVALID;
	input [4:0] sum_5_s_axi_control_AWADDR;
	output wire sum_5_s_axi_control_WREADY;
	input sum_5_s_axi_control_WVALID;
	input [31:0] sum_5_s_axi_control_WDATA;
	input [3:0] sum_5_s_axi_control_WSTRB;
	input sum_5_s_axi_control_BREADY;
	output wire sum_5_s_axi_control_BVALID;
	output wire [1:0] sum_5_s_axi_control_BRESP;
	input sum_6_m_axi_gmem_ARREADY;
	output wire sum_6_m_axi_gmem_ARVALID;
	output wire sum_6_m_axi_gmem_ARID;
	output wire [63:0] sum_6_m_axi_gmem_ARADDR;
	output wire [7:0] sum_6_m_axi_gmem_ARLEN;
	output wire [2:0] sum_6_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_6_m_axi_gmem_ARBURST;
	output wire sum_6_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_6_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_6_m_axi_gmem_ARPROT;
	output wire [3:0] sum_6_m_axi_gmem_ARQOS;
	output wire [3:0] sum_6_m_axi_gmem_ARREGION;
	output wire sum_6_m_axi_gmem_ARUSER;
	output wire sum_6_m_axi_gmem_RREADY;
	input sum_6_m_axi_gmem_RVALID;
	input sum_6_m_axi_gmem_RID;
	input [31:0] sum_6_m_axi_gmem_RDATA;
	input [1:0] sum_6_m_axi_gmem_RRESP;
	input sum_6_m_axi_gmem_RLAST;
	input sum_6_m_axi_gmem_RUSER;
	input sum_6_m_axi_gmem_AWREADY;
	output wire sum_6_m_axi_gmem_AWVALID;
	output wire sum_6_m_axi_gmem_AWID;
	output wire [63:0] sum_6_m_axi_gmem_AWADDR;
	output wire [7:0] sum_6_m_axi_gmem_AWLEN;
	output wire [2:0] sum_6_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_6_m_axi_gmem_AWBURST;
	output wire sum_6_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_6_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_6_m_axi_gmem_AWPROT;
	output wire [3:0] sum_6_m_axi_gmem_AWQOS;
	output wire [3:0] sum_6_m_axi_gmem_AWREGION;
	output wire sum_6_m_axi_gmem_AWUSER;
	input sum_6_m_axi_gmem_WREADY;
	output wire sum_6_m_axi_gmem_WVALID;
	output wire [31:0] sum_6_m_axi_gmem_WDATA;
	output wire [3:0] sum_6_m_axi_gmem_WSTRB;
	output wire sum_6_m_axi_gmem_WLAST;
	output wire sum_6_m_axi_gmem_WUSER;
	output wire sum_6_m_axi_gmem_BREADY;
	input sum_6_m_axi_gmem_BVALID;
	input sum_6_m_axi_gmem_BID;
	input [1:0] sum_6_m_axi_gmem_BRESP;
	input sum_6_m_axi_gmem_BUSER;
	output wire sum_6_s_axi_control_ARREADY;
	input sum_6_s_axi_control_ARVALID;
	input [4:0] sum_6_s_axi_control_ARADDR;
	input sum_6_s_axi_control_RREADY;
	output wire sum_6_s_axi_control_RVALID;
	output wire [31:0] sum_6_s_axi_control_RDATA;
	output wire [1:0] sum_6_s_axi_control_RRESP;
	output wire sum_6_s_axi_control_AWREADY;
	input sum_6_s_axi_control_AWVALID;
	input [4:0] sum_6_s_axi_control_AWADDR;
	output wire sum_6_s_axi_control_WREADY;
	input sum_6_s_axi_control_WVALID;
	input [31:0] sum_6_s_axi_control_WDATA;
	input [3:0] sum_6_s_axi_control_WSTRB;
	input sum_6_s_axi_control_BREADY;
	output wire sum_6_s_axi_control_BVALID;
	output wire [1:0] sum_6_s_axi_control_BRESP;
	input sum_7_m_axi_gmem_ARREADY;
	output wire sum_7_m_axi_gmem_ARVALID;
	output wire sum_7_m_axi_gmem_ARID;
	output wire [63:0] sum_7_m_axi_gmem_ARADDR;
	output wire [7:0] sum_7_m_axi_gmem_ARLEN;
	output wire [2:0] sum_7_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_7_m_axi_gmem_ARBURST;
	output wire sum_7_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_7_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_7_m_axi_gmem_ARPROT;
	output wire [3:0] sum_7_m_axi_gmem_ARQOS;
	output wire [3:0] sum_7_m_axi_gmem_ARREGION;
	output wire sum_7_m_axi_gmem_ARUSER;
	output wire sum_7_m_axi_gmem_RREADY;
	input sum_7_m_axi_gmem_RVALID;
	input sum_7_m_axi_gmem_RID;
	input [31:0] sum_7_m_axi_gmem_RDATA;
	input [1:0] sum_7_m_axi_gmem_RRESP;
	input sum_7_m_axi_gmem_RLAST;
	input sum_7_m_axi_gmem_RUSER;
	input sum_7_m_axi_gmem_AWREADY;
	output wire sum_7_m_axi_gmem_AWVALID;
	output wire sum_7_m_axi_gmem_AWID;
	output wire [63:0] sum_7_m_axi_gmem_AWADDR;
	output wire [7:0] sum_7_m_axi_gmem_AWLEN;
	output wire [2:0] sum_7_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_7_m_axi_gmem_AWBURST;
	output wire sum_7_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_7_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_7_m_axi_gmem_AWPROT;
	output wire [3:0] sum_7_m_axi_gmem_AWQOS;
	output wire [3:0] sum_7_m_axi_gmem_AWREGION;
	output wire sum_7_m_axi_gmem_AWUSER;
	input sum_7_m_axi_gmem_WREADY;
	output wire sum_7_m_axi_gmem_WVALID;
	output wire [31:0] sum_7_m_axi_gmem_WDATA;
	output wire [3:0] sum_7_m_axi_gmem_WSTRB;
	output wire sum_7_m_axi_gmem_WLAST;
	output wire sum_7_m_axi_gmem_WUSER;
	output wire sum_7_m_axi_gmem_BREADY;
	input sum_7_m_axi_gmem_BVALID;
	input sum_7_m_axi_gmem_BID;
	input [1:0] sum_7_m_axi_gmem_BRESP;
	input sum_7_m_axi_gmem_BUSER;
	output wire sum_7_s_axi_control_ARREADY;
	input sum_7_s_axi_control_ARVALID;
	input [4:0] sum_7_s_axi_control_ARADDR;
	input sum_7_s_axi_control_RREADY;
	output wire sum_7_s_axi_control_RVALID;
	output wire [31:0] sum_7_s_axi_control_RDATA;
	output wire [1:0] sum_7_s_axi_control_RRESP;
	output wire sum_7_s_axi_control_AWREADY;
	input sum_7_s_axi_control_AWVALID;
	input [4:0] sum_7_s_axi_control_AWADDR;
	output wire sum_7_s_axi_control_WREADY;
	input sum_7_s_axi_control_WVALID;
	input [31:0] sum_7_s_axi_control_WDATA;
	input [3:0] sum_7_s_axi_control_WSTRB;
	input sum_7_s_axi_control_BREADY;
	output wire sum_7_s_axi_control_BVALID;
	output wire [1:0] sum_7_s_axi_control_BRESP;
	input sum_8_m_axi_gmem_ARREADY;
	output wire sum_8_m_axi_gmem_ARVALID;
	output wire sum_8_m_axi_gmem_ARID;
	output wire [63:0] sum_8_m_axi_gmem_ARADDR;
	output wire [7:0] sum_8_m_axi_gmem_ARLEN;
	output wire [2:0] sum_8_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_8_m_axi_gmem_ARBURST;
	output wire sum_8_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_8_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_8_m_axi_gmem_ARPROT;
	output wire [3:0] sum_8_m_axi_gmem_ARQOS;
	output wire [3:0] sum_8_m_axi_gmem_ARREGION;
	output wire sum_8_m_axi_gmem_ARUSER;
	output wire sum_8_m_axi_gmem_RREADY;
	input sum_8_m_axi_gmem_RVALID;
	input sum_8_m_axi_gmem_RID;
	input [31:0] sum_8_m_axi_gmem_RDATA;
	input [1:0] sum_8_m_axi_gmem_RRESP;
	input sum_8_m_axi_gmem_RLAST;
	input sum_8_m_axi_gmem_RUSER;
	input sum_8_m_axi_gmem_AWREADY;
	output wire sum_8_m_axi_gmem_AWVALID;
	output wire sum_8_m_axi_gmem_AWID;
	output wire [63:0] sum_8_m_axi_gmem_AWADDR;
	output wire [7:0] sum_8_m_axi_gmem_AWLEN;
	output wire [2:0] sum_8_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_8_m_axi_gmem_AWBURST;
	output wire sum_8_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_8_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_8_m_axi_gmem_AWPROT;
	output wire [3:0] sum_8_m_axi_gmem_AWQOS;
	output wire [3:0] sum_8_m_axi_gmem_AWREGION;
	output wire sum_8_m_axi_gmem_AWUSER;
	input sum_8_m_axi_gmem_WREADY;
	output wire sum_8_m_axi_gmem_WVALID;
	output wire [31:0] sum_8_m_axi_gmem_WDATA;
	output wire [3:0] sum_8_m_axi_gmem_WSTRB;
	output wire sum_8_m_axi_gmem_WLAST;
	output wire sum_8_m_axi_gmem_WUSER;
	output wire sum_8_m_axi_gmem_BREADY;
	input sum_8_m_axi_gmem_BVALID;
	input sum_8_m_axi_gmem_BID;
	input [1:0] sum_8_m_axi_gmem_BRESP;
	input sum_8_m_axi_gmem_BUSER;
	output wire sum_8_s_axi_control_ARREADY;
	input sum_8_s_axi_control_ARVALID;
	input [4:0] sum_8_s_axi_control_ARADDR;
	input sum_8_s_axi_control_RREADY;
	output wire sum_8_s_axi_control_RVALID;
	output wire [31:0] sum_8_s_axi_control_RDATA;
	output wire [1:0] sum_8_s_axi_control_RRESP;
	output wire sum_8_s_axi_control_AWREADY;
	input sum_8_s_axi_control_AWVALID;
	input [4:0] sum_8_s_axi_control_AWADDR;
	output wire sum_8_s_axi_control_WREADY;
	input sum_8_s_axi_control_WVALID;
	input [31:0] sum_8_s_axi_control_WDATA;
	input [3:0] sum_8_s_axi_control_WSTRB;
	input sum_8_s_axi_control_BREADY;
	output wire sum_8_s_axi_control_BVALID;
	output wire [1:0] sum_8_s_axi_control_BRESP;
	input sum_9_m_axi_gmem_ARREADY;
	output wire sum_9_m_axi_gmem_ARVALID;
	output wire sum_9_m_axi_gmem_ARID;
	output wire [63:0] sum_9_m_axi_gmem_ARADDR;
	output wire [7:0] sum_9_m_axi_gmem_ARLEN;
	output wire [2:0] sum_9_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_9_m_axi_gmem_ARBURST;
	output wire sum_9_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_9_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_9_m_axi_gmem_ARPROT;
	output wire [3:0] sum_9_m_axi_gmem_ARQOS;
	output wire [3:0] sum_9_m_axi_gmem_ARREGION;
	output wire sum_9_m_axi_gmem_ARUSER;
	output wire sum_9_m_axi_gmem_RREADY;
	input sum_9_m_axi_gmem_RVALID;
	input sum_9_m_axi_gmem_RID;
	input [31:0] sum_9_m_axi_gmem_RDATA;
	input [1:0] sum_9_m_axi_gmem_RRESP;
	input sum_9_m_axi_gmem_RLAST;
	input sum_9_m_axi_gmem_RUSER;
	input sum_9_m_axi_gmem_AWREADY;
	output wire sum_9_m_axi_gmem_AWVALID;
	output wire sum_9_m_axi_gmem_AWID;
	output wire [63:0] sum_9_m_axi_gmem_AWADDR;
	output wire [7:0] sum_9_m_axi_gmem_AWLEN;
	output wire [2:0] sum_9_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_9_m_axi_gmem_AWBURST;
	output wire sum_9_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_9_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_9_m_axi_gmem_AWPROT;
	output wire [3:0] sum_9_m_axi_gmem_AWQOS;
	output wire [3:0] sum_9_m_axi_gmem_AWREGION;
	output wire sum_9_m_axi_gmem_AWUSER;
	input sum_9_m_axi_gmem_WREADY;
	output wire sum_9_m_axi_gmem_WVALID;
	output wire [31:0] sum_9_m_axi_gmem_WDATA;
	output wire [3:0] sum_9_m_axi_gmem_WSTRB;
	output wire sum_9_m_axi_gmem_WLAST;
	output wire sum_9_m_axi_gmem_WUSER;
	output wire sum_9_m_axi_gmem_BREADY;
	input sum_9_m_axi_gmem_BVALID;
	input sum_9_m_axi_gmem_BID;
	input [1:0] sum_9_m_axi_gmem_BRESP;
	input sum_9_m_axi_gmem_BUSER;
	output wire sum_9_s_axi_control_ARREADY;
	input sum_9_s_axi_control_ARVALID;
	input [4:0] sum_9_s_axi_control_ARADDR;
	input sum_9_s_axi_control_RREADY;
	output wire sum_9_s_axi_control_RVALID;
	output wire [31:0] sum_9_s_axi_control_RDATA;
	output wire [1:0] sum_9_s_axi_control_RRESP;
	output wire sum_9_s_axi_control_AWREADY;
	input sum_9_s_axi_control_AWVALID;
	input [4:0] sum_9_s_axi_control_AWADDR;
	output wire sum_9_s_axi_control_WREADY;
	input sum_9_s_axi_control_WVALID;
	input [31:0] sum_9_s_axi_control_WDATA;
	input [3:0] sum_9_s_axi_control_WSTRB;
	input sum_9_s_axi_control_BREADY;
	output wire sum_9_s_axi_control_BVALID;
	output wire [1:0] sum_9_s_axi_control_BRESP;
	input sum_10_m_axi_gmem_ARREADY;
	output wire sum_10_m_axi_gmem_ARVALID;
	output wire sum_10_m_axi_gmem_ARID;
	output wire [63:0] sum_10_m_axi_gmem_ARADDR;
	output wire [7:0] sum_10_m_axi_gmem_ARLEN;
	output wire [2:0] sum_10_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_10_m_axi_gmem_ARBURST;
	output wire sum_10_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_10_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_10_m_axi_gmem_ARPROT;
	output wire [3:0] sum_10_m_axi_gmem_ARQOS;
	output wire [3:0] sum_10_m_axi_gmem_ARREGION;
	output wire sum_10_m_axi_gmem_ARUSER;
	output wire sum_10_m_axi_gmem_RREADY;
	input sum_10_m_axi_gmem_RVALID;
	input sum_10_m_axi_gmem_RID;
	input [31:0] sum_10_m_axi_gmem_RDATA;
	input [1:0] sum_10_m_axi_gmem_RRESP;
	input sum_10_m_axi_gmem_RLAST;
	input sum_10_m_axi_gmem_RUSER;
	input sum_10_m_axi_gmem_AWREADY;
	output wire sum_10_m_axi_gmem_AWVALID;
	output wire sum_10_m_axi_gmem_AWID;
	output wire [63:0] sum_10_m_axi_gmem_AWADDR;
	output wire [7:0] sum_10_m_axi_gmem_AWLEN;
	output wire [2:0] sum_10_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_10_m_axi_gmem_AWBURST;
	output wire sum_10_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_10_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_10_m_axi_gmem_AWPROT;
	output wire [3:0] sum_10_m_axi_gmem_AWQOS;
	output wire [3:0] sum_10_m_axi_gmem_AWREGION;
	output wire sum_10_m_axi_gmem_AWUSER;
	input sum_10_m_axi_gmem_WREADY;
	output wire sum_10_m_axi_gmem_WVALID;
	output wire [31:0] sum_10_m_axi_gmem_WDATA;
	output wire [3:0] sum_10_m_axi_gmem_WSTRB;
	output wire sum_10_m_axi_gmem_WLAST;
	output wire sum_10_m_axi_gmem_WUSER;
	output wire sum_10_m_axi_gmem_BREADY;
	input sum_10_m_axi_gmem_BVALID;
	input sum_10_m_axi_gmem_BID;
	input [1:0] sum_10_m_axi_gmem_BRESP;
	input sum_10_m_axi_gmem_BUSER;
	output wire sum_10_s_axi_control_ARREADY;
	input sum_10_s_axi_control_ARVALID;
	input [4:0] sum_10_s_axi_control_ARADDR;
	input sum_10_s_axi_control_RREADY;
	output wire sum_10_s_axi_control_RVALID;
	output wire [31:0] sum_10_s_axi_control_RDATA;
	output wire [1:0] sum_10_s_axi_control_RRESP;
	output wire sum_10_s_axi_control_AWREADY;
	input sum_10_s_axi_control_AWVALID;
	input [4:0] sum_10_s_axi_control_AWADDR;
	output wire sum_10_s_axi_control_WREADY;
	input sum_10_s_axi_control_WVALID;
	input [31:0] sum_10_s_axi_control_WDATA;
	input [3:0] sum_10_s_axi_control_WSTRB;
	input sum_10_s_axi_control_BREADY;
	output wire sum_10_s_axi_control_BVALID;
	output wire [1:0] sum_10_s_axi_control_BRESP;
	input sum_11_m_axi_gmem_ARREADY;
	output wire sum_11_m_axi_gmem_ARVALID;
	output wire sum_11_m_axi_gmem_ARID;
	output wire [63:0] sum_11_m_axi_gmem_ARADDR;
	output wire [7:0] sum_11_m_axi_gmem_ARLEN;
	output wire [2:0] sum_11_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_11_m_axi_gmem_ARBURST;
	output wire sum_11_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_11_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_11_m_axi_gmem_ARPROT;
	output wire [3:0] sum_11_m_axi_gmem_ARQOS;
	output wire [3:0] sum_11_m_axi_gmem_ARREGION;
	output wire sum_11_m_axi_gmem_ARUSER;
	output wire sum_11_m_axi_gmem_RREADY;
	input sum_11_m_axi_gmem_RVALID;
	input sum_11_m_axi_gmem_RID;
	input [31:0] sum_11_m_axi_gmem_RDATA;
	input [1:0] sum_11_m_axi_gmem_RRESP;
	input sum_11_m_axi_gmem_RLAST;
	input sum_11_m_axi_gmem_RUSER;
	input sum_11_m_axi_gmem_AWREADY;
	output wire sum_11_m_axi_gmem_AWVALID;
	output wire sum_11_m_axi_gmem_AWID;
	output wire [63:0] sum_11_m_axi_gmem_AWADDR;
	output wire [7:0] sum_11_m_axi_gmem_AWLEN;
	output wire [2:0] sum_11_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_11_m_axi_gmem_AWBURST;
	output wire sum_11_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_11_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_11_m_axi_gmem_AWPROT;
	output wire [3:0] sum_11_m_axi_gmem_AWQOS;
	output wire [3:0] sum_11_m_axi_gmem_AWREGION;
	output wire sum_11_m_axi_gmem_AWUSER;
	input sum_11_m_axi_gmem_WREADY;
	output wire sum_11_m_axi_gmem_WVALID;
	output wire [31:0] sum_11_m_axi_gmem_WDATA;
	output wire [3:0] sum_11_m_axi_gmem_WSTRB;
	output wire sum_11_m_axi_gmem_WLAST;
	output wire sum_11_m_axi_gmem_WUSER;
	output wire sum_11_m_axi_gmem_BREADY;
	input sum_11_m_axi_gmem_BVALID;
	input sum_11_m_axi_gmem_BID;
	input [1:0] sum_11_m_axi_gmem_BRESP;
	input sum_11_m_axi_gmem_BUSER;
	output wire sum_11_s_axi_control_ARREADY;
	input sum_11_s_axi_control_ARVALID;
	input [4:0] sum_11_s_axi_control_ARADDR;
	input sum_11_s_axi_control_RREADY;
	output wire sum_11_s_axi_control_RVALID;
	output wire [31:0] sum_11_s_axi_control_RDATA;
	output wire [1:0] sum_11_s_axi_control_RRESP;
	output wire sum_11_s_axi_control_AWREADY;
	input sum_11_s_axi_control_AWVALID;
	input [4:0] sum_11_s_axi_control_AWADDR;
	output wire sum_11_s_axi_control_WREADY;
	input sum_11_s_axi_control_WVALID;
	input [31:0] sum_11_s_axi_control_WDATA;
	input [3:0] sum_11_s_axi_control_WSTRB;
	input sum_11_s_axi_control_BREADY;
	output wire sum_11_s_axi_control_BVALID;
	output wire [1:0] sum_11_s_axi_control_BRESP;
	input sum_12_m_axi_gmem_ARREADY;
	output wire sum_12_m_axi_gmem_ARVALID;
	output wire sum_12_m_axi_gmem_ARID;
	output wire [63:0] sum_12_m_axi_gmem_ARADDR;
	output wire [7:0] sum_12_m_axi_gmem_ARLEN;
	output wire [2:0] sum_12_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_12_m_axi_gmem_ARBURST;
	output wire sum_12_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_12_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_12_m_axi_gmem_ARPROT;
	output wire [3:0] sum_12_m_axi_gmem_ARQOS;
	output wire [3:0] sum_12_m_axi_gmem_ARREGION;
	output wire sum_12_m_axi_gmem_ARUSER;
	output wire sum_12_m_axi_gmem_RREADY;
	input sum_12_m_axi_gmem_RVALID;
	input sum_12_m_axi_gmem_RID;
	input [31:0] sum_12_m_axi_gmem_RDATA;
	input [1:0] sum_12_m_axi_gmem_RRESP;
	input sum_12_m_axi_gmem_RLAST;
	input sum_12_m_axi_gmem_RUSER;
	input sum_12_m_axi_gmem_AWREADY;
	output wire sum_12_m_axi_gmem_AWVALID;
	output wire sum_12_m_axi_gmem_AWID;
	output wire [63:0] sum_12_m_axi_gmem_AWADDR;
	output wire [7:0] sum_12_m_axi_gmem_AWLEN;
	output wire [2:0] sum_12_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_12_m_axi_gmem_AWBURST;
	output wire sum_12_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_12_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_12_m_axi_gmem_AWPROT;
	output wire [3:0] sum_12_m_axi_gmem_AWQOS;
	output wire [3:0] sum_12_m_axi_gmem_AWREGION;
	output wire sum_12_m_axi_gmem_AWUSER;
	input sum_12_m_axi_gmem_WREADY;
	output wire sum_12_m_axi_gmem_WVALID;
	output wire [31:0] sum_12_m_axi_gmem_WDATA;
	output wire [3:0] sum_12_m_axi_gmem_WSTRB;
	output wire sum_12_m_axi_gmem_WLAST;
	output wire sum_12_m_axi_gmem_WUSER;
	output wire sum_12_m_axi_gmem_BREADY;
	input sum_12_m_axi_gmem_BVALID;
	input sum_12_m_axi_gmem_BID;
	input [1:0] sum_12_m_axi_gmem_BRESP;
	input sum_12_m_axi_gmem_BUSER;
	output wire sum_12_s_axi_control_ARREADY;
	input sum_12_s_axi_control_ARVALID;
	input [4:0] sum_12_s_axi_control_ARADDR;
	input sum_12_s_axi_control_RREADY;
	output wire sum_12_s_axi_control_RVALID;
	output wire [31:0] sum_12_s_axi_control_RDATA;
	output wire [1:0] sum_12_s_axi_control_RRESP;
	output wire sum_12_s_axi_control_AWREADY;
	input sum_12_s_axi_control_AWVALID;
	input [4:0] sum_12_s_axi_control_AWADDR;
	output wire sum_12_s_axi_control_WREADY;
	input sum_12_s_axi_control_WVALID;
	input [31:0] sum_12_s_axi_control_WDATA;
	input [3:0] sum_12_s_axi_control_WSTRB;
	input sum_12_s_axi_control_BREADY;
	output wire sum_12_s_axi_control_BVALID;
	output wire [1:0] sum_12_s_axi_control_BRESP;
	input sum_13_m_axi_gmem_ARREADY;
	output wire sum_13_m_axi_gmem_ARVALID;
	output wire sum_13_m_axi_gmem_ARID;
	output wire [63:0] sum_13_m_axi_gmem_ARADDR;
	output wire [7:0] sum_13_m_axi_gmem_ARLEN;
	output wire [2:0] sum_13_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_13_m_axi_gmem_ARBURST;
	output wire sum_13_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_13_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_13_m_axi_gmem_ARPROT;
	output wire [3:0] sum_13_m_axi_gmem_ARQOS;
	output wire [3:0] sum_13_m_axi_gmem_ARREGION;
	output wire sum_13_m_axi_gmem_ARUSER;
	output wire sum_13_m_axi_gmem_RREADY;
	input sum_13_m_axi_gmem_RVALID;
	input sum_13_m_axi_gmem_RID;
	input [31:0] sum_13_m_axi_gmem_RDATA;
	input [1:0] sum_13_m_axi_gmem_RRESP;
	input sum_13_m_axi_gmem_RLAST;
	input sum_13_m_axi_gmem_RUSER;
	input sum_13_m_axi_gmem_AWREADY;
	output wire sum_13_m_axi_gmem_AWVALID;
	output wire sum_13_m_axi_gmem_AWID;
	output wire [63:0] sum_13_m_axi_gmem_AWADDR;
	output wire [7:0] sum_13_m_axi_gmem_AWLEN;
	output wire [2:0] sum_13_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_13_m_axi_gmem_AWBURST;
	output wire sum_13_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_13_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_13_m_axi_gmem_AWPROT;
	output wire [3:0] sum_13_m_axi_gmem_AWQOS;
	output wire [3:0] sum_13_m_axi_gmem_AWREGION;
	output wire sum_13_m_axi_gmem_AWUSER;
	input sum_13_m_axi_gmem_WREADY;
	output wire sum_13_m_axi_gmem_WVALID;
	output wire [31:0] sum_13_m_axi_gmem_WDATA;
	output wire [3:0] sum_13_m_axi_gmem_WSTRB;
	output wire sum_13_m_axi_gmem_WLAST;
	output wire sum_13_m_axi_gmem_WUSER;
	output wire sum_13_m_axi_gmem_BREADY;
	input sum_13_m_axi_gmem_BVALID;
	input sum_13_m_axi_gmem_BID;
	input [1:0] sum_13_m_axi_gmem_BRESP;
	input sum_13_m_axi_gmem_BUSER;
	output wire sum_13_s_axi_control_ARREADY;
	input sum_13_s_axi_control_ARVALID;
	input [4:0] sum_13_s_axi_control_ARADDR;
	input sum_13_s_axi_control_RREADY;
	output wire sum_13_s_axi_control_RVALID;
	output wire [31:0] sum_13_s_axi_control_RDATA;
	output wire [1:0] sum_13_s_axi_control_RRESP;
	output wire sum_13_s_axi_control_AWREADY;
	input sum_13_s_axi_control_AWVALID;
	input [4:0] sum_13_s_axi_control_AWADDR;
	output wire sum_13_s_axi_control_WREADY;
	input sum_13_s_axi_control_WVALID;
	input [31:0] sum_13_s_axi_control_WDATA;
	input [3:0] sum_13_s_axi_control_WSTRB;
	input sum_13_s_axi_control_BREADY;
	output wire sum_13_s_axi_control_BVALID;
	output wire [1:0] sum_13_s_axi_control_BRESP;
	input sum_14_m_axi_gmem_ARREADY;
	output wire sum_14_m_axi_gmem_ARVALID;
	output wire sum_14_m_axi_gmem_ARID;
	output wire [63:0] sum_14_m_axi_gmem_ARADDR;
	output wire [7:0] sum_14_m_axi_gmem_ARLEN;
	output wire [2:0] sum_14_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_14_m_axi_gmem_ARBURST;
	output wire sum_14_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_14_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_14_m_axi_gmem_ARPROT;
	output wire [3:0] sum_14_m_axi_gmem_ARQOS;
	output wire [3:0] sum_14_m_axi_gmem_ARREGION;
	output wire sum_14_m_axi_gmem_ARUSER;
	output wire sum_14_m_axi_gmem_RREADY;
	input sum_14_m_axi_gmem_RVALID;
	input sum_14_m_axi_gmem_RID;
	input [31:0] sum_14_m_axi_gmem_RDATA;
	input [1:0] sum_14_m_axi_gmem_RRESP;
	input sum_14_m_axi_gmem_RLAST;
	input sum_14_m_axi_gmem_RUSER;
	input sum_14_m_axi_gmem_AWREADY;
	output wire sum_14_m_axi_gmem_AWVALID;
	output wire sum_14_m_axi_gmem_AWID;
	output wire [63:0] sum_14_m_axi_gmem_AWADDR;
	output wire [7:0] sum_14_m_axi_gmem_AWLEN;
	output wire [2:0] sum_14_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_14_m_axi_gmem_AWBURST;
	output wire sum_14_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_14_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_14_m_axi_gmem_AWPROT;
	output wire [3:0] sum_14_m_axi_gmem_AWQOS;
	output wire [3:0] sum_14_m_axi_gmem_AWREGION;
	output wire sum_14_m_axi_gmem_AWUSER;
	input sum_14_m_axi_gmem_WREADY;
	output wire sum_14_m_axi_gmem_WVALID;
	output wire [31:0] sum_14_m_axi_gmem_WDATA;
	output wire [3:0] sum_14_m_axi_gmem_WSTRB;
	output wire sum_14_m_axi_gmem_WLAST;
	output wire sum_14_m_axi_gmem_WUSER;
	output wire sum_14_m_axi_gmem_BREADY;
	input sum_14_m_axi_gmem_BVALID;
	input sum_14_m_axi_gmem_BID;
	input [1:0] sum_14_m_axi_gmem_BRESP;
	input sum_14_m_axi_gmem_BUSER;
	output wire sum_14_s_axi_control_ARREADY;
	input sum_14_s_axi_control_ARVALID;
	input [4:0] sum_14_s_axi_control_ARADDR;
	input sum_14_s_axi_control_RREADY;
	output wire sum_14_s_axi_control_RVALID;
	output wire [31:0] sum_14_s_axi_control_RDATA;
	output wire [1:0] sum_14_s_axi_control_RRESP;
	output wire sum_14_s_axi_control_AWREADY;
	input sum_14_s_axi_control_AWVALID;
	input [4:0] sum_14_s_axi_control_AWADDR;
	output wire sum_14_s_axi_control_WREADY;
	input sum_14_s_axi_control_WVALID;
	input [31:0] sum_14_s_axi_control_WDATA;
	input [3:0] sum_14_s_axi_control_WSTRB;
	input sum_14_s_axi_control_BREADY;
	output wire sum_14_s_axi_control_BVALID;
	output wire [1:0] sum_14_s_axi_control_BRESP;
	input sum_15_m_axi_gmem_ARREADY;
	output wire sum_15_m_axi_gmem_ARVALID;
	output wire sum_15_m_axi_gmem_ARID;
	output wire [63:0] sum_15_m_axi_gmem_ARADDR;
	output wire [7:0] sum_15_m_axi_gmem_ARLEN;
	output wire [2:0] sum_15_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_15_m_axi_gmem_ARBURST;
	output wire sum_15_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_15_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_15_m_axi_gmem_ARPROT;
	output wire [3:0] sum_15_m_axi_gmem_ARQOS;
	output wire [3:0] sum_15_m_axi_gmem_ARREGION;
	output wire sum_15_m_axi_gmem_ARUSER;
	output wire sum_15_m_axi_gmem_RREADY;
	input sum_15_m_axi_gmem_RVALID;
	input sum_15_m_axi_gmem_RID;
	input [31:0] sum_15_m_axi_gmem_RDATA;
	input [1:0] sum_15_m_axi_gmem_RRESP;
	input sum_15_m_axi_gmem_RLAST;
	input sum_15_m_axi_gmem_RUSER;
	input sum_15_m_axi_gmem_AWREADY;
	output wire sum_15_m_axi_gmem_AWVALID;
	output wire sum_15_m_axi_gmem_AWID;
	output wire [63:0] sum_15_m_axi_gmem_AWADDR;
	output wire [7:0] sum_15_m_axi_gmem_AWLEN;
	output wire [2:0] sum_15_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_15_m_axi_gmem_AWBURST;
	output wire sum_15_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_15_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_15_m_axi_gmem_AWPROT;
	output wire [3:0] sum_15_m_axi_gmem_AWQOS;
	output wire [3:0] sum_15_m_axi_gmem_AWREGION;
	output wire sum_15_m_axi_gmem_AWUSER;
	input sum_15_m_axi_gmem_WREADY;
	output wire sum_15_m_axi_gmem_WVALID;
	output wire [31:0] sum_15_m_axi_gmem_WDATA;
	output wire [3:0] sum_15_m_axi_gmem_WSTRB;
	output wire sum_15_m_axi_gmem_WLAST;
	output wire sum_15_m_axi_gmem_WUSER;
	output wire sum_15_m_axi_gmem_BREADY;
	input sum_15_m_axi_gmem_BVALID;
	input sum_15_m_axi_gmem_BID;
	input [1:0] sum_15_m_axi_gmem_BRESP;
	input sum_15_m_axi_gmem_BUSER;
	output wire sum_15_s_axi_control_ARREADY;
	input sum_15_s_axi_control_ARVALID;
	input [4:0] sum_15_s_axi_control_ARADDR;
	input sum_15_s_axi_control_RREADY;
	output wire sum_15_s_axi_control_RVALID;
	output wire [31:0] sum_15_s_axi_control_RDATA;
	output wire [1:0] sum_15_s_axi_control_RRESP;
	output wire sum_15_s_axi_control_AWREADY;
	input sum_15_s_axi_control_AWVALID;
	input [4:0] sum_15_s_axi_control_AWADDR;
	output wire sum_15_s_axi_control_WREADY;
	input sum_15_s_axi_control_WVALID;
	input [31:0] sum_15_s_axi_control_WDATA;
	input [3:0] sum_15_s_axi_control_WSTRB;
	input sum_15_s_axi_control_BREADY;
	output wire sum_15_s_axi_control_BVALID;
	output wire [1:0] sum_15_s_axi_control_BRESP;
	input sum_16_m_axi_gmem_ARREADY;
	output wire sum_16_m_axi_gmem_ARVALID;
	output wire sum_16_m_axi_gmem_ARID;
	output wire [63:0] sum_16_m_axi_gmem_ARADDR;
	output wire [7:0] sum_16_m_axi_gmem_ARLEN;
	output wire [2:0] sum_16_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_16_m_axi_gmem_ARBURST;
	output wire sum_16_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_16_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_16_m_axi_gmem_ARPROT;
	output wire [3:0] sum_16_m_axi_gmem_ARQOS;
	output wire [3:0] sum_16_m_axi_gmem_ARREGION;
	output wire sum_16_m_axi_gmem_ARUSER;
	output wire sum_16_m_axi_gmem_RREADY;
	input sum_16_m_axi_gmem_RVALID;
	input sum_16_m_axi_gmem_RID;
	input [31:0] sum_16_m_axi_gmem_RDATA;
	input [1:0] sum_16_m_axi_gmem_RRESP;
	input sum_16_m_axi_gmem_RLAST;
	input sum_16_m_axi_gmem_RUSER;
	input sum_16_m_axi_gmem_AWREADY;
	output wire sum_16_m_axi_gmem_AWVALID;
	output wire sum_16_m_axi_gmem_AWID;
	output wire [63:0] sum_16_m_axi_gmem_AWADDR;
	output wire [7:0] sum_16_m_axi_gmem_AWLEN;
	output wire [2:0] sum_16_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_16_m_axi_gmem_AWBURST;
	output wire sum_16_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_16_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_16_m_axi_gmem_AWPROT;
	output wire [3:0] sum_16_m_axi_gmem_AWQOS;
	output wire [3:0] sum_16_m_axi_gmem_AWREGION;
	output wire sum_16_m_axi_gmem_AWUSER;
	input sum_16_m_axi_gmem_WREADY;
	output wire sum_16_m_axi_gmem_WVALID;
	output wire [31:0] sum_16_m_axi_gmem_WDATA;
	output wire [3:0] sum_16_m_axi_gmem_WSTRB;
	output wire sum_16_m_axi_gmem_WLAST;
	output wire sum_16_m_axi_gmem_WUSER;
	output wire sum_16_m_axi_gmem_BREADY;
	input sum_16_m_axi_gmem_BVALID;
	input sum_16_m_axi_gmem_BID;
	input [1:0] sum_16_m_axi_gmem_BRESP;
	input sum_16_m_axi_gmem_BUSER;
	output wire sum_16_s_axi_control_ARREADY;
	input sum_16_s_axi_control_ARVALID;
	input [4:0] sum_16_s_axi_control_ARADDR;
	input sum_16_s_axi_control_RREADY;
	output wire sum_16_s_axi_control_RVALID;
	output wire [31:0] sum_16_s_axi_control_RDATA;
	output wire [1:0] sum_16_s_axi_control_RRESP;
	output wire sum_16_s_axi_control_AWREADY;
	input sum_16_s_axi_control_AWVALID;
	input [4:0] sum_16_s_axi_control_AWADDR;
	output wire sum_16_s_axi_control_WREADY;
	input sum_16_s_axi_control_WVALID;
	input [31:0] sum_16_s_axi_control_WDATA;
	input [3:0] sum_16_s_axi_control_WSTRB;
	input sum_16_s_axi_control_BREADY;
	output wire sum_16_s_axi_control_BVALID;
	output wire [1:0] sum_16_s_axi_control_BRESP;
	input sum_17_m_axi_gmem_ARREADY;
	output wire sum_17_m_axi_gmem_ARVALID;
	output wire sum_17_m_axi_gmem_ARID;
	output wire [63:0] sum_17_m_axi_gmem_ARADDR;
	output wire [7:0] sum_17_m_axi_gmem_ARLEN;
	output wire [2:0] sum_17_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_17_m_axi_gmem_ARBURST;
	output wire sum_17_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_17_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_17_m_axi_gmem_ARPROT;
	output wire [3:0] sum_17_m_axi_gmem_ARQOS;
	output wire [3:0] sum_17_m_axi_gmem_ARREGION;
	output wire sum_17_m_axi_gmem_ARUSER;
	output wire sum_17_m_axi_gmem_RREADY;
	input sum_17_m_axi_gmem_RVALID;
	input sum_17_m_axi_gmem_RID;
	input [31:0] sum_17_m_axi_gmem_RDATA;
	input [1:0] sum_17_m_axi_gmem_RRESP;
	input sum_17_m_axi_gmem_RLAST;
	input sum_17_m_axi_gmem_RUSER;
	input sum_17_m_axi_gmem_AWREADY;
	output wire sum_17_m_axi_gmem_AWVALID;
	output wire sum_17_m_axi_gmem_AWID;
	output wire [63:0] sum_17_m_axi_gmem_AWADDR;
	output wire [7:0] sum_17_m_axi_gmem_AWLEN;
	output wire [2:0] sum_17_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_17_m_axi_gmem_AWBURST;
	output wire sum_17_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_17_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_17_m_axi_gmem_AWPROT;
	output wire [3:0] sum_17_m_axi_gmem_AWQOS;
	output wire [3:0] sum_17_m_axi_gmem_AWREGION;
	output wire sum_17_m_axi_gmem_AWUSER;
	input sum_17_m_axi_gmem_WREADY;
	output wire sum_17_m_axi_gmem_WVALID;
	output wire [31:0] sum_17_m_axi_gmem_WDATA;
	output wire [3:0] sum_17_m_axi_gmem_WSTRB;
	output wire sum_17_m_axi_gmem_WLAST;
	output wire sum_17_m_axi_gmem_WUSER;
	output wire sum_17_m_axi_gmem_BREADY;
	input sum_17_m_axi_gmem_BVALID;
	input sum_17_m_axi_gmem_BID;
	input [1:0] sum_17_m_axi_gmem_BRESP;
	input sum_17_m_axi_gmem_BUSER;
	output wire sum_17_s_axi_control_ARREADY;
	input sum_17_s_axi_control_ARVALID;
	input [4:0] sum_17_s_axi_control_ARADDR;
	input sum_17_s_axi_control_RREADY;
	output wire sum_17_s_axi_control_RVALID;
	output wire [31:0] sum_17_s_axi_control_RDATA;
	output wire [1:0] sum_17_s_axi_control_RRESP;
	output wire sum_17_s_axi_control_AWREADY;
	input sum_17_s_axi_control_AWVALID;
	input [4:0] sum_17_s_axi_control_AWADDR;
	output wire sum_17_s_axi_control_WREADY;
	input sum_17_s_axi_control_WVALID;
	input [31:0] sum_17_s_axi_control_WDATA;
	input [3:0] sum_17_s_axi_control_WSTRB;
	input sum_17_s_axi_control_BREADY;
	output wire sum_17_s_axi_control_BVALID;
	output wire [1:0] sum_17_s_axi_control_BRESP;
	input sum_18_m_axi_gmem_ARREADY;
	output wire sum_18_m_axi_gmem_ARVALID;
	output wire sum_18_m_axi_gmem_ARID;
	output wire [63:0] sum_18_m_axi_gmem_ARADDR;
	output wire [7:0] sum_18_m_axi_gmem_ARLEN;
	output wire [2:0] sum_18_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_18_m_axi_gmem_ARBURST;
	output wire sum_18_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_18_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_18_m_axi_gmem_ARPROT;
	output wire [3:0] sum_18_m_axi_gmem_ARQOS;
	output wire [3:0] sum_18_m_axi_gmem_ARREGION;
	output wire sum_18_m_axi_gmem_ARUSER;
	output wire sum_18_m_axi_gmem_RREADY;
	input sum_18_m_axi_gmem_RVALID;
	input sum_18_m_axi_gmem_RID;
	input [31:0] sum_18_m_axi_gmem_RDATA;
	input [1:0] sum_18_m_axi_gmem_RRESP;
	input sum_18_m_axi_gmem_RLAST;
	input sum_18_m_axi_gmem_RUSER;
	input sum_18_m_axi_gmem_AWREADY;
	output wire sum_18_m_axi_gmem_AWVALID;
	output wire sum_18_m_axi_gmem_AWID;
	output wire [63:0] sum_18_m_axi_gmem_AWADDR;
	output wire [7:0] sum_18_m_axi_gmem_AWLEN;
	output wire [2:0] sum_18_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_18_m_axi_gmem_AWBURST;
	output wire sum_18_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_18_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_18_m_axi_gmem_AWPROT;
	output wire [3:0] sum_18_m_axi_gmem_AWQOS;
	output wire [3:0] sum_18_m_axi_gmem_AWREGION;
	output wire sum_18_m_axi_gmem_AWUSER;
	input sum_18_m_axi_gmem_WREADY;
	output wire sum_18_m_axi_gmem_WVALID;
	output wire [31:0] sum_18_m_axi_gmem_WDATA;
	output wire [3:0] sum_18_m_axi_gmem_WSTRB;
	output wire sum_18_m_axi_gmem_WLAST;
	output wire sum_18_m_axi_gmem_WUSER;
	output wire sum_18_m_axi_gmem_BREADY;
	input sum_18_m_axi_gmem_BVALID;
	input sum_18_m_axi_gmem_BID;
	input [1:0] sum_18_m_axi_gmem_BRESP;
	input sum_18_m_axi_gmem_BUSER;
	output wire sum_18_s_axi_control_ARREADY;
	input sum_18_s_axi_control_ARVALID;
	input [4:0] sum_18_s_axi_control_ARADDR;
	input sum_18_s_axi_control_RREADY;
	output wire sum_18_s_axi_control_RVALID;
	output wire [31:0] sum_18_s_axi_control_RDATA;
	output wire [1:0] sum_18_s_axi_control_RRESP;
	output wire sum_18_s_axi_control_AWREADY;
	input sum_18_s_axi_control_AWVALID;
	input [4:0] sum_18_s_axi_control_AWADDR;
	output wire sum_18_s_axi_control_WREADY;
	input sum_18_s_axi_control_WVALID;
	input [31:0] sum_18_s_axi_control_WDATA;
	input [3:0] sum_18_s_axi_control_WSTRB;
	input sum_18_s_axi_control_BREADY;
	output wire sum_18_s_axi_control_BVALID;
	output wire [1:0] sum_18_s_axi_control_BRESP;
	input sum_19_m_axi_gmem_ARREADY;
	output wire sum_19_m_axi_gmem_ARVALID;
	output wire sum_19_m_axi_gmem_ARID;
	output wire [63:0] sum_19_m_axi_gmem_ARADDR;
	output wire [7:0] sum_19_m_axi_gmem_ARLEN;
	output wire [2:0] sum_19_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_19_m_axi_gmem_ARBURST;
	output wire sum_19_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_19_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_19_m_axi_gmem_ARPROT;
	output wire [3:0] sum_19_m_axi_gmem_ARQOS;
	output wire [3:0] sum_19_m_axi_gmem_ARREGION;
	output wire sum_19_m_axi_gmem_ARUSER;
	output wire sum_19_m_axi_gmem_RREADY;
	input sum_19_m_axi_gmem_RVALID;
	input sum_19_m_axi_gmem_RID;
	input [31:0] sum_19_m_axi_gmem_RDATA;
	input [1:0] sum_19_m_axi_gmem_RRESP;
	input sum_19_m_axi_gmem_RLAST;
	input sum_19_m_axi_gmem_RUSER;
	input sum_19_m_axi_gmem_AWREADY;
	output wire sum_19_m_axi_gmem_AWVALID;
	output wire sum_19_m_axi_gmem_AWID;
	output wire [63:0] sum_19_m_axi_gmem_AWADDR;
	output wire [7:0] sum_19_m_axi_gmem_AWLEN;
	output wire [2:0] sum_19_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_19_m_axi_gmem_AWBURST;
	output wire sum_19_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_19_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_19_m_axi_gmem_AWPROT;
	output wire [3:0] sum_19_m_axi_gmem_AWQOS;
	output wire [3:0] sum_19_m_axi_gmem_AWREGION;
	output wire sum_19_m_axi_gmem_AWUSER;
	input sum_19_m_axi_gmem_WREADY;
	output wire sum_19_m_axi_gmem_WVALID;
	output wire [31:0] sum_19_m_axi_gmem_WDATA;
	output wire [3:0] sum_19_m_axi_gmem_WSTRB;
	output wire sum_19_m_axi_gmem_WLAST;
	output wire sum_19_m_axi_gmem_WUSER;
	output wire sum_19_m_axi_gmem_BREADY;
	input sum_19_m_axi_gmem_BVALID;
	input sum_19_m_axi_gmem_BID;
	input [1:0] sum_19_m_axi_gmem_BRESP;
	input sum_19_m_axi_gmem_BUSER;
	output wire sum_19_s_axi_control_ARREADY;
	input sum_19_s_axi_control_ARVALID;
	input [4:0] sum_19_s_axi_control_ARADDR;
	input sum_19_s_axi_control_RREADY;
	output wire sum_19_s_axi_control_RVALID;
	output wire [31:0] sum_19_s_axi_control_RDATA;
	output wire [1:0] sum_19_s_axi_control_RRESP;
	output wire sum_19_s_axi_control_AWREADY;
	input sum_19_s_axi_control_AWVALID;
	input [4:0] sum_19_s_axi_control_AWADDR;
	output wire sum_19_s_axi_control_WREADY;
	input sum_19_s_axi_control_WVALID;
	input [31:0] sum_19_s_axi_control_WDATA;
	input [3:0] sum_19_s_axi_control_WSTRB;
	input sum_19_s_axi_control_BREADY;
	output wire sum_19_s_axi_control_BVALID;
	output wire [1:0] sum_19_s_axi_control_BRESP;
	input sum_20_m_axi_gmem_ARREADY;
	output wire sum_20_m_axi_gmem_ARVALID;
	output wire sum_20_m_axi_gmem_ARID;
	output wire [63:0] sum_20_m_axi_gmem_ARADDR;
	output wire [7:0] sum_20_m_axi_gmem_ARLEN;
	output wire [2:0] sum_20_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_20_m_axi_gmem_ARBURST;
	output wire sum_20_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_20_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_20_m_axi_gmem_ARPROT;
	output wire [3:0] sum_20_m_axi_gmem_ARQOS;
	output wire [3:0] sum_20_m_axi_gmem_ARREGION;
	output wire sum_20_m_axi_gmem_ARUSER;
	output wire sum_20_m_axi_gmem_RREADY;
	input sum_20_m_axi_gmem_RVALID;
	input sum_20_m_axi_gmem_RID;
	input [31:0] sum_20_m_axi_gmem_RDATA;
	input [1:0] sum_20_m_axi_gmem_RRESP;
	input sum_20_m_axi_gmem_RLAST;
	input sum_20_m_axi_gmem_RUSER;
	input sum_20_m_axi_gmem_AWREADY;
	output wire sum_20_m_axi_gmem_AWVALID;
	output wire sum_20_m_axi_gmem_AWID;
	output wire [63:0] sum_20_m_axi_gmem_AWADDR;
	output wire [7:0] sum_20_m_axi_gmem_AWLEN;
	output wire [2:0] sum_20_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_20_m_axi_gmem_AWBURST;
	output wire sum_20_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_20_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_20_m_axi_gmem_AWPROT;
	output wire [3:0] sum_20_m_axi_gmem_AWQOS;
	output wire [3:0] sum_20_m_axi_gmem_AWREGION;
	output wire sum_20_m_axi_gmem_AWUSER;
	input sum_20_m_axi_gmem_WREADY;
	output wire sum_20_m_axi_gmem_WVALID;
	output wire [31:0] sum_20_m_axi_gmem_WDATA;
	output wire [3:0] sum_20_m_axi_gmem_WSTRB;
	output wire sum_20_m_axi_gmem_WLAST;
	output wire sum_20_m_axi_gmem_WUSER;
	output wire sum_20_m_axi_gmem_BREADY;
	input sum_20_m_axi_gmem_BVALID;
	input sum_20_m_axi_gmem_BID;
	input [1:0] sum_20_m_axi_gmem_BRESP;
	input sum_20_m_axi_gmem_BUSER;
	output wire sum_20_s_axi_control_ARREADY;
	input sum_20_s_axi_control_ARVALID;
	input [4:0] sum_20_s_axi_control_ARADDR;
	input sum_20_s_axi_control_RREADY;
	output wire sum_20_s_axi_control_RVALID;
	output wire [31:0] sum_20_s_axi_control_RDATA;
	output wire [1:0] sum_20_s_axi_control_RRESP;
	output wire sum_20_s_axi_control_AWREADY;
	input sum_20_s_axi_control_AWVALID;
	input [4:0] sum_20_s_axi_control_AWADDR;
	output wire sum_20_s_axi_control_WREADY;
	input sum_20_s_axi_control_WVALID;
	input [31:0] sum_20_s_axi_control_WDATA;
	input [3:0] sum_20_s_axi_control_WSTRB;
	input sum_20_s_axi_control_BREADY;
	output wire sum_20_s_axi_control_BVALID;
	output wire [1:0] sum_20_s_axi_control_BRESP;
	input sum_21_m_axi_gmem_ARREADY;
	output wire sum_21_m_axi_gmem_ARVALID;
	output wire sum_21_m_axi_gmem_ARID;
	output wire [63:0] sum_21_m_axi_gmem_ARADDR;
	output wire [7:0] sum_21_m_axi_gmem_ARLEN;
	output wire [2:0] sum_21_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_21_m_axi_gmem_ARBURST;
	output wire sum_21_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_21_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_21_m_axi_gmem_ARPROT;
	output wire [3:0] sum_21_m_axi_gmem_ARQOS;
	output wire [3:0] sum_21_m_axi_gmem_ARREGION;
	output wire sum_21_m_axi_gmem_ARUSER;
	output wire sum_21_m_axi_gmem_RREADY;
	input sum_21_m_axi_gmem_RVALID;
	input sum_21_m_axi_gmem_RID;
	input [31:0] sum_21_m_axi_gmem_RDATA;
	input [1:0] sum_21_m_axi_gmem_RRESP;
	input sum_21_m_axi_gmem_RLAST;
	input sum_21_m_axi_gmem_RUSER;
	input sum_21_m_axi_gmem_AWREADY;
	output wire sum_21_m_axi_gmem_AWVALID;
	output wire sum_21_m_axi_gmem_AWID;
	output wire [63:0] sum_21_m_axi_gmem_AWADDR;
	output wire [7:0] sum_21_m_axi_gmem_AWLEN;
	output wire [2:0] sum_21_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_21_m_axi_gmem_AWBURST;
	output wire sum_21_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_21_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_21_m_axi_gmem_AWPROT;
	output wire [3:0] sum_21_m_axi_gmem_AWQOS;
	output wire [3:0] sum_21_m_axi_gmem_AWREGION;
	output wire sum_21_m_axi_gmem_AWUSER;
	input sum_21_m_axi_gmem_WREADY;
	output wire sum_21_m_axi_gmem_WVALID;
	output wire [31:0] sum_21_m_axi_gmem_WDATA;
	output wire [3:0] sum_21_m_axi_gmem_WSTRB;
	output wire sum_21_m_axi_gmem_WLAST;
	output wire sum_21_m_axi_gmem_WUSER;
	output wire sum_21_m_axi_gmem_BREADY;
	input sum_21_m_axi_gmem_BVALID;
	input sum_21_m_axi_gmem_BID;
	input [1:0] sum_21_m_axi_gmem_BRESP;
	input sum_21_m_axi_gmem_BUSER;
	output wire sum_21_s_axi_control_ARREADY;
	input sum_21_s_axi_control_ARVALID;
	input [4:0] sum_21_s_axi_control_ARADDR;
	input sum_21_s_axi_control_RREADY;
	output wire sum_21_s_axi_control_RVALID;
	output wire [31:0] sum_21_s_axi_control_RDATA;
	output wire [1:0] sum_21_s_axi_control_RRESP;
	output wire sum_21_s_axi_control_AWREADY;
	input sum_21_s_axi_control_AWVALID;
	input [4:0] sum_21_s_axi_control_AWADDR;
	output wire sum_21_s_axi_control_WREADY;
	input sum_21_s_axi_control_WVALID;
	input [31:0] sum_21_s_axi_control_WDATA;
	input [3:0] sum_21_s_axi_control_WSTRB;
	input sum_21_s_axi_control_BREADY;
	output wire sum_21_s_axi_control_BVALID;
	output wire [1:0] sum_21_s_axi_control_BRESP;
	input sum_22_m_axi_gmem_ARREADY;
	output wire sum_22_m_axi_gmem_ARVALID;
	output wire sum_22_m_axi_gmem_ARID;
	output wire [63:0] sum_22_m_axi_gmem_ARADDR;
	output wire [7:0] sum_22_m_axi_gmem_ARLEN;
	output wire [2:0] sum_22_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_22_m_axi_gmem_ARBURST;
	output wire sum_22_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_22_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_22_m_axi_gmem_ARPROT;
	output wire [3:0] sum_22_m_axi_gmem_ARQOS;
	output wire [3:0] sum_22_m_axi_gmem_ARREGION;
	output wire sum_22_m_axi_gmem_ARUSER;
	output wire sum_22_m_axi_gmem_RREADY;
	input sum_22_m_axi_gmem_RVALID;
	input sum_22_m_axi_gmem_RID;
	input [31:0] sum_22_m_axi_gmem_RDATA;
	input [1:0] sum_22_m_axi_gmem_RRESP;
	input sum_22_m_axi_gmem_RLAST;
	input sum_22_m_axi_gmem_RUSER;
	input sum_22_m_axi_gmem_AWREADY;
	output wire sum_22_m_axi_gmem_AWVALID;
	output wire sum_22_m_axi_gmem_AWID;
	output wire [63:0] sum_22_m_axi_gmem_AWADDR;
	output wire [7:0] sum_22_m_axi_gmem_AWLEN;
	output wire [2:0] sum_22_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_22_m_axi_gmem_AWBURST;
	output wire sum_22_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_22_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_22_m_axi_gmem_AWPROT;
	output wire [3:0] sum_22_m_axi_gmem_AWQOS;
	output wire [3:0] sum_22_m_axi_gmem_AWREGION;
	output wire sum_22_m_axi_gmem_AWUSER;
	input sum_22_m_axi_gmem_WREADY;
	output wire sum_22_m_axi_gmem_WVALID;
	output wire [31:0] sum_22_m_axi_gmem_WDATA;
	output wire [3:0] sum_22_m_axi_gmem_WSTRB;
	output wire sum_22_m_axi_gmem_WLAST;
	output wire sum_22_m_axi_gmem_WUSER;
	output wire sum_22_m_axi_gmem_BREADY;
	input sum_22_m_axi_gmem_BVALID;
	input sum_22_m_axi_gmem_BID;
	input [1:0] sum_22_m_axi_gmem_BRESP;
	input sum_22_m_axi_gmem_BUSER;
	output wire sum_22_s_axi_control_ARREADY;
	input sum_22_s_axi_control_ARVALID;
	input [4:0] sum_22_s_axi_control_ARADDR;
	input sum_22_s_axi_control_RREADY;
	output wire sum_22_s_axi_control_RVALID;
	output wire [31:0] sum_22_s_axi_control_RDATA;
	output wire [1:0] sum_22_s_axi_control_RRESP;
	output wire sum_22_s_axi_control_AWREADY;
	input sum_22_s_axi_control_AWVALID;
	input [4:0] sum_22_s_axi_control_AWADDR;
	output wire sum_22_s_axi_control_WREADY;
	input sum_22_s_axi_control_WVALID;
	input [31:0] sum_22_s_axi_control_WDATA;
	input [3:0] sum_22_s_axi_control_WSTRB;
	input sum_22_s_axi_control_BREADY;
	output wire sum_22_s_axi_control_BVALID;
	output wire [1:0] sum_22_s_axi_control_BRESP;
	input sum_23_m_axi_gmem_ARREADY;
	output wire sum_23_m_axi_gmem_ARVALID;
	output wire sum_23_m_axi_gmem_ARID;
	output wire [63:0] sum_23_m_axi_gmem_ARADDR;
	output wire [7:0] sum_23_m_axi_gmem_ARLEN;
	output wire [2:0] sum_23_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_23_m_axi_gmem_ARBURST;
	output wire sum_23_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_23_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_23_m_axi_gmem_ARPROT;
	output wire [3:0] sum_23_m_axi_gmem_ARQOS;
	output wire [3:0] sum_23_m_axi_gmem_ARREGION;
	output wire sum_23_m_axi_gmem_ARUSER;
	output wire sum_23_m_axi_gmem_RREADY;
	input sum_23_m_axi_gmem_RVALID;
	input sum_23_m_axi_gmem_RID;
	input [31:0] sum_23_m_axi_gmem_RDATA;
	input [1:0] sum_23_m_axi_gmem_RRESP;
	input sum_23_m_axi_gmem_RLAST;
	input sum_23_m_axi_gmem_RUSER;
	input sum_23_m_axi_gmem_AWREADY;
	output wire sum_23_m_axi_gmem_AWVALID;
	output wire sum_23_m_axi_gmem_AWID;
	output wire [63:0] sum_23_m_axi_gmem_AWADDR;
	output wire [7:0] sum_23_m_axi_gmem_AWLEN;
	output wire [2:0] sum_23_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_23_m_axi_gmem_AWBURST;
	output wire sum_23_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_23_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_23_m_axi_gmem_AWPROT;
	output wire [3:0] sum_23_m_axi_gmem_AWQOS;
	output wire [3:0] sum_23_m_axi_gmem_AWREGION;
	output wire sum_23_m_axi_gmem_AWUSER;
	input sum_23_m_axi_gmem_WREADY;
	output wire sum_23_m_axi_gmem_WVALID;
	output wire [31:0] sum_23_m_axi_gmem_WDATA;
	output wire [3:0] sum_23_m_axi_gmem_WSTRB;
	output wire sum_23_m_axi_gmem_WLAST;
	output wire sum_23_m_axi_gmem_WUSER;
	output wire sum_23_m_axi_gmem_BREADY;
	input sum_23_m_axi_gmem_BVALID;
	input sum_23_m_axi_gmem_BID;
	input [1:0] sum_23_m_axi_gmem_BRESP;
	input sum_23_m_axi_gmem_BUSER;
	output wire sum_23_s_axi_control_ARREADY;
	input sum_23_s_axi_control_ARVALID;
	input [4:0] sum_23_s_axi_control_ARADDR;
	input sum_23_s_axi_control_RREADY;
	output wire sum_23_s_axi_control_RVALID;
	output wire [31:0] sum_23_s_axi_control_RDATA;
	output wire [1:0] sum_23_s_axi_control_RRESP;
	output wire sum_23_s_axi_control_AWREADY;
	input sum_23_s_axi_control_AWVALID;
	input [4:0] sum_23_s_axi_control_AWADDR;
	output wire sum_23_s_axi_control_WREADY;
	input sum_23_s_axi_control_WVALID;
	input [31:0] sum_23_s_axi_control_WDATA;
	input [3:0] sum_23_s_axi_control_WSTRB;
	input sum_23_s_axi_control_BREADY;
	output wire sum_23_s_axi_control_BVALID;
	output wire [1:0] sum_23_s_axi_control_BRESP;
	input sum_24_m_axi_gmem_ARREADY;
	output wire sum_24_m_axi_gmem_ARVALID;
	output wire sum_24_m_axi_gmem_ARID;
	output wire [63:0] sum_24_m_axi_gmem_ARADDR;
	output wire [7:0] sum_24_m_axi_gmem_ARLEN;
	output wire [2:0] sum_24_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_24_m_axi_gmem_ARBURST;
	output wire sum_24_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_24_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_24_m_axi_gmem_ARPROT;
	output wire [3:0] sum_24_m_axi_gmem_ARQOS;
	output wire [3:0] sum_24_m_axi_gmem_ARREGION;
	output wire sum_24_m_axi_gmem_ARUSER;
	output wire sum_24_m_axi_gmem_RREADY;
	input sum_24_m_axi_gmem_RVALID;
	input sum_24_m_axi_gmem_RID;
	input [31:0] sum_24_m_axi_gmem_RDATA;
	input [1:0] sum_24_m_axi_gmem_RRESP;
	input sum_24_m_axi_gmem_RLAST;
	input sum_24_m_axi_gmem_RUSER;
	input sum_24_m_axi_gmem_AWREADY;
	output wire sum_24_m_axi_gmem_AWVALID;
	output wire sum_24_m_axi_gmem_AWID;
	output wire [63:0] sum_24_m_axi_gmem_AWADDR;
	output wire [7:0] sum_24_m_axi_gmem_AWLEN;
	output wire [2:0] sum_24_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_24_m_axi_gmem_AWBURST;
	output wire sum_24_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_24_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_24_m_axi_gmem_AWPROT;
	output wire [3:0] sum_24_m_axi_gmem_AWQOS;
	output wire [3:0] sum_24_m_axi_gmem_AWREGION;
	output wire sum_24_m_axi_gmem_AWUSER;
	input sum_24_m_axi_gmem_WREADY;
	output wire sum_24_m_axi_gmem_WVALID;
	output wire [31:0] sum_24_m_axi_gmem_WDATA;
	output wire [3:0] sum_24_m_axi_gmem_WSTRB;
	output wire sum_24_m_axi_gmem_WLAST;
	output wire sum_24_m_axi_gmem_WUSER;
	output wire sum_24_m_axi_gmem_BREADY;
	input sum_24_m_axi_gmem_BVALID;
	input sum_24_m_axi_gmem_BID;
	input [1:0] sum_24_m_axi_gmem_BRESP;
	input sum_24_m_axi_gmem_BUSER;
	output wire sum_24_s_axi_control_ARREADY;
	input sum_24_s_axi_control_ARVALID;
	input [4:0] sum_24_s_axi_control_ARADDR;
	input sum_24_s_axi_control_RREADY;
	output wire sum_24_s_axi_control_RVALID;
	output wire [31:0] sum_24_s_axi_control_RDATA;
	output wire [1:0] sum_24_s_axi_control_RRESP;
	output wire sum_24_s_axi_control_AWREADY;
	input sum_24_s_axi_control_AWVALID;
	input [4:0] sum_24_s_axi_control_AWADDR;
	output wire sum_24_s_axi_control_WREADY;
	input sum_24_s_axi_control_WVALID;
	input [31:0] sum_24_s_axi_control_WDATA;
	input [3:0] sum_24_s_axi_control_WSTRB;
	input sum_24_s_axi_control_BREADY;
	output wire sum_24_s_axi_control_BVALID;
	output wire [1:0] sum_24_s_axi_control_BRESP;
	input sum_25_m_axi_gmem_ARREADY;
	output wire sum_25_m_axi_gmem_ARVALID;
	output wire sum_25_m_axi_gmem_ARID;
	output wire [63:0] sum_25_m_axi_gmem_ARADDR;
	output wire [7:0] sum_25_m_axi_gmem_ARLEN;
	output wire [2:0] sum_25_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_25_m_axi_gmem_ARBURST;
	output wire sum_25_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_25_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_25_m_axi_gmem_ARPROT;
	output wire [3:0] sum_25_m_axi_gmem_ARQOS;
	output wire [3:0] sum_25_m_axi_gmem_ARREGION;
	output wire sum_25_m_axi_gmem_ARUSER;
	output wire sum_25_m_axi_gmem_RREADY;
	input sum_25_m_axi_gmem_RVALID;
	input sum_25_m_axi_gmem_RID;
	input [31:0] sum_25_m_axi_gmem_RDATA;
	input [1:0] sum_25_m_axi_gmem_RRESP;
	input sum_25_m_axi_gmem_RLAST;
	input sum_25_m_axi_gmem_RUSER;
	input sum_25_m_axi_gmem_AWREADY;
	output wire sum_25_m_axi_gmem_AWVALID;
	output wire sum_25_m_axi_gmem_AWID;
	output wire [63:0] sum_25_m_axi_gmem_AWADDR;
	output wire [7:0] sum_25_m_axi_gmem_AWLEN;
	output wire [2:0] sum_25_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_25_m_axi_gmem_AWBURST;
	output wire sum_25_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_25_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_25_m_axi_gmem_AWPROT;
	output wire [3:0] sum_25_m_axi_gmem_AWQOS;
	output wire [3:0] sum_25_m_axi_gmem_AWREGION;
	output wire sum_25_m_axi_gmem_AWUSER;
	input sum_25_m_axi_gmem_WREADY;
	output wire sum_25_m_axi_gmem_WVALID;
	output wire [31:0] sum_25_m_axi_gmem_WDATA;
	output wire [3:0] sum_25_m_axi_gmem_WSTRB;
	output wire sum_25_m_axi_gmem_WLAST;
	output wire sum_25_m_axi_gmem_WUSER;
	output wire sum_25_m_axi_gmem_BREADY;
	input sum_25_m_axi_gmem_BVALID;
	input sum_25_m_axi_gmem_BID;
	input [1:0] sum_25_m_axi_gmem_BRESP;
	input sum_25_m_axi_gmem_BUSER;
	output wire sum_25_s_axi_control_ARREADY;
	input sum_25_s_axi_control_ARVALID;
	input [4:0] sum_25_s_axi_control_ARADDR;
	input sum_25_s_axi_control_RREADY;
	output wire sum_25_s_axi_control_RVALID;
	output wire [31:0] sum_25_s_axi_control_RDATA;
	output wire [1:0] sum_25_s_axi_control_RRESP;
	output wire sum_25_s_axi_control_AWREADY;
	input sum_25_s_axi_control_AWVALID;
	input [4:0] sum_25_s_axi_control_AWADDR;
	output wire sum_25_s_axi_control_WREADY;
	input sum_25_s_axi_control_WVALID;
	input [31:0] sum_25_s_axi_control_WDATA;
	input [3:0] sum_25_s_axi_control_WSTRB;
	input sum_25_s_axi_control_BREADY;
	output wire sum_25_s_axi_control_BVALID;
	output wire [1:0] sum_25_s_axi_control_BRESP;
	input sum_26_m_axi_gmem_ARREADY;
	output wire sum_26_m_axi_gmem_ARVALID;
	output wire sum_26_m_axi_gmem_ARID;
	output wire [63:0] sum_26_m_axi_gmem_ARADDR;
	output wire [7:0] sum_26_m_axi_gmem_ARLEN;
	output wire [2:0] sum_26_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_26_m_axi_gmem_ARBURST;
	output wire sum_26_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_26_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_26_m_axi_gmem_ARPROT;
	output wire [3:0] sum_26_m_axi_gmem_ARQOS;
	output wire [3:0] sum_26_m_axi_gmem_ARREGION;
	output wire sum_26_m_axi_gmem_ARUSER;
	output wire sum_26_m_axi_gmem_RREADY;
	input sum_26_m_axi_gmem_RVALID;
	input sum_26_m_axi_gmem_RID;
	input [31:0] sum_26_m_axi_gmem_RDATA;
	input [1:0] sum_26_m_axi_gmem_RRESP;
	input sum_26_m_axi_gmem_RLAST;
	input sum_26_m_axi_gmem_RUSER;
	input sum_26_m_axi_gmem_AWREADY;
	output wire sum_26_m_axi_gmem_AWVALID;
	output wire sum_26_m_axi_gmem_AWID;
	output wire [63:0] sum_26_m_axi_gmem_AWADDR;
	output wire [7:0] sum_26_m_axi_gmem_AWLEN;
	output wire [2:0] sum_26_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_26_m_axi_gmem_AWBURST;
	output wire sum_26_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_26_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_26_m_axi_gmem_AWPROT;
	output wire [3:0] sum_26_m_axi_gmem_AWQOS;
	output wire [3:0] sum_26_m_axi_gmem_AWREGION;
	output wire sum_26_m_axi_gmem_AWUSER;
	input sum_26_m_axi_gmem_WREADY;
	output wire sum_26_m_axi_gmem_WVALID;
	output wire [31:0] sum_26_m_axi_gmem_WDATA;
	output wire [3:0] sum_26_m_axi_gmem_WSTRB;
	output wire sum_26_m_axi_gmem_WLAST;
	output wire sum_26_m_axi_gmem_WUSER;
	output wire sum_26_m_axi_gmem_BREADY;
	input sum_26_m_axi_gmem_BVALID;
	input sum_26_m_axi_gmem_BID;
	input [1:0] sum_26_m_axi_gmem_BRESP;
	input sum_26_m_axi_gmem_BUSER;
	output wire sum_26_s_axi_control_ARREADY;
	input sum_26_s_axi_control_ARVALID;
	input [4:0] sum_26_s_axi_control_ARADDR;
	input sum_26_s_axi_control_RREADY;
	output wire sum_26_s_axi_control_RVALID;
	output wire [31:0] sum_26_s_axi_control_RDATA;
	output wire [1:0] sum_26_s_axi_control_RRESP;
	output wire sum_26_s_axi_control_AWREADY;
	input sum_26_s_axi_control_AWVALID;
	input [4:0] sum_26_s_axi_control_AWADDR;
	output wire sum_26_s_axi_control_WREADY;
	input sum_26_s_axi_control_WVALID;
	input [31:0] sum_26_s_axi_control_WDATA;
	input [3:0] sum_26_s_axi_control_WSTRB;
	input sum_26_s_axi_control_BREADY;
	output wire sum_26_s_axi_control_BVALID;
	output wire [1:0] sum_26_s_axi_control_BRESP;
	input sum_27_m_axi_gmem_ARREADY;
	output wire sum_27_m_axi_gmem_ARVALID;
	output wire sum_27_m_axi_gmem_ARID;
	output wire [63:0] sum_27_m_axi_gmem_ARADDR;
	output wire [7:0] sum_27_m_axi_gmem_ARLEN;
	output wire [2:0] sum_27_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_27_m_axi_gmem_ARBURST;
	output wire sum_27_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_27_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_27_m_axi_gmem_ARPROT;
	output wire [3:0] sum_27_m_axi_gmem_ARQOS;
	output wire [3:0] sum_27_m_axi_gmem_ARREGION;
	output wire sum_27_m_axi_gmem_ARUSER;
	output wire sum_27_m_axi_gmem_RREADY;
	input sum_27_m_axi_gmem_RVALID;
	input sum_27_m_axi_gmem_RID;
	input [31:0] sum_27_m_axi_gmem_RDATA;
	input [1:0] sum_27_m_axi_gmem_RRESP;
	input sum_27_m_axi_gmem_RLAST;
	input sum_27_m_axi_gmem_RUSER;
	input sum_27_m_axi_gmem_AWREADY;
	output wire sum_27_m_axi_gmem_AWVALID;
	output wire sum_27_m_axi_gmem_AWID;
	output wire [63:0] sum_27_m_axi_gmem_AWADDR;
	output wire [7:0] sum_27_m_axi_gmem_AWLEN;
	output wire [2:0] sum_27_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_27_m_axi_gmem_AWBURST;
	output wire sum_27_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_27_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_27_m_axi_gmem_AWPROT;
	output wire [3:0] sum_27_m_axi_gmem_AWQOS;
	output wire [3:0] sum_27_m_axi_gmem_AWREGION;
	output wire sum_27_m_axi_gmem_AWUSER;
	input sum_27_m_axi_gmem_WREADY;
	output wire sum_27_m_axi_gmem_WVALID;
	output wire [31:0] sum_27_m_axi_gmem_WDATA;
	output wire [3:0] sum_27_m_axi_gmem_WSTRB;
	output wire sum_27_m_axi_gmem_WLAST;
	output wire sum_27_m_axi_gmem_WUSER;
	output wire sum_27_m_axi_gmem_BREADY;
	input sum_27_m_axi_gmem_BVALID;
	input sum_27_m_axi_gmem_BID;
	input [1:0] sum_27_m_axi_gmem_BRESP;
	input sum_27_m_axi_gmem_BUSER;
	output wire sum_27_s_axi_control_ARREADY;
	input sum_27_s_axi_control_ARVALID;
	input [4:0] sum_27_s_axi_control_ARADDR;
	input sum_27_s_axi_control_RREADY;
	output wire sum_27_s_axi_control_RVALID;
	output wire [31:0] sum_27_s_axi_control_RDATA;
	output wire [1:0] sum_27_s_axi_control_RRESP;
	output wire sum_27_s_axi_control_AWREADY;
	input sum_27_s_axi_control_AWVALID;
	input [4:0] sum_27_s_axi_control_AWADDR;
	output wire sum_27_s_axi_control_WREADY;
	input sum_27_s_axi_control_WVALID;
	input [31:0] sum_27_s_axi_control_WDATA;
	input [3:0] sum_27_s_axi_control_WSTRB;
	input sum_27_s_axi_control_BREADY;
	output wire sum_27_s_axi_control_BVALID;
	output wire [1:0] sum_27_s_axi_control_BRESP;
	input sum_28_m_axi_gmem_ARREADY;
	output wire sum_28_m_axi_gmem_ARVALID;
	output wire sum_28_m_axi_gmem_ARID;
	output wire [63:0] sum_28_m_axi_gmem_ARADDR;
	output wire [7:0] sum_28_m_axi_gmem_ARLEN;
	output wire [2:0] sum_28_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_28_m_axi_gmem_ARBURST;
	output wire sum_28_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_28_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_28_m_axi_gmem_ARPROT;
	output wire [3:0] sum_28_m_axi_gmem_ARQOS;
	output wire [3:0] sum_28_m_axi_gmem_ARREGION;
	output wire sum_28_m_axi_gmem_ARUSER;
	output wire sum_28_m_axi_gmem_RREADY;
	input sum_28_m_axi_gmem_RVALID;
	input sum_28_m_axi_gmem_RID;
	input [31:0] sum_28_m_axi_gmem_RDATA;
	input [1:0] sum_28_m_axi_gmem_RRESP;
	input sum_28_m_axi_gmem_RLAST;
	input sum_28_m_axi_gmem_RUSER;
	input sum_28_m_axi_gmem_AWREADY;
	output wire sum_28_m_axi_gmem_AWVALID;
	output wire sum_28_m_axi_gmem_AWID;
	output wire [63:0] sum_28_m_axi_gmem_AWADDR;
	output wire [7:0] sum_28_m_axi_gmem_AWLEN;
	output wire [2:0] sum_28_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_28_m_axi_gmem_AWBURST;
	output wire sum_28_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_28_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_28_m_axi_gmem_AWPROT;
	output wire [3:0] sum_28_m_axi_gmem_AWQOS;
	output wire [3:0] sum_28_m_axi_gmem_AWREGION;
	output wire sum_28_m_axi_gmem_AWUSER;
	input sum_28_m_axi_gmem_WREADY;
	output wire sum_28_m_axi_gmem_WVALID;
	output wire [31:0] sum_28_m_axi_gmem_WDATA;
	output wire [3:0] sum_28_m_axi_gmem_WSTRB;
	output wire sum_28_m_axi_gmem_WLAST;
	output wire sum_28_m_axi_gmem_WUSER;
	output wire sum_28_m_axi_gmem_BREADY;
	input sum_28_m_axi_gmem_BVALID;
	input sum_28_m_axi_gmem_BID;
	input [1:0] sum_28_m_axi_gmem_BRESP;
	input sum_28_m_axi_gmem_BUSER;
	output wire sum_28_s_axi_control_ARREADY;
	input sum_28_s_axi_control_ARVALID;
	input [4:0] sum_28_s_axi_control_ARADDR;
	input sum_28_s_axi_control_RREADY;
	output wire sum_28_s_axi_control_RVALID;
	output wire [31:0] sum_28_s_axi_control_RDATA;
	output wire [1:0] sum_28_s_axi_control_RRESP;
	output wire sum_28_s_axi_control_AWREADY;
	input sum_28_s_axi_control_AWVALID;
	input [4:0] sum_28_s_axi_control_AWADDR;
	output wire sum_28_s_axi_control_WREADY;
	input sum_28_s_axi_control_WVALID;
	input [31:0] sum_28_s_axi_control_WDATA;
	input [3:0] sum_28_s_axi_control_WSTRB;
	input sum_28_s_axi_control_BREADY;
	output wire sum_28_s_axi_control_BVALID;
	output wire [1:0] sum_28_s_axi_control_BRESP;
	input sum_29_m_axi_gmem_ARREADY;
	output wire sum_29_m_axi_gmem_ARVALID;
	output wire sum_29_m_axi_gmem_ARID;
	output wire [63:0] sum_29_m_axi_gmem_ARADDR;
	output wire [7:0] sum_29_m_axi_gmem_ARLEN;
	output wire [2:0] sum_29_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_29_m_axi_gmem_ARBURST;
	output wire sum_29_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_29_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_29_m_axi_gmem_ARPROT;
	output wire [3:0] sum_29_m_axi_gmem_ARQOS;
	output wire [3:0] sum_29_m_axi_gmem_ARREGION;
	output wire sum_29_m_axi_gmem_ARUSER;
	output wire sum_29_m_axi_gmem_RREADY;
	input sum_29_m_axi_gmem_RVALID;
	input sum_29_m_axi_gmem_RID;
	input [31:0] sum_29_m_axi_gmem_RDATA;
	input [1:0] sum_29_m_axi_gmem_RRESP;
	input sum_29_m_axi_gmem_RLAST;
	input sum_29_m_axi_gmem_RUSER;
	input sum_29_m_axi_gmem_AWREADY;
	output wire sum_29_m_axi_gmem_AWVALID;
	output wire sum_29_m_axi_gmem_AWID;
	output wire [63:0] sum_29_m_axi_gmem_AWADDR;
	output wire [7:0] sum_29_m_axi_gmem_AWLEN;
	output wire [2:0] sum_29_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_29_m_axi_gmem_AWBURST;
	output wire sum_29_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_29_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_29_m_axi_gmem_AWPROT;
	output wire [3:0] sum_29_m_axi_gmem_AWQOS;
	output wire [3:0] sum_29_m_axi_gmem_AWREGION;
	output wire sum_29_m_axi_gmem_AWUSER;
	input sum_29_m_axi_gmem_WREADY;
	output wire sum_29_m_axi_gmem_WVALID;
	output wire [31:0] sum_29_m_axi_gmem_WDATA;
	output wire [3:0] sum_29_m_axi_gmem_WSTRB;
	output wire sum_29_m_axi_gmem_WLAST;
	output wire sum_29_m_axi_gmem_WUSER;
	output wire sum_29_m_axi_gmem_BREADY;
	input sum_29_m_axi_gmem_BVALID;
	input sum_29_m_axi_gmem_BID;
	input [1:0] sum_29_m_axi_gmem_BRESP;
	input sum_29_m_axi_gmem_BUSER;
	output wire sum_29_s_axi_control_ARREADY;
	input sum_29_s_axi_control_ARVALID;
	input [4:0] sum_29_s_axi_control_ARADDR;
	input sum_29_s_axi_control_RREADY;
	output wire sum_29_s_axi_control_RVALID;
	output wire [31:0] sum_29_s_axi_control_RDATA;
	output wire [1:0] sum_29_s_axi_control_RRESP;
	output wire sum_29_s_axi_control_AWREADY;
	input sum_29_s_axi_control_AWVALID;
	input [4:0] sum_29_s_axi_control_AWADDR;
	output wire sum_29_s_axi_control_WREADY;
	input sum_29_s_axi_control_WVALID;
	input [31:0] sum_29_s_axi_control_WDATA;
	input [3:0] sum_29_s_axi_control_WSTRB;
	input sum_29_s_axi_control_BREADY;
	output wire sum_29_s_axi_control_BVALID;
	output wire [1:0] sum_29_s_axi_control_BRESP;
	input sum_30_m_axi_gmem_ARREADY;
	output wire sum_30_m_axi_gmem_ARVALID;
	output wire sum_30_m_axi_gmem_ARID;
	output wire [63:0] sum_30_m_axi_gmem_ARADDR;
	output wire [7:0] sum_30_m_axi_gmem_ARLEN;
	output wire [2:0] sum_30_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_30_m_axi_gmem_ARBURST;
	output wire sum_30_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_30_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_30_m_axi_gmem_ARPROT;
	output wire [3:0] sum_30_m_axi_gmem_ARQOS;
	output wire [3:0] sum_30_m_axi_gmem_ARREGION;
	output wire sum_30_m_axi_gmem_ARUSER;
	output wire sum_30_m_axi_gmem_RREADY;
	input sum_30_m_axi_gmem_RVALID;
	input sum_30_m_axi_gmem_RID;
	input [31:0] sum_30_m_axi_gmem_RDATA;
	input [1:0] sum_30_m_axi_gmem_RRESP;
	input sum_30_m_axi_gmem_RLAST;
	input sum_30_m_axi_gmem_RUSER;
	input sum_30_m_axi_gmem_AWREADY;
	output wire sum_30_m_axi_gmem_AWVALID;
	output wire sum_30_m_axi_gmem_AWID;
	output wire [63:0] sum_30_m_axi_gmem_AWADDR;
	output wire [7:0] sum_30_m_axi_gmem_AWLEN;
	output wire [2:0] sum_30_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_30_m_axi_gmem_AWBURST;
	output wire sum_30_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_30_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_30_m_axi_gmem_AWPROT;
	output wire [3:0] sum_30_m_axi_gmem_AWQOS;
	output wire [3:0] sum_30_m_axi_gmem_AWREGION;
	output wire sum_30_m_axi_gmem_AWUSER;
	input sum_30_m_axi_gmem_WREADY;
	output wire sum_30_m_axi_gmem_WVALID;
	output wire [31:0] sum_30_m_axi_gmem_WDATA;
	output wire [3:0] sum_30_m_axi_gmem_WSTRB;
	output wire sum_30_m_axi_gmem_WLAST;
	output wire sum_30_m_axi_gmem_WUSER;
	output wire sum_30_m_axi_gmem_BREADY;
	input sum_30_m_axi_gmem_BVALID;
	input sum_30_m_axi_gmem_BID;
	input [1:0] sum_30_m_axi_gmem_BRESP;
	input sum_30_m_axi_gmem_BUSER;
	output wire sum_30_s_axi_control_ARREADY;
	input sum_30_s_axi_control_ARVALID;
	input [4:0] sum_30_s_axi_control_ARADDR;
	input sum_30_s_axi_control_RREADY;
	output wire sum_30_s_axi_control_RVALID;
	output wire [31:0] sum_30_s_axi_control_RDATA;
	output wire [1:0] sum_30_s_axi_control_RRESP;
	output wire sum_30_s_axi_control_AWREADY;
	input sum_30_s_axi_control_AWVALID;
	input [4:0] sum_30_s_axi_control_AWADDR;
	output wire sum_30_s_axi_control_WREADY;
	input sum_30_s_axi_control_WVALID;
	input [31:0] sum_30_s_axi_control_WDATA;
	input [3:0] sum_30_s_axi_control_WSTRB;
	input sum_30_s_axi_control_BREADY;
	output wire sum_30_s_axi_control_BVALID;
	output wire [1:0] sum_30_s_axi_control_BRESP;
	input sum_31_m_axi_gmem_ARREADY;
	output wire sum_31_m_axi_gmem_ARVALID;
	output wire sum_31_m_axi_gmem_ARID;
	output wire [63:0] sum_31_m_axi_gmem_ARADDR;
	output wire [7:0] sum_31_m_axi_gmem_ARLEN;
	output wire [2:0] sum_31_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_31_m_axi_gmem_ARBURST;
	output wire sum_31_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_31_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_31_m_axi_gmem_ARPROT;
	output wire [3:0] sum_31_m_axi_gmem_ARQOS;
	output wire [3:0] sum_31_m_axi_gmem_ARREGION;
	output wire sum_31_m_axi_gmem_ARUSER;
	output wire sum_31_m_axi_gmem_RREADY;
	input sum_31_m_axi_gmem_RVALID;
	input sum_31_m_axi_gmem_RID;
	input [31:0] sum_31_m_axi_gmem_RDATA;
	input [1:0] sum_31_m_axi_gmem_RRESP;
	input sum_31_m_axi_gmem_RLAST;
	input sum_31_m_axi_gmem_RUSER;
	input sum_31_m_axi_gmem_AWREADY;
	output wire sum_31_m_axi_gmem_AWVALID;
	output wire sum_31_m_axi_gmem_AWID;
	output wire [63:0] sum_31_m_axi_gmem_AWADDR;
	output wire [7:0] sum_31_m_axi_gmem_AWLEN;
	output wire [2:0] sum_31_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_31_m_axi_gmem_AWBURST;
	output wire sum_31_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_31_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_31_m_axi_gmem_AWPROT;
	output wire [3:0] sum_31_m_axi_gmem_AWQOS;
	output wire [3:0] sum_31_m_axi_gmem_AWREGION;
	output wire sum_31_m_axi_gmem_AWUSER;
	input sum_31_m_axi_gmem_WREADY;
	output wire sum_31_m_axi_gmem_WVALID;
	output wire [31:0] sum_31_m_axi_gmem_WDATA;
	output wire [3:0] sum_31_m_axi_gmem_WSTRB;
	output wire sum_31_m_axi_gmem_WLAST;
	output wire sum_31_m_axi_gmem_WUSER;
	output wire sum_31_m_axi_gmem_BREADY;
	input sum_31_m_axi_gmem_BVALID;
	input sum_31_m_axi_gmem_BID;
	input [1:0] sum_31_m_axi_gmem_BRESP;
	input sum_31_m_axi_gmem_BUSER;
	output wire sum_31_s_axi_control_ARREADY;
	input sum_31_s_axi_control_ARVALID;
	input [4:0] sum_31_s_axi_control_ARADDR;
	input sum_31_s_axi_control_RREADY;
	output wire sum_31_s_axi_control_RVALID;
	output wire [31:0] sum_31_s_axi_control_RDATA;
	output wire [1:0] sum_31_s_axi_control_RRESP;
	output wire sum_31_s_axi_control_AWREADY;
	input sum_31_s_axi_control_AWVALID;
	input [4:0] sum_31_s_axi_control_AWADDR;
	output wire sum_31_s_axi_control_WREADY;
	input sum_31_s_axi_control_WVALID;
	input [31:0] sum_31_s_axi_control_WDATA;
	input [3:0] sum_31_s_axi_control_WSTRB;
	input sum_31_s_axi_control_BREADY;
	output wire sum_31_s_axi_control_BVALID;
	output wire [1:0] sum_31_s_axi_control_BRESP;
	input sum_32_m_axi_gmem_ARREADY;
	output wire sum_32_m_axi_gmem_ARVALID;
	output wire sum_32_m_axi_gmem_ARID;
	output wire [63:0] sum_32_m_axi_gmem_ARADDR;
	output wire [7:0] sum_32_m_axi_gmem_ARLEN;
	output wire [2:0] sum_32_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_32_m_axi_gmem_ARBURST;
	output wire sum_32_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_32_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_32_m_axi_gmem_ARPROT;
	output wire [3:0] sum_32_m_axi_gmem_ARQOS;
	output wire [3:0] sum_32_m_axi_gmem_ARREGION;
	output wire sum_32_m_axi_gmem_ARUSER;
	output wire sum_32_m_axi_gmem_RREADY;
	input sum_32_m_axi_gmem_RVALID;
	input sum_32_m_axi_gmem_RID;
	input [31:0] sum_32_m_axi_gmem_RDATA;
	input [1:0] sum_32_m_axi_gmem_RRESP;
	input sum_32_m_axi_gmem_RLAST;
	input sum_32_m_axi_gmem_RUSER;
	input sum_32_m_axi_gmem_AWREADY;
	output wire sum_32_m_axi_gmem_AWVALID;
	output wire sum_32_m_axi_gmem_AWID;
	output wire [63:0] sum_32_m_axi_gmem_AWADDR;
	output wire [7:0] sum_32_m_axi_gmem_AWLEN;
	output wire [2:0] sum_32_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_32_m_axi_gmem_AWBURST;
	output wire sum_32_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_32_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_32_m_axi_gmem_AWPROT;
	output wire [3:0] sum_32_m_axi_gmem_AWQOS;
	output wire [3:0] sum_32_m_axi_gmem_AWREGION;
	output wire sum_32_m_axi_gmem_AWUSER;
	input sum_32_m_axi_gmem_WREADY;
	output wire sum_32_m_axi_gmem_WVALID;
	output wire [31:0] sum_32_m_axi_gmem_WDATA;
	output wire [3:0] sum_32_m_axi_gmem_WSTRB;
	output wire sum_32_m_axi_gmem_WLAST;
	output wire sum_32_m_axi_gmem_WUSER;
	output wire sum_32_m_axi_gmem_BREADY;
	input sum_32_m_axi_gmem_BVALID;
	input sum_32_m_axi_gmem_BID;
	input [1:0] sum_32_m_axi_gmem_BRESP;
	input sum_32_m_axi_gmem_BUSER;
	output wire sum_32_s_axi_control_ARREADY;
	input sum_32_s_axi_control_ARVALID;
	input [4:0] sum_32_s_axi_control_ARADDR;
	input sum_32_s_axi_control_RREADY;
	output wire sum_32_s_axi_control_RVALID;
	output wire [31:0] sum_32_s_axi_control_RDATA;
	output wire [1:0] sum_32_s_axi_control_RRESP;
	output wire sum_32_s_axi_control_AWREADY;
	input sum_32_s_axi_control_AWVALID;
	input [4:0] sum_32_s_axi_control_AWADDR;
	output wire sum_32_s_axi_control_WREADY;
	input sum_32_s_axi_control_WVALID;
	input [31:0] sum_32_s_axi_control_WDATA;
	input [3:0] sum_32_s_axi_control_WSTRB;
	input sum_32_s_axi_control_BREADY;
	output wire sum_32_s_axi_control_BVALID;
	output wire [1:0] sum_32_s_axi_control_BRESP;
	input sum_33_m_axi_gmem_ARREADY;
	output wire sum_33_m_axi_gmem_ARVALID;
	output wire sum_33_m_axi_gmem_ARID;
	output wire [63:0] sum_33_m_axi_gmem_ARADDR;
	output wire [7:0] sum_33_m_axi_gmem_ARLEN;
	output wire [2:0] sum_33_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_33_m_axi_gmem_ARBURST;
	output wire sum_33_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_33_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_33_m_axi_gmem_ARPROT;
	output wire [3:0] sum_33_m_axi_gmem_ARQOS;
	output wire [3:0] sum_33_m_axi_gmem_ARREGION;
	output wire sum_33_m_axi_gmem_ARUSER;
	output wire sum_33_m_axi_gmem_RREADY;
	input sum_33_m_axi_gmem_RVALID;
	input sum_33_m_axi_gmem_RID;
	input [31:0] sum_33_m_axi_gmem_RDATA;
	input [1:0] sum_33_m_axi_gmem_RRESP;
	input sum_33_m_axi_gmem_RLAST;
	input sum_33_m_axi_gmem_RUSER;
	input sum_33_m_axi_gmem_AWREADY;
	output wire sum_33_m_axi_gmem_AWVALID;
	output wire sum_33_m_axi_gmem_AWID;
	output wire [63:0] sum_33_m_axi_gmem_AWADDR;
	output wire [7:0] sum_33_m_axi_gmem_AWLEN;
	output wire [2:0] sum_33_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_33_m_axi_gmem_AWBURST;
	output wire sum_33_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_33_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_33_m_axi_gmem_AWPROT;
	output wire [3:0] sum_33_m_axi_gmem_AWQOS;
	output wire [3:0] sum_33_m_axi_gmem_AWREGION;
	output wire sum_33_m_axi_gmem_AWUSER;
	input sum_33_m_axi_gmem_WREADY;
	output wire sum_33_m_axi_gmem_WVALID;
	output wire [31:0] sum_33_m_axi_gmem_WDATA;
	output wire [3:0] sum_33_m_axi_gmem_WSTRB;
	output wire sum_33_m_axi_gmem_WLAST;
	output wire sum_33_m_axi_gmem_WUSER;
	output wire sum_33_m_axi_gmem_BREADY;
	input sum_33_m_axi_gmem_BVALID;
	input sum_33_m_axi_gmem_BID;
	input [1:0] sum_33_m_axi_gmem_BRESP;
	input sum_33_m_axi_gmem_BUSER;
	output wire sum_33_s_axi_control_ARREADY;
	input sum_33_s_axi_control_ARVALID;
	input [4:0] sum_33_s_axi_control_ARADDR;
	input sum_33_s_axi_control_RREADY;
	output wire sum_33_s_axi_control_RVALID;
	output wire [31:0] sum_33_s_axi_control_RDATA;
	output wire [1:0] sum_33_s_axi_control_RRESP;
	output wire sum_33_s_axi_control_AWREADY;
	input sum_33_s_axi_control_AWVALID;
	input [4:0] sum_33_s_axi_control_AWADDR;
	output wire sum_33_s_axi_control_WREADY;
	input sum_33_s_axi_control_WVALID;
	input [31:0] sum_33_s_axi_control_WDATA;
	input [3:0] sum_33_s_axi_control_WSTRB;
	input sum_33_s_axi_control_BREADY;
	output wire sum_33_s_axi_control_BVALID;
	output wire [1:0] sum_33_s_axi_control_BRESP;
	input sum_34_m_axi_gmem_ARREADY;
	output wire sum_34_m_axi_gmem_ARVALID;
	output wire sum_34_m_axi_gmem_ARID;
	output wire [63:0] sum_34_m_axi_gmem_ARADDR;
	output wire [7:0] sum_34_m_axi_gmem_ARLEN;
	output wire [2:0] sum_34_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_34_m_axi_gmem_ARBURST;
	output wire sum_34_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_34_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_34_m_axi_gmem_ARPROT;
	output wire [3:0] sum_34_m_axi_gmem_ARQOS;
	output wire [3:0] sum_34_m_axi_gmem_ARREGION;
	output wire sum_34_m_axi_gmem_ARUSER;
	output wire sum_34_m_axi_gmem_RREADY;
	input sum_34_m_axi_gmem_RVALID;
	input sum_34_m_axi_gmem_RID;
	input [31:0] sum_34_m_axi_gmem_RDATA;
	input [1:0] sum_34_m_axi_gmem_RRESP;
	input sum_34_m_axi_gmem_RLAST;
	input sum_34_m_axi_gmem_RUSER;
	input sum_34_m_axi_gmem_AWREADY;
	output wire sum_34_m_axi_gmem_AWVALID;
	output wire sum_34_m_axi_gmem_AWID;
	output wire [63:0] sum_34_m_axi_gmem_AWADDR;
	output wire [7:0] sum_34_m_axi_gmem_AWLEN;
	output wire [2:0] sum_34_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_34_m_axi_gmem_AWBURST;
	output wire sum_34_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_34_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_34_m_axi_gmem_AWPROT;
	output wire [3:0] sum_34_m_axi_gmem_AWQOS;
	output wire [3:0] sum_34_m_axi_gmem_AWREGION;
	output wire sum_34_m_axi_gmem_AWUSER;
	input sum_34_m_axi_gmem_WREADY;
	output wire sum_34_m_axi_gmem_WVALID;
	output wire [31:0] sum_34_m_axi_gmem_WDATA;
	output wire [3:0] sum_34_m_axi_gmem_WSTRB;
	output wire sum_34_m_axi_gmem_WLAST;
	output wire sum_34_m_axi_gmem_WUSER;
	output wire sum_34_m_axi_gmem_BREADY;
	input sum_34_m_axi_gmem_BVALID;
	input sum_34_m_axi_gmem_BID;
	input [1:0] sum_34_m_axi_gmem_BRESP;
	input sum_34_m_axi_gmem_BUSER;
	output wire sum_34_s_axi_control_ARREADY;
	input sum_34_s_axi_control_ARVALID;
	input [4:0] sum_34_s_axi_control_ARADDR;
	input sum_34_s_axi_control_RREADY;
	output wire sum_34_s_axi_control_RVALID;
	output wire [31:0] sum_34_s_axi_control_RDATA;
	output wire [1:0] sum_34_s_axi_control_RRESP;
	output wire sum_34_s_axi_control_AWREADY;
	input sum_34_s_axi_control_AWVALID;
	input [4:0] sum_34_s_axi_control_AWADDR;
	output wire sum_34_s_axi_control_WREADY;
	input sum_34_s_axi_control_WVALID;
	input [31:0] sum_34_s_axi_control_WDATA;
	input [3:0] sum_34_s_axi_control_WSTRB;
	input sum_34_s_axi_control_BREADY;
	output wire sum_34_s_axi_control_BVALID;
	output wire [1:0] sum_34_s_axi_control_BRESP;
	input sum_35_m_axi_gmem_ARREADY;
	output wire sum_35_m_axi_gmem_ARVALID;
	output wire sum_35_m_axi_gmem_ARID;
	output wire [63:0] sum_35_m_axi_gmem_ARADDR;
	output wire [7:0] sum_35_m_axi_gmem_ARLEN;
	output wire [2:0] sum_35_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_35_m_axi_gmem_ARBURST;
	output wire sum_35_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_35_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_35_m_axi_gmem_ARPROT;
	output wire [3:0] sum_35_m_axi_gmem_ARQOS;
	output wire [3:0] sum_35_m_axi_gmem_ARREGION;
	output wire sum_35_m_axi_gmem_ARUSER;
	output wire sum_35_m_axi_gmem_RREADY;
	input sum_35_m_axi_gmem_RVALID;
	input sum_35_m_axi_gmem_RID;
	input [31:0] sum_35_m_axi_gmem_RDATA;
	input [1:0] sum_35_m_axi_gmem_RRESP;
	input sum_35_m_axi_gmem_RLAST;
	input sum_35_m_axi_gmem_RUSER;
	input sum_35_m_axi_gmem_AWREADY;
	output wire sum_35_m_axi_gmem_AWVALID;
	output wire sum_35_m_axi_gmem_AWID;
	output wire [63:0] sum_35_m_axi_gmem_AWADDR;
	output wire [7:0] sum_35_m_axi_gmem_AWLEN;
	output wire [2:0] sum_35_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_35_m_axi_gmem_AWBURST;
	output wire sum_35_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_35_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_35_m_axi_gmem_AWPROT;
	output wire [3:0] sum_35_m_axi_gmem_AWQOS;
	output wire [3:0] sum_35_m_axi_gmem_AWREGION;
	output wire sum_35_m_axi_gmem_AWUSER;
	input sum_35_m_axi_gmem_WREADY;
	output wire sum_35_m_axi_gmem_WVALID;
	output wire [31:0] sum_35_m_axi_gmem_WDATA;
	output wire [3:0] sum_35_m_axi_gmem_WSTRB;
	output wire sum_35_m_axi_gmem_WLAST;
	output wire sum_35_m_axi_gmem_WUSER;
	output wire sum_35_m_axi_gmem_BREADY;
	input sum_35_m_axi_gmem_BVALID;
	input sum_35_m_axi_gmem_BID;
	input [1:0] sum_35_m_axi_gmem_BRESP;
	input sum_35_m_axi_gmem_BUSER;
	output wire sum_35_s_axi_control_ARREADY;
	input sum_35_s_axi_control_ARVALID;
	input [4:0] sum_35_s_axi_control_ARADDR;
	input sum_35_s_axi_control_RREADY;
	output wire sum_35_s_axi_control_RVALID;
	output wire [31:0] sum_35_s_axi_control_RDATA;
	output wire [1:0] sum_35_s_axi_control_RRESP;
	output wire sum_35_s_axi_control_AWREADY;
	input sum_35_s_axi_control_AWVALID;
	input [4:0] sum_35_s_axi_control_AWADDR;
	output wire sum_35_s_axi_control_WREADY;
	input sum_35_s_axi_control_WVALID;
	input [31:0] sum_35_s_axi_control_WDATA;
	input [3:0] sum_35_s_axi_control_WSTRB;
	input sum_35_s_axi_control_BREADY;
	output wire sum_35_s_axi_control_BVALID;
	output wire [1:0] sum_35_s_axi_control_BRESP;
	input sum_36_m_axi_gmem_ARREADY;
	output wire sum_36_m_axi_gmem_ARVALID;
	output wire sum_36_m_axi_gmem_ARID;
	output wire [63:0] sum_36_m_axi_gmem_ARADDR;
	output wire [7:0] sum_36_m_axi_gmem_ARLEN;
	output wire [2:0] sum_36_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_36_m_axi_gmem_ARBURST;
	output wire sum_36_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_36_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_36_m_axi_gmem_ARPROT;
	output wire [3:0] sum_36_m_axi_gmem_ARQOS;
	output wire [3:0] sum_36_m_axi_gmem_ARREGION;
	output wire sum_36_m_axi_gmem_ARUSER;
	output wire sum_36_m_axi_gmem_RREADY;
	input sum_36_m_axi_gmem_RVALID;
	input sum_36_m_axi_gmem_RID;
	input [31:0] sum_36_m_axi_gmem_RDATA;
	input [1:0] sum_36_m_axi_gmem_RRESP;
	input sum_36_m_axi_gmem_RLAST;
	input sum_36_m_axi_gmem_RUSER;
	input sum_36_m_axi_gmem_AWREADY;
	output wire sum_36_m_axi_gmem_AWVALID;
	output wire sum_36_m_axi_gmem_AWID;
	output wire [63:0] sum_36_m_axi_gmem_AWADDR;
	output wire [7:0] sum_36_m_axi_gmem_AWLEN;
	output wire [2:0] sum_36_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_36_m_axi_gmem_AWBURST;
	output wire sum_36_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_36_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_36_m_axi_gmem_AWPROT;
	output wire [3:0] sum_36_m_axi_gmem_AWQOS;
	output wire [3:0] sum_36_m_axi_gmem_AWREGION;
	output wire sum_36_m_axi_gmem_AWUSER;
	input sum_36_m_axi_gmem_WREADY;
	output wire sum_36_m_axi_gmem_WVALID;
	output wire [31:0] sum_36_m_axi_gmem_WDATA;
	output wire [3:0] sum_36_m_axi_gmem_WSTRB;
	output wire sum_36_m_axi_gmem_WLAST;
	output wire sum_36_m_axi_gmem_WUSER;
	output wire sum_36_m_axi_gmem_BREADY;
	input sum_36_m_axi_gmem_BVALID;
	input sum_36_m_axi_gmem_BID;
	input [1:0] sum_36_m_axi_gmem_BRESP;
	input sum_36_m_axi_gmem_BUSER;
	output wire sum_36_s_axi_control_ARREADY;
	input sum_36_s_axi_control_ARVALID;
	input [4:0] sum_36_s_axi_control_ARADDR;
	input sum_36_s_axi_control_RREADY;
	output wire sum_36_s_axi_control_RVALID;
	output wire [31:0] sum_36_s_axi_control_RDATA;
	output wire [1:0] sum_36_s_axi_control_RRESP;
	output wire sum_36_s_axi_control_AWREADY;
	input sum_36_s_axi_control_AWVALID;
	input [4:0] sum_36_s_axi_control_AWADDR;
	output wire sum_36_s_axi_control_WREADY;
	input sum_36_s_axi_control_WVALID;
	input [31:0] sum_36_s_axi_control_WDATA;
	input [3:0] sum_36_s_axi_control_WSTRB;
	input sum_36_s_axi_control_BREADY;
	output wire sum_36_s_axi_control_BVALID;
	output wire [1:0] sum_36_s_axi_control_BRESP;
	input sum_37_m_axi_gmem_ARREADY;
	output wire sum_37_m_axi_gmem_ARVALID;
	output wire sum_37_m_axi_gmem_ARID;
	output wire [63:0] sum_37_m_axi_gmem_ARADDR;
	output wire [7:0] sum_37_m_axi_gmem_ARLEN;
	output wire [2:0] sum_37_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_37_m_axi_gmem_ARBURST;
	output wire sum_37_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_37_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_37_m_axi_gmem_ARPROT;
	output wire [3:0] sum_37_m_axi_gmem_ARQOS;
	output wire [3:0] sum_37_m_axi_gmem_ARREGION;
	output wire sum_37_m_axi_gmem_ARUSER;
	output wire sum_37_m_axi_gmem_RREADY;
	input sum_37_m_axi_gmem_RVALID;
	input sum_37_m_axi_gmem_RID;
	input [31:0] sum_37_m_axi_gmem_RDATA;
	input [1:0] sum_37_m_axi_gmem_RRESP;
	input sum_37_m_axi_gmem_RLAST;
	input sum_37_m_axi_gmem_RUSER;
	input sum_37_m_axi_gmem_AWREADY;
	output wire sum_37_m_axi_gmem_AWVALID;
	output wire sum_37_m_axi_gmem_AWID;
	output wire [63:0] sum_37_m_axi_gmem_AWADDR;
	output wire [7:0] sum_37_m_axi_gmem_AWLEN;
	output wire [2:0] sum_37_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_37_m_axi_gmem_AWBURST;
	output wire sum_37_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_37_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_37_m_axi_gmem_AWPROT;
	output wire [3:0] sum_37_m_axi_gmem_AWQOS;
	output wire [3:0] sum_37_m_axi_gmem_AWREGION;
	output wire sum_37_m_axi_gmem_AWUSER;
	input sum_37_m_axi_gmem_WREADY;
	output wire sum_37_m_axi_gmem_WVALID;
	output wire [31:0] sum_37_m_axi_gmem_WDATA;
	output wire [3:0] sum_37_m_axi_gmem_WSTRB;
	output wire sum_37_m_axi_gmem_WLAST;
	output wire sum_37_m_axi_gmem_WUSER;
	output wire sum_37_m_axi_gmem_BREADY;
	input sum_37_m_axi_gmem_BVALID;
	input sum_37_m_axi_gmem_BID;
	input [1:0] sum_37_m_axi_gmem_BRESP;
	input sum_37_m_axi_gmem_BUSER;
	output wire sum_37_s_axi_control_ARREADY;
	input sum_37_s_axi_control_ARVALID;
	input [4:0] sum_37_s_axi_control_ARADDR;
	input sum_37_s_axi_control_RREADY;
	output wire sum_37_s_axi_control_RVALID;
	output wire [31:0] sum_37_s_axi_control_RDATA;
	output wire [1:0] sum_37_s_axi_control_RRESP;
	output wire sum_37_s_axi_control_AWREADY;
	input sum_37_s_axi_control_AWVALID;
	input [4:0] sum_37_s_axi_control_AWADDR;
	output wire sum_37_s_axi_control_WREADY;
	input sum_37_s_axi_control_WVALID;
	input [31:0] sum_37_s_axi_control_WDATA;
	input [3:0] sum_37_s_axi_control_WSTRB;
	input sum_37_s_axi_control_BREADY;
	output wire sum_37_s_axi_control_BVALID;
	output wire [1:0] sum_37_s_axi_control_BRESP;
	input sum_38_m_axi_gmem_ARREADY;
	output wire sum_38_m_axi_gmem_ARVALID;
	output wire sum_38_m_axi_gmem_ARID;
	output wire [63:0] sum_38_m_axi_gmem_ARADDR;
	output wire [7:0] sum_38_m_axi_gmem_ARLEN;
	output wire [2:0] sum_38_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_38_m_axi_gmem_ARBURST;
	output wire sum_38_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_38_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_38_m_axi_gmem_ARPROT;
	output wire [3:0] sum_38_m_axi_gmem_ARQOS;
	output wire [3:0] sum_38_m_axi_gmem_ARREGION;
	output wire sum_38_m_axi_gmem_ARUSER;
	output wire sum_38_m_axi_gmem_RREADY;
	input sum_38_m_axi_gmem_RVALID;
	input sum_38_m_axi_gmem_RID;
	input [31:0] sum_38_m_axi_gmem_RDATA;
	input [1:0] sum_38_m_axi_gmem_RRESP;
	input sum_38_m_axi_gmem_RLAST;
	input sum_38_m_axi_gmem_RUSER;
	input sum_38_m_axi_gmem_AWREADY;
	output wire sum_38_m_axi_gmem_AWVALID;
	output wire sum_38_m_axi_gmem_AWID;
	output wire [63:0] sum_38_m_axi_gmem_AWADDR;
	output wire [7:0] sum_38_m_axi_gmem_AWLEN;
	output wire [2:0] sum_38_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_38_m_axi_gmem_AWBURST;
	output wire sum_38_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_38_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_38_m_axi_gmem_AWPROT;
	output wire [3:0] sum_38_m_axi_gmem_AWQOS;
	output wire [3:0] sum_38_m_axi_gmem_AWREGION;
	output wire sum_38_m_axi_gmem_AWUSER;
	input sum_38_m_axi_gmem_WREADY;
	output wire sum_38_m_axi_gmem_WVALID;
	output wire [31:0] sum_38_m_axi_gmem_WDATA;
	output wire [3:0] sum_38_m_axi_gmem_WSTRB;
	output wire sum_38_m_axi_gmem_WLAST;
	output wire sum_38_m_axi_gmem_WUSER;
	output wire sum_38_m_axi_gmem_BREADY;
	input sum_38_m_axi_gmem_BVALID;
	input sum_38_m_axi_gmem_BID;
	input [1:0] sum_38_m_axi_gmem_BRESP;
	input sum_38_m_axi_gmem_BUSER;
	output wire sum_38_s_axi_control_ARREADY;
	input sum_38_s_axi_control_ARVALID;
	input [4:0] sum_38_s_axi_control_ARADDR;
	input sum_38_s_axi_control_RREADY;
	output wire sum_38_s_axi_control_RVALID;
	output wire [31:0] sum_38_s_axi_control_RDATA;
	output wire [1:0] sum_38_s_axi_control_RRESP;
	output wire sum_38_s_axi_control_AWREADY;
	input sum_38_s_axi_control_AWVALID;
	input [4:0] sum_38_s_axi_control_AWADDR;
	output wire sum_38_s_axi_control_WREADY;
	input sum_38_s_axi_control_WVALID;
	input [31:0] sum_38_s_axi_control_WDATA;
	input [3:0] sum_38_s_axi_control_WSTRB;
	input sum_38_s_axi_control_BREADY;
	output wire sum_38_s_axi_control_BVALID;
	output wire [1:0] sum_38_s_axi_control_BRESP;
	input sum_39_m_axi_gmem_ARREADY;
	output wire sum_39_m_axi_gmem_ARVALID;
	output wire sum_39_m_axi_gmem_ARID;
	output wire [63:0] sum_39_m_axi_gmem_ARADDR;
	output wire [7:0] sum_39_m_axi_gmem_ARLEN;
	output wire [2:0] sum_39_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_39_m_axi_gmem_ARBURST;
	output wire sum_39_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_39_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_39_m_axi_gmem_ARPROT;
	output wire [3:0] sum_39_m_axi_gmem_ARQOS;
	output wire [3:0] sum_39_m_axi_gmem_ARREGION;
	output wire sum_39_m_axi_gmem_ARUSER;
	output wire sum_39_m_axi_gmem_RREADY;
	input sum_39_m_axi_gmem_RVALID;
	input sum_39_m_axi_gmem_RID;
	input [31:0] sum_39_m_axi_gmem_RDATA;
	input [1:0] sum_39_m_axi_gmem_RRESP;
	input sum_39_m_axi_gmem_RLAST;
	input sum_39_m_axi_gmem_RUSER;
	input sum_39_m_axi_gmem_AWREADY;
	output wire sum_39_m_axi_gmem_AWVALID;
	output wire sum_39_m_axi_gmem_AWID;
	output wire [63:0] sum_39_m_axi_gmem_AWADDR;
	output wire [7:0] sum_39_m_axi_gmem_AWLEN;
	output wire [2:0] sum_39_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_39_m_axi_gmem_AWBURST;
	output wire sum_39_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_39_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_39_m_axi_gmem_AWPROT;
	output wire [3:0] sum_39_m_axi_gmem_AWQOS;
	output wire [3:0] sum_39_m_axi_gmem_AWREGION;
	output wire sum_39_m_axi_gmem_AWUSER;
	input sum_39_m_axi_gmem_WREADY;
	output wire sum_39_m_axi_gmem_WVALID;
	output wire [31:0] sum_39_m_axi_gmem_WDATA;
	output wire [3:0] sum_39_m_axi_gmem_WSTRB;
	output wire sum_39_m_axi_gmem_WLAST;
	output wire sum_39_m_axi_gmem_WUSER;
	output wire sum_39_m_axi_gmem_BREADY;
	input sum_39_m_axi_gmem_BVALID;
	input sum_39_m_axi_gmem_BID;
	input [1:0] sum_39_m_axi_gmem_BRESP;
	input sum_39_m_axi_gmem_BUSER;
	output wire sum_39_s_axi_control_ARREADY;
	input sum_39_s_axi_control_ARVALID;
	input [4:0] sum_39_s_axi_control_ARADDR;
	input sum_39_s_axi_control_RREADY;
	output wire sum_39_s_axi_control_RVALID;
	output wire [31:0] sum_39_s_axi_control_RDATA;
	output wire [1:0] sum_39_s_axi_control_RRESP;
	output wire sum_39_s_axi_control_AWREADY;
	input sum_39_s_axi_control_AWVALID;
	input [4:0] sum_39_s_axi_control_AWADDR;
	output wire sum_39_s_axi_control_WREADY;
	input sum_39_s_axi_control_WVALID;
	input [31:0] sum_39_s_axi_control_WDATA;
	input [3:0] sum_39_s_axi_control_WSTRB;
	input sum_39_s_axi_control_BREADY;
	output wire sum_39_s_axi_control_BVALID;
	output wire [1:0] sum_39_s_axi_control_BRESP;
	input sum_40_m_axi_gmem_ARREADY;
	output wire sum_40_m_axi_gmem_ARVALID;
	output wire sum_40_m_axi_gmem_ARID;
	output wire [63:0] sum_40_m_axi_gmem_ARADDR;
	output wire [7:0] sum_40_m_axi_gmem_ARLEN;
	output wire [2:0] sum_40_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_40_m_axi_gmem_ARBURST;
	output wire sum_40_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_40_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_40_m_axi_gmem_ARPROT;
	output wire [3:0] sum_40_m_axi_gmem_ARQOS;
	output wire [3:0] sum_40_m_axi_gmem_ARREGION;
	output wire sum_40_m_axi_gmem_ARUSER;
	output wire sum_40_m_axi_gmem_RREADY;
	input sum_40_m_axi_gmem_RVALID;
	input sum_40_m_axi_gmem_RID;
	input [31:0] sum_40_m_axi_gmem_RDATA;
	input [1:0] sum_40_m_axi_gmem_RRESP;
	input sum_40_m_axi_gmem_RLAST;
	input sum_40_m_axi_gmem_RUSER;
	input sum_40_m_axi_gmem_AWREADY;
	output wire sum_40_m_axi_gmem_AWVALID;
	output wire sum_40_m_axi_gmem_AWID;
	output wire [63:0] sum_40_m_axi_gmem_AWADDR;
	output wire [7:0] sum_40_m_axi_gmem_AWLEN;
	output wire [2:0] sum_40_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_40_m_axi_gmem_AWBURST;
	output wire sum_40_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_40_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_40_m_axi_gmem_AWPROT;
	output wire [3:0] sum_40_m_axi_gmem_AWQOS;
	output wire [3:0] sum_40_m_axi_gmem_AWREGION;
	output wire sum_40_m_axi_gmem_AWUSER;
	input sum_40_m_axi_gmem_WREADY;
	output wire sum_40_m_axi_gmem_WVALID;
	output wire [31:0] sum_40_m_axi_gmem_WDATA;
	output wire [3:0] sum_40_m_axi_gmem_WSTRB;
	output wire sum_40_m_axi_gmem_WLAST;
	output wire sum_40_m_axi_gmem_WUSER;
	output wire sum_40_m_axi_gmem_BREADY;
	input sum_40_m_axi_gmem_BVALID;
	input sum_40_m_axi_gmem_BID;
	input [1:0] sum_40_m_axi_gmem_BRESP;
	input sum_40_m_axi_gmem_BUSER;
	output wire sum_40_s_axi_control_ARREADY;
	input sum_40_s_axi_control_ARVALID;
	input [4:0] sum_40_s_axi_control_ARADDR;
	input sum_40_s_axi_control_RREADY;
	output wire sum_40_s_axi_control_RVALID;
	output wire [31:0] sum_40_s_axi_control_RDATA;
	output wire [1:0] sum_40_s_axi_control_RRESP;
	output wire sum_40_s_axi_control_AWREADY;
	input sum_40_s_axi_control_AWVALID;
	input [4:0] sum_40_s_axi_control_AWADDR;
	output wire sum_40_s_axi_control_WREADY;
	input sum_40_s_axi_control_WVALID;
	input [31:0] sum_40_s_axi_control_WDATA;
	input [3:0] sum_40_s_axi_control_WSTRB;
	input sum_40_s_axi_control_BREADY;
	output wire sum_40_s_axi_control_BVALID;
	output wire [1:0] sum_40_s_axi_control_BRESP;
	input sum_41_m_axi_gmem_ARREADY;
	output wire sum_41_m_axi_gmem_ARVALID;
	output wire sum_41_m_axi_gmem_ARID;
	output wire [63:0] sum_41_m_axi_gmem_ARADDR;
	output wire [7:0] sum_41_m_axi_gmem_ARLEN;
	output wire [2:0] sum_41_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_41_m_axi_gmem_ARBURST;
	output wire sum_41_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_41_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_41_m_axi_gmem_ARPROT;
	output wire [3:0] sum_41_m_axi_gmem_ARQOS;
	output wire [3:0] sum_41_m_axi_gmem_ARREGION;
	output wire sum_41_m_axi_gmem_ARUSER;
	output wire sum_41_m_axi_gmem_RREADY;
	input sum_41_m_axi_gmem_RVALID;
	input sum_41_m_axi_gmem_RID;
	input [31:0] sum_41_m_axi_gmem_RDATA;
	input [1:0] sum_41_m_axi_gmem_RRESP;
	input sum_41_m_axi_gmem_RLAST;
	input sum_41_m_axi_gmem_RUSER;
	input sum_41_m_axi_gmem_AWREADY;
	output wire sum_41_m_axi_gmem_AWVALID;
	output wire sum_41_m_axi_gmem_AWID;
	output wire [63:0] sum_41_m_axi_gmem_AWADDR;
	output wire [7:0] sum_41_m_axi_gmem_AWLEN;
	output wire [2:0] sum_41_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_41_m_axi_gmem_AWBURST;
	output wire sum_41_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_41_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_41_m_axi_gmem_AWPROT;
	output wire [3:0] sum_41_m_axi_gmem_AWQOS;
	output wire [3:0] sum_41_m_axi_gmem_AWREGION;
	output wire sum_41_m_axi_gmem_AWUSER;
	input sum_41_m_axi_gmem_WREADY;
	output wire sum_41_m_axi_gmem_WVALID;
	output wire [31:0] sum_41_m_axi_gmem_WDATA;
	output wire [3:0] sum_41_m_axi_gmem_WSTRB;
	output wire sum_41_m_axi_gmem_WLAST;
	output wire sum_41_m_axi_gmem_WUSER;
	output wire sum_41_m_axi_gmem_BREADY;
	input sum_41_m_axi_gmem_BVALID;
	input sum_41_m_axi_gmem_BID;
	input [1:0] sum_41_m_axi_gmem_BRESP;
	input sum_41_m_axi_gmem_BUSER;
	output wire sum_41_s_axi_control_ARREADY;
	input sum_41_s_axi_control_ARVALID;
	input [4:0] sum_41_s_axi_control_ARADDR;
	input sum_41_s_axi_control_RREADY;
	output wire sum_41_s_axi_control_RVALID;
	output wire [31:0] sum_41_s_axi_control_RDATA;
	output wire [1:0] sum_41_s_axi_control_RRESP;
	output wire sum_41_s_axi_control_AWREADY;
	input sum_41_s_axi_control_AWVALID;
	input [4:0] sum_41_s_axi_control_AWADDR;
	output wire sum_41_s_axi_control_WREADY;
	input sum_41_s_axi_control_WVALID;
	input [31:0] sum_41_s_axi_control_WDATA;
	input [3:0] sum_41_s_axi_control_WSTRB;
	input sum_41_s_axi_control_BREADY;
	output wire sum_41_s_axi_control_BVALID;
	output wire [1:0] sum_41_s_axi_control_BRESP;
	input sum_42_m_axi_gmem_ARREADY;
	output wire sum_42_m_axi_gmem_ARVALID;
	output wire sum_42_m_axi_gmem_ARID;
	output wire [63:0] sum_42_m_axi_gmem_ARADDR;
	output wire [7:0] sum_42_m_axi_gmem_ARLEN;
	output wire [2:0] sum_42_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_42_m_axi_gmem_ARBURST;
	output wire sum_42_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_42_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_42_m_axi_gmem_ARPROT;
	output wire [3:0] sum_42_m_axi_gmem_ARQOS;
	output wire [3:0] sum_42_m_axi_gmem_ARREGION;
	output wire sum_42_m_axi_gmem_ARUSER;
	output wire sum_42_m_axi_gmem_RREADY;
	input sum_42_m_axi_gmem_RVALID;
	input sum_42_m_axi_gmem_RID;
	input [31:0] sum_42_m_axi_gmem_RDATA;
	input [1:0] sum_42_m_axi_gmem_RRESP;
	input sum_42_m_axi_gmem_RLAST;
	input sum_42_m_axi_gmem_RUSER;
	input sum_42_m_axi_gmem_AWREADY;
	output wire sum_42_m_axi_gmem_AWVALID;
	output wire sum_42_m_axi_gmem_AWID;
	output wire [63:0] sum_42_m_axi_gmem_AWADDR;
	output wire [7:0] sum_42_m_axi_gmem_AWLEN;
	output wire [2:0] sum_42_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_42_m_axi_gmem_AWBURST;
	output wire sum_42_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_42_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_42_m_axi_gmem_AWPROT;
	output wire [3:0] sum_42_m_axi_gmem_AWQOS;
	output wire [3:0] sum_42_m_axi_gmem_AWREGION;
	output wire sum_42_m_axi_gmem_AWUSER;
	input sum_42_m_axi_gmem_WREADY;
	output wire sum_42_m_axi_gmem_WVALID;
	output wire [31:0] sum_42_m_axi_gmem_WDATA;
	output wire [3:0] sum_42_m_axi_gmem_WSTRB;
	output wire sum_42_m_axi_gmem_WLAST;
	output wire sum_42_m_axi_gmem_WUSER;
	output wire sum_42_m_axi_gmem_BREADY;
	input sum_42_m_axi_gmem_BVALID;
	input sum_42_m_axi_gmem_BID;
	input [1:0] sum_42_m_axi_gmem_BRESP;
	input sum_42_m_axi_gmem_BUSER;
	output wire sum_42_s_axi_control_ARREADY;
	input sum_42_s_axi_control_ARVALID;
	input [4:0] sum_42_s_axi_control_ARADDR;
	input sum_42_s_axi_control_RREADY;
	output wire sum_42_s_axi_control_RVALID;
	output wire [31:0] sum_42_s_axi_control_RDATA;
	output wire [1:0] sum_42_s_axi_control_RRESP;
	output wire sum_42_s_axi_control_AWREADY;
	input sum_42_s_axi_control_AWVALID;
	input [4:0] sum_42_s_axi_control_AWADDR;
	output wire sum_42_s_axi_control_WREADY;
	input sum_42_s_axi_control_WVALID;
	input [31:0] sum_42_s_axi_control_WDATA;
	input [3:0] sum_42_s_axi_control_WSTRB;
	input sum_42_s_axi_control_BREADY;
	output wire sum_42_s_axi_control_BVALID;
	output wire [1:0] sum_42_s_axi_control_BRESP;
	input sum_43_m_axi_gmem_ARREADY;
	output wire sum_43_m_axi_gmem_ARVALID;
	output wire sum_43_m_axi_gmem_ARID;
	output wire [63:0] sum_43_m_axi_gmem_ARADDR;
	output wire [7:0] sum_43_m_axi_gmem_ARLEN;
	output wire [2:0] sum_43_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_43_m_axi_gmem_ARBURST;
	output wire sum_43_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_43_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_43_m_axi_gmem_ARPROT;
	output wire [3:0] sum_43_m_axi_gmem_ARQOS;
	output wire [3:0] sum_43_m_axi_gmem_ARREGION;
	output wire sum_43_m_axi_gmem_ARUSER;
	output wire sum_43_m_axi_gmem_RREADY;
	input sum_43_m_axi_gmem_RVALID;
	input sum_43_m_axi_gmem_RID;
	input [31:0] sum_43_m_axi_gmem_RDATA;
	input [1:0] sum_43_m_axi_gmem_RRESP;
	input sum_43_m_axi_gmem_RLAST;
	input sum_43_m_axi_gmem_RUSER;
	input sum_43_m_axi_gmem_AWREADY;
	output wire sum_43_m_axi_gmem_AWVALID;
	output wire sum_43_m_axi_gmem_AWID;
	output wire [63:0] sum_43_m_axi_gmem_AWADDR;
	output wire [7:0] sum_43_m_axi_gmem_AWLEN;
	output wire [2:0] sum_43_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_43_m_axi_gmem_AWBURST;
	output wire sum_43_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_43_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_43_m_axi_gmem_AWPROT;
	output wire [3:0] sum_43_m_axi_gmem_AWQOS;
	output wire [3:0] sum_43_m_axi_gmem_AWREGION;
	output wire sum_43_m_axi_gmem_AWUSER;
	input sum_43_m_axi_gmem_WREADY;
	output wire sum_43_m_axi_gmem_WVALID;
	output wire [31:0] sum_43_m_axi_gmem_WDATA;
	output wire [3:0] sum_43_m_axi_gmem_WSTRB;
	output wire sum_43_m_axi_gmem_WLAST;
	output wire sum_43_m_axi_gmem_WUSER;
	output wire sum_43_m_axi_gmem_BREADY;
	input sum_43_m_axi_gmem_BVALID;
	input sum_43_m_axi_gmem_BID;
	input [1:0] sum_43_m_axi_gmem_BRESP;
	input sum_43_m_axi_gmem_BUSER;
	output wire sum_43_s_axi_control_ARREADY;
	input sum_43_s_axi_control_ARVALID;
	input [4:0] sum_43_s_axi_control_ARADDR;
	input sum_43_s_axi_control_RREADY;
	output wire sum_43_s_axi_control_RVALID;
	output wire [31:0] sum_43_s_axi_control_RDATA;
	output wire [1:0] sum_43_s_axi_control_RRESP;
	output wire sum_43_s_axi_control_AWREADY;
	input sum_43_s_axi_control_AWVALID;
	input [4:0] sum_43_s_axi_control_AWADDR;
	output wire sum_43_s_axi_control_WREADY;
	input sum_43_s_axi_control_WVALID;
	input [31:0] sum_43_s_axi_control_WDATA;
	input [3:0] sum_43_s_axi_control_WSTRB;
	input sum_43_s_axi_control_BREADY;
	output wire sum_43_s_axi_control_BVALID;
	output wire [1:0] sum_43_s_axi_control_BRESP;
	input sum_44_m_axi_gmem_ARREADY;
	output wire sum_44_m_axi_gmem_ARVALID;
	output wire sum_44_m_axi_gmem_ARID;
	output wire [63:0] sum_44_m_axi_gmem_ARADDR;
	output wire [7:0] sum_44_m_axi_gmem_ARLEN;
	output wire [2:0] sum_44_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_44_m_axi_gmem_ARBURST;
	output wire sum_44_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_44_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_44_m_axi_gmem_ARPROT;
	output wire [3:0] sum_44_m_axi_gmem_ARQOS;
	output wire [3:0] sum_44_m_axi_gmem_ARREGION;
	output wire sum_44_m_axi_gmem_ARUSER;
	output wire sum_44_m_axi_gmem_RREADY;
	input sum_44_m_axi_gmem_RVALID;
	input sum_44_m_axi_gmem_RID;
	input [31:0] sum_44_m_axi_gmem_RDATA;
	input [1:0] sum_44_m_axi_gmem_RRESP;
	input sum_44_m_axi_gmem_RLAST;
	input sum_44_m_axi_gmem_RUSER;
	input sum_44_m_axi_gmem_AWREADY;
	output wire sum_44_m_axi_gmem_AWVALID;
	output wire sum_44_m_axi_gmem_AWID;
	output wire [63:0] sum_44_m_axi_gmem_AWADDR;
	output wire [7:0] sum_44_m_axi_gmem_AWLEN;
	output wire [2:0] sum_44_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_44_m_axi_gmem_AWBURST;
	output wire sum_44_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_44_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_44_m_axi_gmem_AWPROT;
	output wire [3:0] sum_44_m_axi_gmem_AWQOS;
	output wire [3:0] sum_44_m_axi_gmem_AWREGION;
	output wire sum_44_m_axi_gmem_AWUSER;
	input sum_44_m_axi_gmem_WREADY;
	output wire sum_44_m_axi_gmem_WVALID;
	output wire [31:0] sum_44_m_axi_gmem_WDATA;
	output wire [3:0] sum_44_m_axi_gmem_WSTRB;
	output wire sum_44_m_axi_gmem_WLAST;
	output wire sum_44_m_axi_gmem_WUSER;
	output wire sum_44_m_axi_gmem_BREADY;
	input sum_44_m_axi_gmem_BVALID;
	input sum_44_m_axi_gmem_BID;
	input [1:0] sum_44_m_axi_gmem_BRESP;
	input sum_44_m_axi_gmem_BUSER;
	output wire sum_44_s_axi_control_ARREADY;
	input sum_44_s_axi_control_ARVALID;
	input [4:0] sum_44_s_axi_control_ARADDR;
	input sum_44_s_axi_control_RREADY;
	output wire sum_44_s_axi_control_RVALID;
	output wire [31:0] sum_44_s_axi_control_RDATA;
	output wire [1:0] sum_44_s_axi_control_RRESP;
	output wire sum_44_s_axi_control_AWREADY;
	input sum_44_s_axi_control_AWVALID;
	input [4:0] sum_44_s_axi_control_AWADDR;
	output wire sum_44_s_axi_control_WREADY;
	input sum_44_s_axi_control_WVALID;
	input [31:0] sum_44_s_axi_control_WDATA;
	input [3:0] sum_44_s_axi_control_WSTRB;
	input sum_44_s_axi_control_BREADY;
	output wire sum_44_s_axi_control_BVALID;
	output wire [1:0] sum_44_s_axi_control_BRESP;
	input sum_45_m_axi_gmem_ARREADY;
	output wire sum_45_m_axi_gmem_ARVALID;
	output wire sum_45_m_axi_gmem_ARID;
	output wire [63:0] sum_45_m_axi_gmem_ARADDR;
	output wire [7:0] sum_45_m_axi_gmem_ARLEN;
	output wire [2:0] sum_45_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_45_m_axi_gmem_ARBURST;
	output wire sum_45_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_45_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_45_m_axi_gmem_ARPROT;
	output wire [3:0] sum_45_m_axi_gmem_ARQOS;
	output wire [3:0] sum_45_m_axi_gmem_ARREGION;
	output wire sum_45_m_axi_gmem_ARUSER;
	output wire sum_45_m_axi_gmem_RREADY;
	input sum_45_m_axi_gmem_RVALID;
	input sum_45_m_axi_gmem_RID;
	input [31:0] sum_45_m_axi_gmem_RDATA;
	input [1:0] sum_45_m_axi_gmem_RRESP;
	input sum_45_m_axi_gmem_RLAST;
	input sum_45_m_axi_gmem_RUSER;
	input sum_45_m_axi_gmem_AWREADY;
	output wire sum_45_m_axi_gmem_AWVALID;
	output wire sum_45_m_axi_gmem_AWID;
	output wire [63:0] sum_45_m_axi_gmem_AWADDR;
	output wire [7:0] sum_45_m_axi_gmem_AWLEN;
	output wire [2:0] sum_45_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_45_m_axi_gmem_AWBURST;
	output wire sum_45_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_45_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_45_m_axi_gmem_AWPROT;
	output wire [3:0] sum_45_m_axi_gmem_AWQOS;
	output wire [3:0] sum_45_m_axi_gmem_AWREGION;
	output wire sum_45_m_axi_gmem_AWUSER;
	input sum_45_m_axi_gmem_WREADY;
	output wire sum_45_m_axi_gmem_WVALID;
	output wire [31:0] sum_45_m_axi_gmem_WDATA;
	output wire [3:0] sum_45_m_axi_gmem_WSTRB;
	output wire sum_45_m_axi_gmem_WLAST;
	output wire sum_45_m_axi_gmem_WUSER;
	output wire sum_45_m_axi_gmem_BREADY;
	input sum_45_m_axi_gmem_BVALID;
	input sum_45_m_axi_gmem_BID;
	input [1:0] sum_45_m_axi_gmem_BRESP;
	input sum_45_m_axi_gmem_BUSER;
	output wire sum_45_s_axi_control_ARREADY;
	input sum_45_s_axi_control_ARVALID;
	input [4:0] sum_45_s_axi_control_ARADDR;
	input sum_45_s_axi_control_RREADY;
	output wire sum_45_s_axi_control_RVALID;
	output wire [31:0] sum_45_s_axi_control_RDATA;
	output wire [1:0] sum_45_s_axi_control_RRESP;
	output wire sum_45_s_axi_control_AWREADY;
	input sum_45_s_axi_control_AWVALID;
	input [4:0] sum_45_s_axi_control_AWADDR;
	output wire sum_45_s_axi_control_WREADY;
	input sum_45_s_axi_control_WVALID;
	input [31:0] sum_45_s_axi_control_WDATA;
	input [3:0] sum_45_s_axi_control_WSTRB;
	input sum_45_s_axi_control_BREADY;
	output wire sum_45_s_axi_control_BVALID;
	output wire [1:0] sum_45_s_axi_control_BRESP;
	input sum_46_m_axi_gmem_ARREADY;
	output wire sum_46_m_axi_gmem_ARVALID;
	output wire sum_46_m_axi_gmem_ARID;
	output wire [63:0] sum_46_m_axi_gmem_ARADDR;
	output wire [7:0] sum_46_m_axi_gmem_ARLEN;
	output wire [2:0] sum_46_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_46_m_axi_gmem_ARBURST;
	output wire sum_46_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_46_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_46_m_axi_gmem_ARPROT;
	output wire [3:0] sum_46_m_axi_gmem_ARQOS;
	output wire [3:0] sum_46_m_axi_gmem_ARREGION;
	output wire sum_46_m_axi_gmem_ARUSER;
	output wire sum_46_m_axi_gmem_RREADY;
	input sum_46_m_axi_gmem_RVALID;
	input sum_46_m_axi_gmem_RID;
	input [31:0] sum_46_m_axi_gmem_RDATA;
	input [1:0] sum_46_m_axi_gmem_RRESP;
	input sum_46_m_axi_gmem_RLAST;
	input sum_46_m_axi_gmem_RUSER;
	input sum_46_m_axi_gmem_AWREADY;
	output wire sum_46_m_axi_gmem_AWVALID;
	output wire sum_46_m_axi_gmem_AWID;
	output wire [63:0] sum_46_m_axi_gmem_AWADDR;
	output wire [7:0] sum_46_m_axi_gmem_AWLEN;
	output wire [2:0] sum_46_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_46_m_axi_gmem_AWBURST;
	output wire sum_46_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_46_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_46_m_axi_gmem_AWPROT;
	output wire [3:0] sum_46_m_axi_gmem_AWQOS;
	output wire [3:0] sum_46_m_axi_gmem_AWREGION;
	output wire sum_46_m_axi_gmem_AWUSER;
	input sum_46_m_axi_gmem_WREADY;
	output wire sum_46_m_axi_gmem_WVALID;
	output wire [31:0] sum_46_m_axi_gmem_WDATA;
	output wire [3:0] sum_46_m_axi_gmem_WSTRB;
	output wire sum_46_m_axi_gmem_WLAST;
	output wire sum_46_m_axi_gmem_WUSER;
	output wire sum_46_m_axi_gmem_BREADY;
	input sum_46_m_axi_gmem_BVALID;
	input sum_46_m_axi_gmem_BID;
	input [1:0] sum_46_m_axi_gmem_BRESP;
	input sum_46_m_axi_gmem_BUSER;
	output wire sum_46_s_axi_control_ARREADY;
	input sum_46_s_axi_control_ARVALID;
	input [4:0] sum_46_s_axi_control_ARADDR;
	input sum_46_s_axi_control_RREADY;
	output wire sum_46_s_axi_control_RVALID;
	output wire [31:0] sum_46_s_axi_control_RDATA;
	output wire [1:0] sum_46_s_axi_control_RRESP;
	output wire sum_46_s_axi_control_AWREADY;
	input sum_46_s_axi_control_AWVALID;
	input [4:0] sum_46_s_axi_control_AWADDR;
	output wire sum_46_s_axi_control_WREADY;
	input sum_46_s_axi_control_WVALID;
	input [31:0] sum_46_s_axi_control_WDATA;
	input [3:0] sum_46_s_axi_control_WSTRB;
	input sum_46_s_axi_control_BREADY;
	output wire sum_46_s_axi_control_BVALID;
	output wire [1:0] sum_46_s_axi_control_BRESP;
	input sum_47_m_axi_gmem_ARREADY;
	output wire sum_47_m_axi_gmem_ARVALID;
	output wire sum_47_m_axi_gmem_ARID;
	output wire [63:0] sum_47_m_axi_gmem_ARADDR;
	output wire [7:0] sum_47_m_axi_gmem_ARLEN;
	output wire [2:0] sum_47_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_47_m_axi_gmem_ARBURST;
	output wire sum_47_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_47_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_47_m_axi_gmem_ARPROT;
	output wire [3:0] sum_47_m_axi_gmem_ARQOS;
	output wire [3:0] sum_47_m_axi_gmem_ARREGION;
	output wire sum_47_m_axi_gmem_ARUSER;
	output wire sum_47_m_axi_gmem_RREADY;
	input sum_47_m_axi_gmem_RVALID;
	input sum_47_m_axi_gmem_RID;
	input [31:0] sum_47_m_axi_gmem_RDATA;
	input [1:0] sum_47_m_axi_gmem_RRESP;
	input sum_47_m_axi_gmem_RLAST;
	input sum_47_m_axi_gmem_RUSER;
	input sum_47_m_axi_gmem_AWREADY;
	output wire sum_47_m_axi_gmem_AWVALID;
	output wire sum_47_m_axi_gmem_AWID;
	output wire [63:0] sum_47_m_axi_gmem_AWADDR;
	output wire [7:0] sum_47_m_axi_gmem_AWLEN;
	output wire [2:0] sum_47_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_47_m_axi_gmem_AWBURST;
	output wire sum_47_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_47_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_47_m_axi_gmem_AWPROT;
	output wire [3:0] sum_47_m_axi_gmem_AWQOS;
	output wire [3:0] sum_47_m_axi_gmem_AWREGION;
	output wire sum_47_m_axi_gmem_AWUSER;
	input sum_47_m_axi_gmem_WREADY;
	output wire sum_47_m_axi_gmem_WVALID;
	output wire [31:0] sum_47_m_axi_gmem_WDATA;
	output wire [3:0] sum_47_m_axi_gmem_WSTRB;
	output wire sum_47_m_axi_gmem_WLAST;
	output wire sum_47_m_axi_gmem_WUSER;
	output wire sum_47_m_axi_gmem_BREADY;
	input sum_47_m_axi_gmem_BVALID;
	input sum_47_m_axi_gmem_BID;
	input [1:0] sum_47_m_axi_gmem_BRESP;
	input sum_47_m_axi_gmem_BUSER;
	output wire sum_47_s_axi_control_ARREADY;
	input sum_47_s_axi_control_ARVALID;
	input [4:0] sum_47_s_axi_control_ARADDR;
	input sum_47_s_axi_control_RREADY;
	output wire sum_47_s_axi_control_RVALID;
	output wire [31:0] sum_47_s_axi_control_RDATA;
	output wire [1:0] sum_47_s_axi_control_RRESP;
	output wire sum_47_s_axi_control_AWREADY;
	input sum_47_s_axi_control_AWVALID;
	input [4:0] sum_47_s_axi_control_AWADDR;
	output wire sum_47_s_axi_control_WREADY;
	input sum_47_s_axi_control_WVALID;
	input [31:0] sum_47_s_axi_control_WDATA;
	input [3:0] sum_47_s_axi_control_WSTRB;
	input sum_47_s_axi_control_BREADY;
	output wire sum_47_s_axi_control_BVALID;
	output wire [1:0] sum_47_s_axi_control_BRESP;
	input sum_48_m_axi_gmem_ARREADY;
	output wire sum_48_m_axi_gmem_ARVALID;
	output wire sum_48_m_axi_gmem_ARID;
	output wire [63:0] sum_48_m_axi_gmem_ARADDR;
	output wire [7:0] sum_48_m_axi_gmem_ARLEN;
	output wire [2:0] sum_48_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_48_m_axi_gmem_ARBURST;
	output wire sum_48_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_48_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_48_m_axi_gmem_ARPROT;
	output wire [3:0] sum_48_m_axi_gmem_ARQOS;
	output wire [3:0] sum_48_m_axi_gmem_ARREGION;
	output wire sum_48_m_axi_gmem_ARUSER;
	output wire sum_48_m_axi_gmem_RREADY;
	input sum_48_m_axi_gmem_RVALID;
	input sum_48_m_axi_gmem_RID;
	input [31:0] sum_48_m_axi_gmem_RDATA;
	input [1:0] sum_48_m_axi_gmem_RRESP;
	input sum_48_m_axi_gmem_RLAST;
	input sum_48_m_axi_gmem_RUSER;
	input sum_48_m_axi_gmem_AWREADY;
	output wire sum_48_m_axi_gmem_AWVALID;
	output wire sum_48_m_axi_gmem_AWID;
	output wire [63:0] sum_48_m_axi_gmem_AWADDR;
	output wire [7:0] sum_48_m_axi_gmem_AWLEN;
	output wire [2:0] sum_48_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_48_m_axi_gmem_AWBURST;
	output wire sum_48_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_48_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_48_m_axi_gmem_AWPROT;
	output wire [3:0] sum_48_m_axi_gmem_AWQOS;
	output wire [3:0] sum_48_m_axi_gmem_AWREGION;
	output wire sum_48_m_axi_gmem_AWUSER;
	input sum_48_m_axi_gmem_WREADY;
	output wire sum_48_m_axi_gmem_WVALID;
	output wire [31:0] sum_48_m_axi_gmem_WDATA;
	output wire [3:0] sum_48_m_axi_gmem_WSTRB;
	output wire sum_48_m_axi_gmem_WLAST;
	output wire sum_48_m_axi_gmem_WUSER;
	output wire sum_48_m_axi_gmem_BREADY;
	input sum_48_m_axi_gmem_BVALID;
	input sum_48_m_axi_gmem_BID;
	input [1:0] sum_48_m_axi_gmem_BRESP;
	input sum_48_m_axi_gmem_BUSER;
	output wire sum_48_s_axi_control_ARREADY;
	input sum_48_s_axi_control_ARVALID;
	input [4:0] sum_48_s_axi_control_ARADDR;
	input sum_48_s_axi_control_RREADY;
	output wire sum_48_s_axi_control_RVALID;
	output wire [31:0] sum_48_s_axi_control_RDATA;
	output wire [1:0] sum_48_s_axi_control_RRESP;
	output wire sum_48_s_axi_control_AWREADY;
	input sum_48_s_axi_control_AWVALID;
	input [4:0] sum_48_s_axi_control_AWADDR;
	output wire sum_48_s_axi_control_WREADY;
	input sum_48_s_axi_control_WVALID;
	input [31:0] sum_48_s_axi_control_WDATA;
	input [3:0] sum_48_s_axi_control_WSTRB;
	input sum_48_s_axi_control_BREADY;
	output wire sum_48_s_axi_control_BVALID;
	output wire [1:0] sum_48_s_axi_control_BRESP;
	input sum_49_m_axi_gmem_ARREADY;
	output wire sum_49_m_axi_gmem_ARVALID;
	output wire sum_49_m_axi_gmem_ARID;
	output wire [63:0] sum_49_m_axi_gmem_ARADDR;
	output wire [7:0] sum_49_m_axi_gmem_ARLEN;
	output wire [2:0] sum_49_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_49_m_axi_gmem_ARBURST;
	output wire sum_49_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_49_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_49_m_axi_gmem_ARPROT;
	output wire [3:0] sum_49_m_axi_gmem_ARQOS;
	output wire [3:0] sum_49_m_axi_gmem_ARREGION;
	output wire sum_49_m_axi_gmem_ARUSER;
	output wire sum_49_m_axi_gmem_RREADY;
	input sum_49_m_axi_gmem_RVALID;
	input sum_49_m_axi_gmem_RID;
	input [31:0] sum_49_m_axi_gmem_RDATA;
	input [1:0] sum_49_m_axi_gmem_RRESP;
	input sum_49_m_axi_gmem_RLAST;
	input sum_49_m_axi_gmem_RUSER;
	input sum_49_m_axi_gmem_AWREADY;
	output wire sum_49_m_axi_gmem_AWVALID;
	output wire sum_49_m_axi_gmem_AWID;
	output wire [63:0] sum_49_m_axi_gmem_AWADDR;
	output wire [7:0] sum_49_m_axi_gmem_AWLEN;
	output wire [2:0] sum_49_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_49_m_axi_gmem_AWBURST;
	output wire sum_49_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_49_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_49_m_axi_gmem_AWPROT;
	output wire [3:0] sum_49_m_axi_gmem_AWQOS;
	output wire [3:0] sum_49_m_axi_gmem_AWREGION;
	output wire sum_49_m_axi_gmem_AWUSER;
	input sum_49_m_axi_gmem_WREADY;
	output wire sum_49_m_axi_gmem_WVALID;
	output wire [31:0] sum_49_m_axi_gmem_WDATA;
	output wire [3:0] sum_49_m_axi_gmem_WSTRB;
	output wire sum_49_m_axi_gmem_WLAST;
	output wire sum_49_m_axi_gmem_WUSER;
	output wire sum_49_m_axi_gmem_BREADY;
	input sum_49_m_axi_gmem_BVALID;
	input sum_49_m_axi_gmem_BID;
	input [1:0] sum_49_m_axi_gmem_BRESP;
	input sum_49_m_axi_gmem_BUSER;
	output wire sum_49_s_axi_control_ARREADY;
	input sum_49_s_axi_control_ARVALID;
	input [4:0] sum_49_s_axi_control_ARADDR;
	input sum_49_s_axi_control_RREADY;
	output wire sum_49_s_axi_control_RVALID;
	output wire [31:0] sum_49_s_axi_control_RDATA;
	output wire [1:0] sum_49_s_axi_control_RRESP;
	output wire sum_49_s_axi_control_AWREADY;
	input sum_49_s_axi_control_AWVALID;
	input [4:0] sum_49_s_axi_control_AWADDR;
	output wire sum_49_s_axi_control_WREADY;
	input sum_49_s_axi_control_WVALID;
	input [31:0] sum_49_s_axi_control_WDATA;
	input [3:0] sum_49_s_axi_control_WSTRB;
	input sum_49_s_axi_control_BREADY;
	output wire sum_49_s_axi_control_BVALID;
	output wire [1:0] sum_49_s_axi_control_BRESP;
	input sum_50_m_axi_gmem_ARREADY;
	output wire sum_50_m_axi_gmem_ARVALID;
	output wire sum_50_m_axi_gmem_ARID;
	output wire [63:0] sum_50_m_axi_gmem_ARADDR;
	output wire [7:0] sum_50_m_axi_gmem_ARLEN;
	output wire [2:0] sum_50_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_50_m_axi_gmem_ARBURST;
	output wire sum_50_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_50_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_50_m_axi_gmem_ARPROT;
	output wire [3:0] sum_50_m_axi_gmem_ARQOS;
	output wire [3:0] sum_50_m_axi_gmem_ARREGION;
	output wire sum_50_m_axi_gmem_ARUSER;
	output wire sum_50_m_axi_gmem_RREADY;
	input sum_50_m_axi_gmem_RVALID;
	input sum_50_m_axi_gmem_RID;
	input [31:0] sum_50_m_axi_gmem_RDATA;
	input [1:0] sum_50_m_axi_gmem_RRESP;
	input sum_50_m_axi_gmem_RLAST;
	input sum_50_m_axi_gmem_RUSER;
	input sum_50_m_axi_gmem_AWREADY;
	output wire sum_50_m_axi_gmem_AWVALID;
	output wire sum_50_m_axi_gmem_AWID;
	output wire [63:0] sum_50_m_axi_gmem_AWADDR;
	output wire [7:0] sum_50_m_axi_gmem_AWLEN;
	output wire [2:0] sum_50_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_50_m_axi_gmem_AWBURST;
	output wire sum_50_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_50_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_50_m_axi_gmem_AWPROT;
	output wire [3:0] sum_50_m_axi_gmem_AWQOS;
	output wire [3:0] sum_50_m_axi_gmem_AWREGION;
	output wire sum_50_m_axi_gmem_AWUSER;
	input sum_50_m_axi_gmem_WREADY;
	output wire sum_50_m_axi_gmem_WVALID;
	output wire [31:0] sum_50_m_axi_gmem_WDATA;
	output wire [3:0] sum_50_m_axi_gmem_WSTRB;
	output wire sum_50_m_axi_gmem_WLAST;
	output wire sum_50_m_axi_gmem_WUSER;
	output wire sum_50_m_axi_gmem_BREADY;
	input sum_50_m_axi_gmem_BVALID;
	input sum_50_m_axi_gmem_BID;
	input [1:0] sum_50_m_axi_gmem_BRESP;
	input sum_50_m_axi_gmem_BUSER;
	output wire sum_50_s_axi_control_ARREADY;
	input sum_50_s_axi_control_ARVALID;
	input [4:0] sum_50_s_axi_control_ARADDR;
	input sum_50_s_axi_control_RREADY;
	output wire sum_50_s_axi_control_RVALID;
	output wire [31:0] sum_50_s_axi_control_RDATA;
	output wire [1:0] sum_50_s_axi_control_RRESP;
	output wire sum_50_s_axi_control_AWREADY;
	input sum_50_s_axi_control_AWVALID;
	input [4:0] sum_50_s_axi_control_AWADDR;
	output wire sum_50_s_axi_control_WREADY;
	input sum_50_s_axi_control_WVALID;
	input [31:0] sum_50_s_axi_control_WDATA;
	input [3:0] sum_50_s_axi_control_WSTRB;
	input sum_50_s_axi_control_BREADY;
	output wire sum_50_s_axi_control_BVALID;
	output wire [1:0] sum_50_s_axi_control_BRESP;
	input sum_51_m_axi_gmem_ARREADY;
	output wire sum_51_m_axi_gmem_ARVALID;
	output wire sum_51_m_axi_gmem_ARID;
	output wire [63:0] sum_51_m_axi_gmem_ARADDR;
	output wire [7:0] sum_51_m_axi_gmem_ARLEN;
	output wire [2:0] sum_51_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_51_m_axi_gmem_ARBURST;
	output wire sum_51_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_51_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_51_m_axi_gmem_ARPROT;
	output wire [3:0] sum_51_m_axi_gmem_ARQOS;
	output wire [3:0] sum_51_m_axi_gmem_ARREGION;
	output wire sum_51_m_axi_gmem_ARUSER;
	output wire sum_51_m_axi_gmem_RREADY;
	input sum_51_m_axi_gmem_RVALID;
	input sum_51_m_axi_gmem_RID;
	input [31:0] sum_51_m_axi_gmem_RDATA;
	input [1:0] sum_51_m_axi_gmem_RRESP;
	input sum_51_m_axi_gmem_RLAST;
	input sum_51_m_axi_gmem_RUSER;
	input sum_51_m_axi_gmem_AWREADY;
	output wire sum_51_m_axi_gmem_AWVALID;
	output wire sum_51_m_axi_gmem_AWID;
	output wire [63:0] sum_51_m_axi_gmem_AWADDR;
	output wire [7:0] sum_51_m_axi_gmem_AWLEN;
	output wire [2:0] sum_51_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_51_m_axi_gmem_AWBURST;
	output wire sum_51_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_51_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_51_m_axi_gmem_AWPROT;
	output wire [3:0] sum_51_m_axi_gmem_AWQOS;
	output wire [3:0] sum_51_m_axi_gmem_AWREGION;
	output wire sum_51_m_axi_gmem_AWUSER;
	input sum_51_m_axi_gmem_WREADY;
	output wire sum_51_m_axi_gmem_WVALID;
	output wire [31:0] sum_51_m_axi_gmem_WDATA;
	output wire [3:0] sum_51_m_axi_gmem_WSTRB;
	output wire sum_51_m_axi_gmem_WLAST;
	output wire sum_51_m_axi_gmem_WUSER;
	output wire sum_51_m_axi_gmem_BREADY;
	input sum_51_m_axi_gmem_BVALID;
	input sum_51_m_axi_gmem_BID;
	input [1:0] sum_51_m_axi_gmem_BRESP;
	input sum_51_m_axi_gmem_BUSER;
	output wire sum_51_s_axi_control_ARREADY;
	input sum_51_s_axi_control_ARVALID;
	input [4:0] sum_51_s_axi_control_ARADDR;
	input sum_51_s_axi_control_RREADY;
	output wire sum_51_s_axi_control_RVALID;
	output wire [31:0] sum_51_s_axi_control_RDATA;
	output wire [1:0] sum_51_s_axi_control_RRESP;
	output wire sum_51_s_axi_control_AWREADY;
	input sum_51_s_axi_control_AWVALID;
	input [4:0] sum_51_s_axi_control_AWADDR;
	output wire sum_51_s_axi_control_WREADY;
	input sum_51_s_axi_control_WVALID;
	input [31:0] sum_51_s_axi_control_WDATA;
	input [3:0] sum_51_s_axi_control_WSTRB;
	input sum_51_s_axi_control_BREADY;
	output wire sum_51_s_axi_control_BVALID;
	output wire [1:0] sum_51_s_axi_control_BRESP;
	input sum_52_m_axi_gmem_ARREADY;
	output wire sum_52_m_axi_gmem_ARVALID;
	output wire sum_52_m_axi_gmem_ARID;
	output wire [63:0] sum_52_m_axi_gmem_ARADDR;
	output wire [7:0] sum_52_m_axi_gmem_ARLEN;
	output wire [2:0] sum_52_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_52_m_axi_gmem_ARBURST;
	output wire sum_52_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_52_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_52_m_axi_gmem_ARPROT;
	output wire [3:0] sum_52_m_axi_gmem_ARQOS;
	output wire [3:0] sum_52_m_axi_gmem_ARREGION;
	output wire sum_52_m_axi_gmem_ARUSER;
	output wire sum_52_m_axi_gmem_RREADY;
	input sum_52_m_axi_gmem_RVALID;
	input sum_52_m_axi_gmem_RID;
	input [31:0] sum_52_m_axi_gmem_RDATA;
	input [1:0] sum_52_m_axi_gmem_RRESP;
	input sum_52_m_axi_gmem_RLAST;
	input sum_52_m_axi_gmem_RUSER;
	input sum_52_m_axi_gmem_AWREADY;
	output wire sum_52_m_axi_gmem_AWVALID;
	output wire sum_52_m_axi_gmem_AWID;
	output wire [63:0] sum_52_m_axi_gmem_AWADDR;
	output wire [7:0] sum_52_m_axi_gmem_AWLEN;
	output wire [2:0] sum_52_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_52_m_axi_gmem_AWBURST;
	output wire sum_52_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_52_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_52_m_axi_gmem_AWPROT;
	output wire [3:0] sum_52_m_axi_gmem_AWQOS;
	output wire [3:0] sum_52_m_axi_gmem_AWREGION;
	output wire sum_52_m_axi_gmem_AWUSER;
	input sum_52_m_axi_gmem_WREADY;
	output wire sum_52_m_axi_gmem_WVALID;
	output wire [31:0] sum_52_m_axi_gmem_WDATA;
	output wire [3:0] sum_52_m_axi_gmem_WSTRB;
	output wire sum_52_m_axi_gmem_WLAST;
	output wire sum_52_m_axi_gmem_WUSER;
	output wire sum_52_m_axi_gmem_BREADY;
	input sum_52_m_axi_gmem_BVALID;
	input sum_52_m_axi_gmem_BID;
	input [1:0] sum_52_m_axi_gmem_BRESP;
	input sum_52_m_axi_gmem_BUSER;
	output wire sum_52_s_axi_control_ARREADY;
	input sum_52_s_axi_control_ARVALID;
	input [4:0] sum_52_s_axi_control_ARADDR;
	input sum_52_s_axi_control_RREADY;
	output wire sum_52_s_axi_control_RVALID;
	output wire [31:0] sum_52_s_axi_control_RDATA;
	output wire [1:0] sum_52_s_axi_control_RRESP;
	output wire sum_52_s_axi_control_AWREADY;
	input sum_52_s_axi_control_AWVALID;
	input [4:0] sum_52_s_axi_control_AWADDR;
	output wire sum_52_s_axi_control_WREADY;
	input sum_52_s_axi_control_WVALID;
	input [31:0] sum_52_s_axi_control_WDATA;
	input [3:0] sum_52_s_axi_control_WSTRB;
	input sum_52_s_axi_control_BREADY;
	output wire sum_52_s_axi_control_BVALID;
	output wire [1:0] sum_52_s_axi_control_BRESP;
	input sum_53_m_axi_gmem_ARREADY;
	output wire sum_53_m_axi_gmem_ARVALID;
	output wire sum_53_m_axi_gmem_ARID;
	output wire [63:0] sum_53_m_axi_gmem_ARADDR;
	output wire [7:0] sum_53_m_axi_gmem_ARLEN;
	output wire [2:0] sum_53_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_53_m_axi_gmem_ARBURST;
	output wire sum_53_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_53_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_53_m_axi_gmem_ARPROT;
	output wire [3:0] sum_53_m_axi_gmem_ARQOS;
	output wire [3:0] sum_53_m_axi_gmem_ARREGION;
	output wire sum_53_m_axi_gmem_ARUSER;
	output wire sum_53_m_axi_gmem_RREADY;
	input sum_53_m_axi_gmem_RVALID;
	input sum_53_m_axi_gmem_RID;
	input [31:0] sum_53_m_axi_gmem_RDATA;
	input [1:0] sum_53_m_axi_gmem_RRESP;
	input sum_53_m_axi_gmem_RLAST;
	input sum_53_m_axi_gmem_RUSER;
	input sum_53_m_axi_gmem_AWREADY;
	output wire sum_53_m_axi_gmem_AWVALID;
	output wire sum_53_m_axi_gmem_AWID;
	output wire [63:0] sum_53_m_axi_gmem_AWADDR;
	output wire [7:0] sum_53_m_axi_gmem_AWLEN;
	output wire [2:0] sum_53_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_53_m_axi_gmem_AWBURST;
	output wire sum_53_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_53_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_53_m_axi_gmem_AWPROT;
	output wire [3:0] sum_53_m_axi_gmem_AWQOS;
	output wire [3:0] sum_53_m_axi_gmem_AWREGION;
	output wire sum_53_m_axi_gmem_AWUSER;
	input sum_53_m_axi_gmem_WREADY;
	output wire sum_53_m_axi_gmem_WVALID;
	output wire [31:0] sum_53_m_axi_gmem_WDATA;
	output wire [3:0] sum_53_m_axi_gmem_WSTRB;
	output wire sum_53_m_axi_gmem_WLAST;
	output wire sum_53_m_axi_gmem_WUSER;
	output wire sum_53_m_axi_gmem_BREADY;
	input sum_53_m_axi_gmem_BVALID;
	input sum_53_m_axi_gmem_BID;
	input [1:0] sum_53_m_axi_gmem_BRESP;
	input sum_53_m_axi_gmem_BUSER;
	output wire sum_53_s_axi_control_ARREADY;
	input sum_53_s_axi_control_ARVALID;
	input [4:0] sum_53_s_axi_control_ARADDR;
	input sum_53_s_axi_control_RREADY;
	output wire sum_53_s_axi_control_RVALID;
	output wire [31:0] sum_53_s_axi_control_RDATA;
	output wire [1:0] sum_53_s_axi_control_RRESP;
	output wire sum_53_s_axi_control_AWREADY;
	input sum_53_s_axi_control_AWVALID;
	input [4:0] sum_53_s_axi_control_AWADDR;
	output wire sum_53_s_axi_control_WREADY;
	input sum_53_s_axi_control_WVALID;
	input [31:0] sum_53_s_axi_control_WDATA;
	input [3:0] sum_53_s_axi_control_WSTRB;
	input sum_53_s_axi_control_BREADY;
	output wire sum_53_s_axi_control_BVALID;
	output wire [1:0] sum_53_s_axi_control_BRESP;
	input sum_54_m_axi_gmem_ARREADY;
	output wire sum_54_m_axi_gmem_ARVALID;
	output wire sum_54_m_axi_gmem_ARID;
	output wire [63:0] sum_54_m_axi_gmem_ARADDR;
	output wire [7:0] sum_54_m_axi_gmem_ARLEN;
	output wire [2:0] sum_54_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_54_m_axi_gmem_ARBURST;
	output wire sum_54_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_54_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_54_m_axi_gmem_ARPROT;
	output wire [3:0] sum_54_m_axi_gmem_ARQOS;
	output wire [3:0] sum_54_m_axi_gmem_ARREGION;
	output wire sum_54_m_axi_gmem_ARUSER;
	output wire sum_54_m_axi_gmem_RREADY;
	input sum_54_m_axi_gmem_RVALID;
	input sum_54_m_axi_gmem_RID;
	input [31:0] sum_54_m_axi_gmem_RDATA;
	input [1:0] sum_54_m_axi_gmem_RRESP;
	input sum_54_m_axi_gmem_RLAST;
	input sum_54_m_axi_gmem_RUSER;
	input sum_54_m_axi_gmem_AWREADY;
	output wire sum_54_m_axi_gmem_AWVALID;
	output wire sum_54_m_axi_gmem_AWID;
	output wire [63:0] sum_54_m_axi_gmem_AWADDR;
	output wire [7:0] sum_54_m_axi_gmem_AWLEN;
	output wire [2:0] sum_54_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_54_m_axi_gmem_AWBURST;
	output wire sum_54_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_54_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_54_m_axi_gmem_AWPROT;
	output wire [3:0] sum_54_m_axi_gmem_AWQOS;
	output wire [3:0] sum_54_m_axi_gmem_AWREGION;
	output wire sum_54_m_axi_gmem_AWUSER;
	input sum_54_m_axi_gmem_WREADY;
	output wire sum_54_m_axi_gmem_WVALID;
	output wire [31:0] sum_54_m_axi_gmem_WDATA;
	output wire [3:0] sum_54_m_axi_gmem_WSTRB;
	output wire sum_54_m_axi_gmem_WLAST;
	output wire sum_54_m_axi_gmem_WUSER;
	output wire sum_54_m_axi_gmem_BREADY;
	input sum_54_m_axi_gmem_BVALID;
	input sum_54_m_axi_gmem_BID;
	input [1:0] sum_54_m_axi_gmem_BRESP;
	input sum_54_m_axi_gmem_BUSER;
	output wire sum_54_s_axi_control_ARREADY;
	input sum_54_s_axi_control_ARVALID;
	input [4:0] sum_54_s_axi_control_ARADDR;
	input sum_54_s_axi_control_RREADY;
	output wire sum_54_s_axi_control_RVALID;
	output wire [31:0] sum_54_s_axi_control_RDATA;
	output wire [1:0] sum_54_s_axi_control_RRESP;
	output wire sum_54_s_axi_control_AWREADY;
	input sum_54_s_axi_control_AWVALID;
	input [4:0] sum_54_s_axi_control_AWADDR;
	output wire sum_54_s_axi_control_WREADY;
	input sum_54_s_axi_control_WVALID;
	input [31:0] sum_54_s_axi_control_WDATA;
	input [3:0] sum_54_s_axi_control_WSTRB;
	input sum_54_s_axi_control_BREADY;
	output wire sum_54_s_axi_control_BVALID;
	output wire [1:0] sum_54_s_axi_control_BRESP;
	input sum_55_m_axi_gmem_ARREADY;
	output wire sum_55_m_axi_gmem_ARVALID;
	output wire sum_55_m_axi_gmem_ARID;
	output wire [63:0] sum_55_m_axi_gmem_ARADDR;
	output wire [7:0] sum_55_m_axi_gmem_ARLEN;
	output wire [2:0] sum_55_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_55_m_axi_gmem_ARBURST;
	output wire sum_55_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_55_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_55_m_axi_gmem_ARPROT;
	output wire [3:0] sum_55_m_axi_gmem_ARQOS;
	output wire [3:0] sum_55_m_axi_gmem_ARREGION;
	output wire sum_55_m_axi_gmem_ARUSER;
	output wire sum_55_m_axi_gmem_RREADY;
	input sum_55_m_axi_gmem_RVALID;
	input sum_55_m_axi_gmem_RID;
	input [31:0] sum_55_m_axi_gmem_RDATA;
	input [1:0] sum_55_m_axi_gmem_RRESP;
	input sum_55_m_axi_gmem_RLAST;
	input sum_55_m_axi_gmem_RUSER;
	input sum_55_m_axi_gmem_AWREADY;
	output wire sum_55_m_axi_gmem_AWVALID;
	output wire sum_55_m_axi_gmem_AWID;
	output wire [63:0] sum_55_m_axi_gmem_AWADDR;
	output wire [7:0] sum_55_m_axi_gmem_AWLEN;
	output wire [2:0] sum_55_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_55_m_axi_gmem_AWBURST;
	output wire sum_55_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_55_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_55_m_axi_gmem_AWPROT;
	output wire [3:0] sum_55_m_axi_gmem_AWQOS;
	output wire [3:0] sum_55_m_axi_gmem_AWREGION;
	output wire sum_55_m_axi_gmem_AWUSER;
	input sum_55_m_axi_gmem_WREADY;
	output wire sum_55_m_axi_gmem_WVALID;
	output wire [31:0] sum_55_m_axi_gmem_WDATA;
	output wire [3:0] sum_55_m_axi_gmem_WSTRB;
	output wire sum_55_m_axi_gmem_WLAST;
	output wire sum_55_m_axi_gmem_WUSER;
	output wire sum_55_m_axi_gmem_BREADY;
	input sum_55_m_axi_gmem_BVALID;
	input sum_55_m_axi_gmem_BID;
	input [1:0] sum_55_m_axi_gmem_BRESP;
	input sum_55_m_axi_gmem_BUSER;
	output wire sum_55_s_axi_control_ARREADY;
	input sum_55_s_axi_control_ARVALID;
	input [4:0] sum_55_s_axi_control_ARADDR;
	input sum_55_s_axi_control_RREADY;
	output wire sum_55_s_axi_control_RVALID;
	output wire [31:0] sum_55_s_axi_control_RDATA;
	output wire [1:0] sum_55_s_axi_control_RRESP;
	output wire sum_55_s_axi_control_AWREADY;
	input sum_55_s_axi_control_AWVALID;
	input [4:0] sum_55_s_axi_control_AWADDR;
	output wire sum_55_s_axi_control_WREADY;
	input sum_55_s_axi_control_WVALID;
	input [31:0] sum_55_s_axi_control_WDATA;
	input [3:0] sum_55_s_axi_control_WSTRB;
	input sum_55_s_axi_control_BREADY;
	output wire sum_55_s_axi_control_BVALID;
	output wire [1:0] sum_55_s_axi_control_BRESP;
	input sum_56_m_axi_gmem_ARREADY;
	output wire sum_56_m_axi_gmem_ARVALID;
	output wire sum_56_m_axi_gmem_ARID;
	output wire [63:0] sum_56_m_axi_gmem_ARADDR;
	output wire [7:0] sum_56_m_axi_gmem_ARLEN;
	output wire [2:0] sum_56_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_56_m_axi_gmem_ARBURST;
	output wire sum_56_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_56_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_56_m_axi_gmem_ARPROT;
	output wire [3:0] sum_56_m_axi_gmem_ARQOS;
	output wire [3:0] sum_56_m_axi_gmem_ARREGION;
	output wire sum_56_m_axi_gmem_ARUSER;
	output wire sum_56_m_axi_gmem_RREADY;
	input sum_56_m_axi_gmem_RVALID;
	input sum_56_m_axi_gmem_RID;
	input [31:0] sum_56_m_axi_gmem_RDATA;
	input [1:0] sum_56_m_axi_gmem_RRESP;
	input sum_56_m_axi_gmem_RLAST;
	input sum_56_m_axi_gmem_RUSER;
	input sum_56_m_axi_gmem_AWREADY;
	output wire sum_56_m_axi_gmem_AWVALID;
	output wire sum_56_m_axi_gmem_AWID;
	output wire [63:0] sum_56_m_axi_gmem_AWADDR;
	output wire [7:0] sum_56_m_axi_gmem_AWLEN;
	output wire [2:0] sum_56_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_56_m_axi_gmem_AWBURST;
	output wire sum_56_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_56_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_56_m_axi_gmem_AWPROT;
	output wire [3:0] sum_56_m_axi_gmem_AWQOS;
	output wire [3:0] sum_56_m_axi_gmem_AWREGION;
	output wire sum_56_m_axi_gmem_AWUSER;
	input sum_56_m_axi_gmem_WREADY;
	output wire sum_56_m_axi_gmem_WVALID;
	output wire [31:0] sum_56_m_axi_gmem_WDATA;
	output wire [3:0] sum_56_m_axi_gmem_WSTRB;
	output wire sum_56_m_axi_gmem_WLAST;
	output wire sum_56_m_axi_gmem_WUSER;
	output wire sum_56_m_axi_gmem_BREADY;
	input sum_56_m_axi_gmem_BVALID;
	input sum_56_m_axi_gmem_BID;
	input [1:0] sum_56_m_axi_gmem_BRESP;
	input sum_56_m_axi_gmem_BUSER;
	output wire sum_56_s_axi_control_ARREADY;
	input sum_56_s_axi_control_ARVALID;
	input [4:0] sum_56_s_axi_control_ARADDR;
	input sum_56_s_axi_control_RREADY;
	output wire sum_56_s_axi_control_RVALID;
	output wire [31:0] sum_56_s_axi_control_RDATA;
	output wire [1:0] sum_56_s_axi_control_RRESP;
	output wire sum_56_s_axi_control_AWREADY;
	input sum_56_s_axi_control_AWVALID;
	input [4:0] sum_56_s_axi_control_AWADDR;
	output wire sum_56_s_axi_control_WREADY;
	input sum_56_s_axi_control_WVALID;
	input [31:0] sum_56_s_axi_control_WDATA;
	input [3:0] sum_56_s_axi_control_WSTRB;
	input sum_56_s_axi_control_BREADY;
	output wire sum_56_s_axi_control_BVALID;
	output wire [1:0] sum_56_s_axi_control_BRESP;
	input sum_57_m_axi_gmem_ARREADY;
	output wire sum_57_m_axi_gmem_ARVALID;
	output wire sum_57_m_axi_gmem_ARID;
	output wire [63:0] sum_57_m_axi_gmem_ARADDR;
	output wire [7:0] sum_57_m_axi_gmem_ARLEN;
	output wire [2:0] sum_57_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_57_m_axi_gmem_ARBURST;
	output wire sum_57_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_57_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_57_m_axi_gmem_ARPROT;
	output wire [3:0] sum_57_m_axi_gmem_ARQOS;
	output wire [3:0] sum_57_m_axi_gmem_ARREGION;
	output wire sum_57_m_axi_gmem_ARUSER;
	output wire sum_57_m_axi_gmem_RREADY;
	input sum_57_m_axi_gmem_RVALID;
	input sum_57_m_axi_gmem_RID;
	input [31:0] sum_57_m_axi_gmem_RDATA;
	input [1:0] sum_57_m_axi_gmem_RRESP;
	input sum_57_m_axi_gmem_RLAST;
	input sum_57_m_axi_gmem_RUSER;
	input sum_57_m_axi_gmem_AWREADY;
	output wire sum_57_m_axi_gmem_AWVALID;
	output wire sum_57_m_axi_gmem_AWID;
	output wire [63:0] sum_57_m_axi_gmem_AWADDR;
	output wire [7:0] sum_57_m_axi_gmem_AWLEN;
	output wire [2:0] sum_57_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_57_m_axi_gmem_AWBURST;
	output wire sum_57_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_57_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_57_m_axi_gmem_AWPROT;
	output wire [3:0] sum_57_m_axi_gmem_AWQOS;
	output wire [3:0] sum_57_m_axi_gmem_AWREGION;
	output wire sum_57_m_axi_gmem_AWUSER;
	input sum_57_m_axi_gmem_WREADY;
	output wire sum_57_m_axi_gmem_WVALID;
	output wire [31:0] sum_57_m_axi_gmem_WDATA;
	output wire [3:0] sum_57_m_axi_gmem_WSTRB;
	output wire sum_57_m_axi_gmem_WLAST;
	output wire sum_57_m_axi_gmem_WUSER;
	output wire sum_57_m_axi_gmem_BREADY;
	input sum_57_m_axi_gmem_BVALID;
	input sum_57_m_axi_gmem_BID;
	input [1:0] sum_57_m_axi_gmem_BRESP;
	input sum_57_m_axi_gmem_BUSER;
	output wire sum_57_s_axi_control_ARREADY;
	input sum_57_s_axi_control_ARVALID;
	input [4:0] sum_57_s_axi_control_ARADDR;
	input sum_57_s_axi_control_RREADY;
	output wire sum_57_s_axi_control_RVALID;
	output wire [31:0] sum_57_s_axi_control_RDATA;
	output wire [1:0] sum_57_s_axi_control_RRESP;
	output wire sum_57_s_axi_control_AWREADY;
	input sum_57_s_axi_control_AWVALID;
	input [4:0] sum_57_s_axi_control_AWADDR;
	output wire sum_57_s_axi_control_WREADY;
	input sum_57_s_axi_control_WVALID;
	input [31:0] sum_57_s_axi_control_WDATA;
	input [3:0] sum_57_s_axi_control_WSTRB;
	input sum_57_s_axi_control_BREADY;
	output wire sum_57_s_axi_control_BVALID;
	output wire [1:0] sum_57_s_axi_control_BRESP;
	input sum_58_m_axi_gmem_ARREADY;
	output wire sum_58_m_axi_gmem_ARVALID;
	output wire sum_58_m_axi_gmem_ARID;
	output wire [63:0] sum_58_m_axi_gmem_ARADDR;
	output wire [7:0] sum_58_m_axi_gmem_ARLEN;
	output wire [2:0] sum_58_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_58_m_axi_gmem_ARBURST;
	output wire sum_58_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_58_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_58_m_axi_gmem_ARPROT;
	output wire [3:0] sum_58_m_axi_gmem_ARQOS;
	output wire [3:0] sum_58_m_axi_gmem_ARREGION;
	output wire sum_58_m_axi_gmem_ARUSER;
	output wire sum_58_m_axi_gmem_RREADY;
	input sum_58_m_axi_gmem_RVALID;
	input sum_58_m_axi_gmem_RID;
	input [31:0] sum_58_m_axi_gmem_RDATA;
	input [1:0] sum_58_m_axi_gmem_RRESP;
	input sum_58_m_axi_gmem_RLAST;
	input sum_58_m_axi_gmem_RUSER;
	input sum_58_m_axi_gmem_AWREADY;
	output wire sum_58_m_axi_gmem_AWVALID;
	output wire sum_58_m_axi_gmem_AWID;
	output wire [63:0] sum_58_m_axi_gmem_AWADDR;
	output wire [7:0] sum_58_m_axi_gmem_AWLEN;
	output wire [2:0] sum_58_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_58_m_axi_gmem_AWBURST;
	output wire sum_58_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_58_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_58_m_axi_gmem_AWPROT;
	output wire [3:0] sum_58_m_axi_gmem_AWQOS;
	output wire [3:0] sum_58_m_axi_gmem_AWREGION;
	output wire sum_58_m_axi_gmem_AWUSER;
	input sum_58_m_axi_gmem_WREADY;
	output wire sum_58_m_axi_gmem_WVALID;
	output wire [31:0] sum_58_m_axi_gmem_WDATA;
	output wire [3:0] sum_58_m_axi_gmem_WSTRB;
	output wire sum_58_m_axi_gmem_WLAST;
	output wire sum_58_m_axi_gmem_WUSER;
	output wire sum_58_m_axi_gmem_BREADY;
	input sum_58_m_axi_gmem_BVALID;
	input sum_58_m_axi_gmem_BID;
	input [1:0] sum_58_m_axi_gmem_BRESP;
	input sum_58_m_axi_gmem_BUSER;
	output wire sum_58_s_axi_control_ARREADY;
	input sum_58_s_axi_control_ARVALID;
	input [4:0] sum_58_s_axi_control_ARADDR;
	input sum_58_s_axi_control_RREADY;
	output wire sum_58_s_axi_control_RVALID;
	output wire [31:0] sum_58_s_axi_control_RDATA;
	output wire [1:0] sum_58_s_axi_control_RRESP;
	output wire sum_58_s_axi_control_AWREADY;
	input sum_58_s_axi_control_AWVALID;
	input [4:0] sum_58_s_axi_control_AWADDR;
	output wire sum_58_s_axi_control_WREADY;
	input sum_58_s_axi_control_WVALID;
	input [31:0] sum_58_s_axi_control_WDATA;
	input [3:0] sum_58_s_axi_control_WSTRB;
	input sum_58_s_axi_control_BREADY;
	output wire sum_58_s_axi_control_BVALID;
	output wire [1:0] sum_58_s_axi_control_BRESP;
	input sum_59_m_axi_gmem_ARREADY;
	output wire sum_59_m_axi_gmem_ARVALID;
	output wire sum_59_m_axi_gmem_ARID;
	output wire [63:0] sum_59_m_axi_gmem_ARADDR;
	output wire [7:0] sum_59_m_axi_gmem_ARLEN;
	output wire [2:0] sum_59_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_59_m_axi_gmem_ARBURST;
	output wire sum_59_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_59_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_59_m_axi_gmem_ARPROT;
	output wire [3:0] sum_59_m_axi_gmem_ARQOS;
	output wire [3:0] sum_59_m_axi_gmem_ARREGION;
	output wire sum_59_m_axi_gmem_ARUSER;
	output wire sum_59_m_axi_gmem_RREADY;
	input sum_59_m_axi_gmem_RVALID;
	input sum_59_m_axi_gmem_RID;
	input [31:0] sum_59_m_axi_gmem_RDATA;
	input [1:0] sum_59_m_axi_gmem_RRESP;
	input sum_59_m_axi_gmem_RLAST;
	input sum_59_m_axi_gmem_RUSER;
	input sum_59_m_axi_gmem_AWREADY;
	output wire sum_59_m_axi_gmem_AWVALID;
	output wire sum_59_m_axi_gmem_AWID;
	output wire [63:0] sum_59_m_axi_gmem_AWADDR;
	output wire [7:0] sum_59_m_axi_gmem_AWLEN;
	output wire [2:0] sum_59_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_59_m_axi_gmem_AWBURST;
	output wire sum_59_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_59_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_59_m_axi_gmem_AWPROT;
	output wire [3:0] sum_59_m_axi_gmem_AWQOS;
	output wire [3:0] sum_59_m_axi_gmem_AWREGION;
	output wire sum_59_m_axi_gmem_AWUSER;
	input sum_59_m_axi_gmem_WREADY;
	output wire sum_59_m_axi_gmem_WVALID;
	output wire [31:0] sum_59_m_axi_gmem_WDATA;
	output wire [3:0] sum_59_m_axi_gmem_WSTRB;
	output wire sum_59_m_axi_gmem_WLAST;
	output wire sum_59_m_axi_gmem_WUSER;
	output wire sum_59_m_axi_gmem_BREADY;
	input sum_59_m_axi_gmem_BVALID;
	input sum_59_m_axi_gmem_BID;
	input [1:0] sum_59_m_axi_gmem_BRESP;
	input sum_59_m_axi_gmem_BUSER;
	output wire sum_59_s_axi_control_ARREADY;
	input sum_59_s_axi_control_ARVALID;
	input [4:0] sum_59_s_axi_control_ARADDR;
	input sum_59_s_axi_control_RREADY;
	output wire sum_59_s_axi_control_RVALID;
	output wire [31:0] sum_59_s_axi_control_RDATA;
	output wire [1:0] sum_59_s_axi_control_RRESP;
	output wire sum_59_s_axi_control_AWREADY;
	input sum_59_s_axi_control_AWVALID;
	input [4:0] sum_59_s_axi_control_AWADDR;
	output wire sum_59_s_axi_control_WREADY;
	input sum_59_s_axi_control_WVALID;
	input [31:0] sum_59_s_axi_control_WDATA;
	input [3:0] sum_59_s_axi_control_WSTRB;
	input sum_59_s_axi_control_BREADY;
	output wire sum_59_s_axi_control_BVALID;
	output wire [1:0] sum_59_s_axi_control_BRESP;
	input sum_60_m_axi_gmem_ARREADY;
	output wire sum_60_m_axi_gmem_ARVALID;
	output wire sum_60_m_axi_gmem_ARID;
	output wire [63:0] sum_60_m_axi_gmem_ARADDR;
	output wire [7:0] sum_60_m_axi_gmem_ARLEN;
	output wire [2:0] sum_60_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_60_m_axi_gmem_ARBURST;
	output wire sum_60_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_60_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_60_m_axi_gmem_ARPROT;
	output wire [3:0] sum_60_m_axi_gmem_ARQOS;
	output wire [3:0] sum_60_m_axi_gmem_ARREGION;
	output wire sum_60_m_axi_gmem_ARUSER;
	output wire sum_60_m_axi_gmem_RREADY;
	input sum_60_m_axi_gmem_RVALID;
	input sum_60_m_axi_gmem_RID;
	input [31:0] sum_60_m_axi_gmem_RDATA;
	input [1:0] sum_60_m_axi_gmem_RRESP;
	input sum_60_m_axi_gmem_RLAST;
	input sum_60_m_axi_gmem_RUSER;
	input sum_60_m_axi_gmem_AWREADY;
	output wire sum_60_m_axi_gmem_AWVALID;
	output wire sum_60_m_axi_gmem_AWID;
	output wire [63:0] sum_60_m_axi_gmem_AWADDR;
	output wire [7:0] sum_60_m_axi_gmem_AWLEN;
	output wire [2:0] sum_60_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_60_m_axi_gmem_AWBURST;
	output wire sum_60_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_60_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_60_m_axi_gmem_AWPROT;
	output wire [3:0] sum_60_m_axi_gmem_AWQOS;
	output wire [3:0] sum_60_m_axi_gmem_AWREGION;
	output wire sum_60_m_axi_gmem_AWUSER;
	input sum_60_m_axi_gmem_WREADY;
	output wire sum_60_m_axi_gmem_WVALID;
	output wire [31:0] sum_60_m_axi_gmem_WDATA;
	output wire [3:0] sum_60_m_axi_gmem_WSTRB;
	output wire sum_60_m_axi_gmem_WLAST;
	output wire sum_60_m_axi_gmem_WUSER;
	output wire sum_60_m_axi_gmem_BREADY;
	input sum_60_m_axi_gmem_BVALID;
	input sum_60_m_axi_gmem_BID;
	input [1:0] sum_60_m_axi_gmem_BRESP;
	input sum_60_m_axi_gmem_BUSER;
	output wire sum_60_s_axi_control_ARREADY;
	input sum_60_s_axi_control_ARVALID;
	input [4:0] sum_60_s_axi_control_ARADDR;
	input sum_60_s_axi_control_RREADY;
	output wire sum_60_s_axi_control_RVALID;
	output wire [31:0] sum_60_s_axi_control_RDATA;
	output wire [1:0] sum_60_s_axi_control_RRESP;
	output wire sum_60_s_axi_control_AWREADY;
	input sum_60_s_axi_control_AWVALID;
	input [4:0] sum_60_s_axi_control_AWADDR;
	output wire sum_60_s_axi_control_WREADY;
	input sum_60_s_axi_control_WVALID;
	input [31:0] sum_60_s_axi_control_WDATA;
	input [3:0] sum_60_s_axi_control_WSTRB;
	input sum_60_s_axi_control_BREADY;
	output wire sum_60_s_axi_control_BVALID;
	output wire [1:0] sum_60_s_axi_control_BRESP;
	input sum_61_m_axi_gmem_ARREADY;
	output wire sum_61_m_axi_gmem_ARVALID;
	output wire sum_61_m_axi_gmem_ARID;
	output wire [63:0] sum_61_m_axi_gmem_ARADDR;
	output wire [7:0] sum_61_m_axi_gmem_ARLEN;
	output wire [2:0] sum_61_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_61_m_axi_gmem_ARBURST;
	output wire sum_61_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_61_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_61_m_axi_gmem_ARPROT;
	output wire [3:0] sum_61_m_axi_gmem_ARQOS;
	output wire [3:0] sum_61_m_axi_gmem_ARREGION;
	output wire sum_61_m_axi_gmem_ARUSER;
	output wire sum_61_m_axi_gmem_RREADY;
	input sum_61_m_axi_gmem_RVALID;
	input sum_61_m_axi_gmem_RID;
	input [31:0] sum_61_m_axi_gmem_RDATA;
	input [1:0] sum_61_m_axi_gmem_RRESP;
	input sum_61_m_axi_gmem_RLAST;
	input sum_61_m_axi_gmem_RUSER;
	input sum_61_m_axi_gmem_AWREADY;
	output wire sum_61_m_axi_gmem_AWVALID;
	output wire sum_61_m_axi_gmem_AWID;
	output wire [63:0] sum_61_m_axi_gmem_AWADDR;
	output wire [7:0] sum_61_m_axi_gmem_AWLEN;
	output wire [2:0] sum_61_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_61_m_axi_gmem_AWBURST;
	output wire sum_61_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_61_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_61_m_axi_gmem_AWPROT;
	output wire [3:0] sum_61_m_axi_gmem_AWQOS;
	output wire [3:0] sum_61_m_axi_gmem_AWREGION;
	output wire sum_61_m_axi_gmem_AWUSER;
	input sum_61_m_axi_gmem_WREADY;
	output wire sum_61_m_axi_gmem_WVALID;
	output wire [31:0] sum_61_m_axi_gmem_WDATA;
	output wire [3:0] sum_61_m_axi_gmem_WSTRB;
	output wire sum_61_m_axi_gmem_WLAST;
	output wire sum_61_m_axi_gmem_WUSER;
	output wire sum_61_m_axi_gmem_BREADY;
	input sum_61_m_axi_gmem_BVALID;
	input sum_61_m_axi_gmem_BID;
	input [1:0] sum_61_m_axi_gmem_BRESP;
	input sum_61_m_axi_gmem_BUSER;
	output wire sum_61_s_axi_control_ARREADY;
	input sum_61_s_axi_control_ARVALID;
	input [4:0] sum_61_s_axi_control_ARADDR;
	input sum_61_s_axi_control_RREADY;
	output wire sum_61_s_axi_control_RVALID;
	output wire [31:0] sum_61_s_axi_control_RDATA;
	output wire [1:0] sum_61_s_axi_control_RRESP;
	output wire sum_61_s_axi_control_AWREADY;
	input sum_61_s_axi_control_AWVALID;
	input [4:0] sum_61_s_axi_control_AWADDR;
	output wire sum_61_s_axi_control_WREADY;
	input sum_61_s_axi_control_WVALID;
	input [31:0] sum_61_s_axi_control_WDATA;
	input [3:0] sum_61_s_axi_control_WSTRB;
	input sum_61_s_axi_control_BREADY;
	output wire sum_61_s_axi_control_BVALID;
	output wire [1:0] sum_61_s_axi_control_BRESP;
	input sum_62_m_axi_gmem_ARREADY;
	output wire sum_62_m_axi_gmem_ARVALID;
	output wire sum_62_m_axi_gmem_ARID;
	output wire [63:0] sum_62_m_axi_gmem_ARADDR;
	output wire [7:0] sum_62_m_axi_gmem_ARLEN;
	output wire [2:0] sum_62_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_62_m_axi_gmem_ARBURST;
	output wire sum_62_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_62_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_62_m_axi_gmem_ARPROT;
	output wire [3:0] sum_62_m_axi_gmem_ARQOS;
	output wire [3:0] sum_62_m_axi_gmem_ARREGION;
	output wire sum_62_m_axi_gmem_ARUSER;
	output wire sum_62_m_axi_gmem_RREADY;
	input sum_62_m_axi_gmem_RVALID;
	input sum_62_m_axi_gmem_RID;
	input [31:0] sum_62_m_axi_gmem_RDATA;
	input [1:0] sum_62_m_axi_gmem_RRESP;
	input sum_62_m_axi_gmem_RLAST;
	input sum_62_m_axi_gmem_RUSER;
	input sum_62_m_axi_gmem_AWREADY;
	output wire sum_62_m_axi_gmem_AWVALID;
	output wire sum_62_m_axi_gmem_AWID;
	output wire [63:0] sum_62_m_axi_gmem_AWADDR;
	output wire [7:0] sum_62_m_axi_gmem_AWLEN;
	output wire [2:0] sum_62_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_62_m_axi_gmem_AWBURST;
	output wire sum_62_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_62_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_62_m_axi_gmem_AWPROT;
	output wire [3:0] sum_62_m_axi_gmem_AWQOS;
	output wire [3:0] sum_62_m_axi_gmem_AWREGION;
	output wire sum_62_m_axi_gmem_AWUSER;
	input sum_62_m_axi_gmem_WREADY;
	output wire sum_62_m_axi_gmem_WVALID;
	output wire [31:0] sum_62_m_axi_gmem_WDATA;
	output wire [3:0] sum_62_m_axi_gmem_WSTRB;
	output wire sum_62_m_axi_gmem_WLAST;
	output wire sum_62_m_axi_gmem_WUSER;
	output wire sum_62_m_axi_gmem_BREADY;
	input sum_62_m_axi_gmem_BVALID;
	input sum_62_m_axi_gmem_BID;
	input [1:0] sum_62_m_axi_gmem_BRESP;
	input sum_62_m_axi_gmem_BUSER;
	output wire sum_62_s_axi_control_ARREADY;
	input sum_62_s_axi_control_ARVALID;
	input [4:0] sum_62_s_axi_control_ARADDR;
	input sum_62_s_axi_control_RREADY;
	output wire sum_62_s_axi_control_RVALID;
	output wire [31:0] sum_62_s_axi_control_RDATA;
	output wire [1:0] sum_62_s_axi_control_RRESP;
	output wire sum_62_s_axi_control_AWREADY;
	input sum_62_s_axi_control_AWVALID;
	input [4:0] sum_62_s_axi_control_AWADDR;
	output wire sum_62_s_axi_control_WREADY;
	input sum_62_s_axi_control_WVALID;
	input [31:0] sum_62_s_axi_control_WDATA;
	input [3:0] sum_62_s_axi_control_WSTRB;
	input sum_62_s_axi_control_BREADY;
	output wire sum_62_s_axi_control_BVALID;
	output wire [1:0] sum_62_s_axi_control_BRESP;
	input sum_63_m_axi_gmem_ARREADY;
	output wire sum_63_m_axi_gmem_ARVALID;
	output wire sum_63_m_axi_gmem_ARID;
	output wire [63:0] sum_63_m_axi_gmem_ARADDR;
	output wire [7:0] sum_63_m_axi_gmem_ARLEN;
	output wire [2:0] sum_63_m_axi_gmem_ARSIZE;
	output wire [1:0] sum_63_m_axi_gmem_ARBURST;
	output wire sum_63_m_axi_gmem_ARLOCK;
	output wire [3:0] sum_63_m_axi_gmem_ARCACHE;
	output wire [2:0] sum_63_m_axi_gmem_ARPROT;
	output wire [3:0] sum_63_m_axi_gmem_ARQOS;
	output wire [3:0] sum_63_m_axi_gmem_ARREGION;
	output wire sum_63_m_axi_gmem_ARUSER;
	output wire sum_63_m_axi_gmem_RREADY;
	input sum_63_m_axi_gmem_RVALID;
	input sum_63_m_axi_gmem_RID;
	input [31:0] sum_63_m_axi_gmem_RDATA;
	input [1:0] sum_63_m_axi_gmem_RRESP;
	input sum_63_m_axi_gmem_RLAST;
	input sum_63_m_axi_gmem_RUSER;
	input sum_63_m_axi_gmem_AWREADY;
	output wire sum_63_m_axi_gmem_AWVALID;
	output wire sum_63_m_axi_gmem_AWID;
	output wire [63:0] sum_63_m_axi_gmem_AWADDR;
	output wire [7:0] sum_63_m_axi_gmem_AWLEN;
	output wire [2:0] sum_63_m_axi_gmem_AWSIZE;
	output wire [1:0] sum_63_m_axi_gmem_AWBURST;
	output wire sum_63_m_axi_gmem_AWLOCK;
	output wire [3:0] sum_63_m_axi_gmem_AWCACHE;
	output wire [2:0] sum_63_m_axi_gmem_AWPROT;
	output wire [3:0] sum_63_m_axi_gmem_AWQOS;
	output wire [3:0] sum_63_m_axi_gmem_AWREGION;
	output wire sum_63_m_axi_gmem_AWUSER;
	input sum_63_m_axi_gmem_WREADY;
	output wire sum_63_m_axi_gmem_WVALID;
	output wire [31:0] sum_63_m_axi_gmem_WDATA;
	output wire [3:0] sum_63_m_axi_gmem_WSTRB;
	output wire sum_63_m_axi_gmem_WLAST;
	output wire sum_63_m_axi_gmem_WUSER;
	output wire sum_63_m_axi_gmem_BREADY;
	input sum_63_m_axi_gmem_BVALID;
	input sum_63_m_axi_gmem_BID;
	input [1:0] sum_63_m_axi_gmem_BRESP;
	input sum_63_m_axi_gmem_BUSER;
	output wire sum_63_s_axi_control_ARREADY;
	input sum_63_s_axi_control_ARVALID;
	input [4:0] sum_63_s_axi_control_ARADDR;
	input sum_63_s_axi_control_RREADY;
	output wire sum_63_s_axi_control_RVALID;
	output wire [31:0] sum_63_s_axi_control_RDATA;
	output wire [1:0] sum_63_s_axi_control_RRESP;
	output wire sum_63_s_axi_control_AWREADY;
	input sum_63_s_axi_control_AWVALID;
	input [4:0] sum_63_s_axi_control_AWADDR;
	output wire sum_63_s_axi_control_WREADY;
	input sum_63_s_axi_control_WVALID;
	input [31:0] sum_63_s_axi_control_WDATA;
	input [3:0] sum_63_s_axi_control_WSTRB;
	input sum_63_s_axi_control_BREADY;
	output wire sum_63_s_axi_control_BVALID;
	output wire [1:0] sum_63_s_axi_control_BRESP;
	input sum_schedulerAXI_0_ARREADY;
	output wire sum_schedulerAXI_0_ARVALID;
	output wire [1:0] sum_schedulerAXI_0_ARID;
	output wire [63:0] sum_schedulerAXI_0_ARADDR;
	output wire [7:0] sum_schedulerAXI_0_ARLEN;
	output wire [2:0] sum_schedulerAXI_0_ARSIZE;
	output wire [1:0] sum_schedulerAXI_0_ARBURST;
	output wire sum_schedulerAXI_0_ARLOCK;
	output wire [3:0] sum_schedulerAXI_0_ARCACHE;
	output wire [2:0] sum_schedulerAXI_0_ARPROT;
	output wire [3:0] sum_schedulerAXI_0_ARQOS;
	output wire [3:0] sum_schedulerAXI_0_ARREGION;
	output wire sum_schedulerAXI_0_RREADY;
	input sum_schedulerAXI_0_RVALID;
	input [1:0] sum_schedulerAXI_0_RID;
	input [255:0] sum_schedulerAXI_0_RDATA;
	input [1:0] sum_schedulerAXI_0_RRESP;
	input sum_schedulerAXI_0_RLAST;
	input sum_schedulerAXI_0_AWREADY;
	output wire sum_schedulerAXI_0_AWVALID;
	output wire [1:0] sum_schedulerAXI_0_AWID;
	output wire [63:0] sum_schedulerAXI_0_AWADDR;
	output wire [7:0] sum_schedulerAXI_0_AWLEN;
	output wire [2:0] sum_schedulerAXI_0_AWSIZE;
	output wire [1:0] sum_schedulerAXI_0_AWBURST;
	output wire sum_schedulerAXI_0_AWLOCK;
	output wire [3:0] sum_schedulerAXI_0_AWCACHE;
	output wire [2:0] sum_schedulerAXI_0_AWPROT;
	output wire [3:0] sum_schedulerAXI_0_AWQOS;
	output wire [3:0] sum_schedulerAXI_0_AWREGION;
	input sum_schedulerAXI_0_WREADY;
	output wire sum_schedulerAXI_0_WVALID;
	output wire [255:0] sum_schedulerAXI_0_WDATA;
	output wire [31:0] sum_schedulerAXI_0_WSTRB;
	output wire sum_schedulerAXI_0_WLAST;
	output wire sum_schedulerAXI_0_BREADY;
	input sum_schedulerAXI_0_BVALID;
	input [1:0] sum_schedulerAXI_0_BID;
	input [1:0] sum_schedulerAXI_0_BRESP;
	input sum_closureAllocatorAXI_0_ARREADY;
	output wire sum_closureAllocatorAXI_0_ARVALID;
	output wire [6:0] sum_closureAllocatorAXI_0_ARID;
	output wire [63:0] sum_closureAllocatorAXI_0_ARADDR;
	output wire [7:0] sum_closureAllocatorAXI_0_ARLEN;
	output wire [2:0] sum_closureAllocatorAXI_0_ARSIZE;
	output wire [1:0] sum_closureAllocatorAXI_0_ARBURST;
	output wire sum_closureAllocatorAXI_0_ARLOCK;
	output wire [3:0] sum_closureAllocatorAXI_0_ARCACHE;
	output wire [2:0] sum_closureAllocatorAXI_0_ARPROT;
	output wire [3:0] sum_closureAllocatorAXI_0_ARQOS;
	output wire [3:0] sum_closureAllocatorAXI_0_ARREGION;
	output wire sum_closureAllocatorAXI_0_RREADY;
	input sum_closureAllocatorAXI_0_RVALID;
	input [6:0] sum_closureAllocatorAXI_0_RID;
	input [63:0] sum_closureAllocatorAXI_0_RDATA;
	input [1:0] sum_closureAllocatorAXI_0_RRESP;
	input sum_closureAllocatorAXI_0_RLAST;
	input sum_closureAllocatorAXI_0_AWREADY;
	output wire sum_closureAllocatorAXI_0_AWVALID;
	output wire [6:0] sum_closureAllocatorAXI_0_AWID;
	output wire [63:0] sum_closureAllocatorAXI_0_AWADDR;
	output wire [7:0] sum_closureAllocatorAXI_0_AWLEN;
	output wire [2:0] sum_closureAllocatorAXI_0_AWSIZE;
	output wire [1:0] sum_closureAllocatorAXI_0_AWBURST;
	output wire sum_closureAllocatorAXI_0_AWLOCK;
	output wire [3:0] sum_closureAllocatorAXI_0_AWCACHE;
	output wire [2:0] sum_closureAllocatorAXI_0_AWPROT;
	output wire [3:0] sum_closureAllocatorAXI_0_AWQOS;
	output wire [3:0] sum_closureAllocatorAXI_0_AWREGION;
	input sum_closureAllocatorAXI_0_WREADY;
	output wire sum_closureAllocatorAXI_0_WVALID;
	output wire [63:0] sum_closureAllocatorAXI_0_WDATA;
	output wire [7:0] sum_closureAllocatorAXI_0_WSTRB;
	output wire sum_closureAllocatorAXI_0_WLAST;
	output wire sum_closureAllocatorAXI_0_BREADY;
	input sum_closureAllocatorAXI_0_BVALID;
	input [6:0] sum_closureAllocatorAXI_0_BID;
	input [1:0] sum_closureAllocatorAXI_0_BRESP;
	input sum_argumentNotifierAXI_0_ARREADY;
	output wire sum_argumentNotifierAXI_0_ARVALID;
	output wire [4:0] sum_argumentNotifierAXI_0_ARID;
	output wire [63:0] sum_argumentNotifierAXI_0_ARADDR;
	output wire [7:0] sum_argumentNotifierAXI_0_ARLEN;
	output wire [2:0] sum_argumentNotifierAXI_0_ARSIZE;
	output wire [1:0] sum_argumentNotifierAXI_0_ARBURST;
	output wire sum_argumentNotifierAXI_0_ARLOCK;
	output wire [3:0] sum_argumentNotifierAXI_0_ARCACHE;
	output wire [2:0] sum_argumentNotifierAXI_0_ARPROT;
	output wire [3:0] sum_argumentNotifierAXI_0_ARQOS;
	output wire [3:0] sum_argumentNotifierAXI_0_ARREGION;
	output wire sum_argumentNotifierAXI_0_RREADY;
	input sum_argumentNotifierAXI_0_RVALID;
	input [4:0] sum_argumentNotifierAXI_0_RID;
	input [31:0] sum_argumentNotifierAXI_0_RDATA;
	input [1:0] sum_argumentNotifierAXI_0_RRESP;
	input sum_argumentNotifierAXI_0_RLAST;
	input sum_argumentNotifierAXI_0_AWREADY;
	output wire sum_argumentNotifierAXI_0_AWVALID;
	output wire [4:0] sum_argumentNotifierAXI_0_AWID;
	output wire [63:0] sum_argumentNotifierAXI_0_AWADDR;
	output wire [7:0] sum_argumentNotifierAXI_0_AWLEN;
	output wire [2:0] sum_argumentNotifierAXI_0_AWSIZE;
	output wire [1:0] sum_argumentNotifierAXI_0_AWBURST;
	output wire sum_argumentNotifierAXI_0_AWLOCK;
	output wire [3:0] sum_argumentNotifierAXI_0_AWCACHE;
	output wire [2:0] sum_argumentNotifierAXI_0_AWPROT;
	output wire [3:0] sum_argumentNotifierAXI_0_AWQOS;
	output wire [3:0] sum_argumentNotifierAXI_0_AWREGION;
	input sum_argumentNotifierAXI_0_WREADY;
	output wire sum_argumentNotifierAXI_0_WVALID;
	output wire [31:0] sum_argumentNotifierAXI_0_WDATA;
	output wire [3:0] sum_argumentNotifierAXI_0_WSTRB;
	output wire sum_argumentNotifierAXI_0_WLAST;
	output wire sum_argumentNotifierAXI_0_BREADY;
	input sum_argumentNotifierAXI_0_BVALID;
	input [4:0] sum_argumentNotifierAXI_0_BID;
	input [1:0] sum_argumentNotifierAXI_0_BRESP;
	wire _ArgumentNotifier_io_export_argIn_0_TREADY;
	wire _ArgumentNotifier_io_export_argIn_1_TREADY;
	wire _ArgumentNotifier_io_export_argIn_2_TREADY;
	wire _ArgumentNotifier_io_export_argIn_3_TREADY;
	wire _ArgumentNotifier_io_export_argIn_4_TREADY;
	wire _ArgumentNotifier_io_export_argIn_5_TREADY;
	wire _ArgumentNotifier_io_export_argIn_6_TREADY;
	wire _ArgumentNotifier_io_export_argIn_7_TREADY;
	wire _ArgumentNotifier_io_export_argIn_8_TREADY;
	wire _ArgumentNotifier_io_export_argIn_9_TREADY;
	wire _ArgumentNotifier_io_export_argIn_10_TREADY;
	wire _ArgumentNotifier_io_export_argIn_11_TREADY;
	wire _ArgumentNotifier_io_export_argIn_12_TREADY;
	wire _ArgumentNotifier_io_export_argIn_13_TREADY;
	wire _ArgumentNotifier_io_export_argIn_14_TREADY;
	wire _ArgumentNotifier_io_export_argIn_15_TREADY;
	wire _ArgumentNotifier_io_export_argIn_16_TREADY;
	wire _ArgumentNotifier_io_export_argIn_17_TREADY;
	wire _ArgumentNotifier_io_export_argIn_18_TREADY;
	wire _ArgumentNotifier_io_export_argIn_19_TREADY;
	wire _ArgumentNotifier_io_export_argIn_20_TREADY;
	wire _ArgumentNotifier_io_export_argIn_21_TREADY;
	wire _ArgumentNotifier_io_export_argIn_22_TREADY;
	wire _ArgumentNotifier_io_export_argIn_23_TREADY;
	wire _ArgumentNotifier_io_export_argIn_24_TREADY;
	wire _ArgumentNotifier_io_export_argIn_25_TREADY;
	wire _ArgumentNotifier_io_export_argIn_26_TREADY;
	wire _ArgumentNotifier_io_export_argIn_27_TREADY;
	wire _ArgumentNotifier_io_export_argIn_28_TREADY;
	wire _ArgumentNotifier_io_export_argIn_29_TREADY;
	wire _ArgumentNotifier_io_export_argIn_30_TREADY;
	wire _ArgumentNotifier_io_export_argIn_31_TREADY;
	wire _ArgumentNotifier_io_export_argIn_32_TREADY;
	wire _ArgumentNotifier_io_export_argIn_33_TREADY;
	wire _ArgumentNotifier_io_export_argIn_34_TREADY;
	wire _ArgumentNotifier_io_export_argIn_35_TREADY;
	wire _ArgumentNotifier_io_export_argIn_36_TREADY;
	wire _ArgumentNotifier_io_export_argIn_37_TREADY;
	wire _ArgumentNotifier_io_export_argIn_38_TREADY;
	wire _ArgumentNotifier_io_export_argIn_39_TREADY;
	wire _ArgumentNotifier_io_export_argIn_40_TREADY;
	wire _ArgumentNotifier_io_export_argIn_41_TREADY;
	wire _ArgumentNotifier_io_export_argIn_42_TREADY;
	wire _ArgumentNotifier_io_export_argIn_43_TREADY;
	wire _ArgumentNotifier_io_export_argIn_44_TREADY;
	wire _ArgumentNotifier_io_export_argIn_45_TREADY;
	wire _ArgumentNotifier_io_export_argIn_46_TREADY;
	wire _ArgumentNotifier_io_export_argIn_47_TREADY;
	wire _ArgumentNotifier_io_export_argIn_48_TREADY;
	wire _ArgumentNotifier_io_export_argIn_49_TREADY;
	wire _ArgumentNotifier_io_export_argIn_50_TREADY;
	wire _ArgumentNotifier_io_export_argIn_51_TREADY;
	wire _ArgumentNotifier_io_export_argIn_52_TREADY;
	wire _ArgumentNotifier_io_export_argIn_53_TREADY;
	wire _ArgumentNotifier_io_export_argIn_54_TREADY;
	wire _ArgumentNotifier_io_export_argIn_55_TREADY;
	wire _ArgumentNotifier_io_export_argIn_56_TREADY;
	wire _ArgumentNotifier_io_export_argIn_57_TREADY;
	wire _ArgumentNotifier_io_export_argIn_58_TREADY;
	wire _ArgumentNotifier_io_export_argIn_59_TREADY;
	wire _ArgumentNotifier_io_export_argIn_60_TREADY;
	wire _ArgumentNotifier_io_export_argIn_61_TREADY;
	wire _ArgumentNotifier_io_export_argIn_62_TREADY;
	wire _ArgumentNotifier_io_export_argIn_63_TREADY;
	wire _ArgumentNotifier_io_export_argIn_64_TREADY;
	wire _ArgumentNotifier_io_export_argIn_65_TREADY;
	wire _ArgumentNotifier_io_export_argIn_66_TREADY;
	wire _ArgumentNotifier_io_export_argIn_67_TREADY;
	wire _ArgumentNotifier_io_export_argIn_68_TREADY;
	wire _ArgumentNotifier_io_export_argIn_69_TREADY;
	wire _ArgumentNotifier_io_export_argIn_70_TREADY;
	wire _ArgumentNotifier_io_export_argIn_71_TREADY;
	wire _ArgumentNotifier_io_export_argIn_72_TREADY;
	wire _ArgumentNotifier_io_export_argIn_73_TREADY;
	wire _ArgumentNotifier_io_export_argIn_74_TREADY;
	wire _ArgumentNotifier_io_export_argIn_75_TREADY;
	wire _ArgumentNotifier_io_export_argIn_76_TREADY;
	wire _ArgumentNotifier_io_export_argIn_77_TREADY;
	wire _ArgumentNotifier_io_export_argIn_78_TREADY;
	wire _ArgumentNotifier_io_export_argIn_79_TREADY;
	wire _ArgumentNotifier_io_export_argIn_80_TREADY;
	wire _ArgumentNotifier_io_export_argIn_81_TREADY;
	wire _ArgumentNotifier_io_export_argIn_82_TREADY;
	wire _ArgumentNotifier_io_export_argIn_83_TREADY;
	wire _ArgumentNotifier_io_export_argIn_84_TREADY;
	wire _ArgumentNotifier_io_export_argIn_85_TREADY;
	wire _ArgumentNotifier_io_export_argIn_86_TREADY;
	wire _ArgumentNotifier_io_export_argIn_87_TREADY;
	wire _ArgumentNotifier_io_export_argIn_88_TREADY;
	wire _ArgumentNotifier_io_export_argIn_89_TREADY;
	wire _ArgumentNotifier_io_export_argIn_90_TREADY;
	wire _ArgumentNotifier_io_export_argIn_91_TREADY;
	wire _ArgumentNotifier_io_export_argIn_92_TREADY;
	wire _ArgumentNotifier_io_export_argIn_93_TREADY;
	wire _ArgumentNotifier_io_export_argIn_94_TREADY;
	wire _ArgumentNotifier_io_export_argIn_95_TREADY;
	wire _ArgumentNotifier_io_export_argIn_96_TREADY;
	wire _ArgumentNotifier_io_export_argIn_97_TREADY;
	wire _ArgumentNotifier_io_export_argIn_98_TREADY;
	wire _ArgumentNotifier_io_export_argIn_99_TREADY;
	wire _ArgumentNotifier_io_export_argIn_100_TREADY;
	wire _ArgumentNotifier_io_export_argIn_101_TREADY;
	wire _ArgumentNotifier_io_export_argIn_102_TREADY;
	wire _ArgumentNotifier_io_export_argIn_103_TREADY;
	wire _ArgumentNotifier_io_export_argIn_104_TREADY;
	wire _ArgumentNotifier_io_export_argIn_105_TREADY;
	wire _ArgumentNotifier_io_export_argIn_106_TREADY;
	wire _ArgumentNotifier_io_export_argIn_107_TREADY;
	wire _ArgumentNotifier_io_export_argIn_108_TREADY;
	wire _ArgumentNotifier_io_export_argIn_109_TREADY;
	wire _ArgumentNotifier_io_export_argIn_110_TREADY;
	wire _ArgumentNotifier_io_export_argIn_111_TREADY;
	wire _ArgumentNotifier_io_export_argIn_112_TREADY;
	wire _ArgumentNotifier_io_export_argIn_113_TREADY;
	wire _ArgumentNotifier_io_export_argIn_114_TREADY;
	wire _ArgumentNotifier_io_export_argIn_115_TREADY;
	wire _ArgumentNotifier_io_export_argIn_116_TREADY;
	wire _ArgumentNotifier_io_export_argIn_117_TREADY;
	wire _ArgumentNotifier_io_export_argIn_118_TREADY;
	wire _ArgumentNotifier_io_export_argIn_119_TREADY;
	wire _ArgumentNotifier_io_export_argIn_120_TREADY;
	wire _ArgumentNotifier_io_export_argIn_121_TREADY;
	wire _ArgumentNotifier_io_export_argIn_122_TREADY;
	wire _ArgumentNotifier_io_export_argIn_123_TREADY;
	wire _ArgumentNotifier_io_export_argIn_124_TREADY;
	wire _ArgumentNotifier_io_export_argIn_125_TREADY;
	wire _ArgumentNotifier_io_export_argIn_126_TREADY;
	wire _ArgumentNotifier_io_export_argIn_127_TREADY;
	wire _ArgumentNotifier_connStealNtw_0_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_0_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_0_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_1_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_1_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_1_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_2_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_2_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_2_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_3_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_3_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_3_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_4_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_4_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_4_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_5_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_5_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_5_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_6_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_6_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_6_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_7_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_7_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_7_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_8_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_8_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_8_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_9_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_9_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_9_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_10_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_10_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_10_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_11_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_11_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_11_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_12_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_12_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_12_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_13_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_13_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_13_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_14_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_14_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_14_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_15_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_15_data_qOutTask_valid;
	wire [255:0] _ArgumentNotifier_connStealNtw_15_data_qOutTask_bits;
	wire _Allocator_io_export_closureOut_0_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_0_TDATA;
	wire _Allocator_io_export_closureOut_1_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_1_TDATA;
	wire _Allocator_io_export_closureOut_2_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_2_TDATA;
	wire _Allocator_io_export_closureOut_3_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_3_TDATA;
	wire _Allocator_io_export_closureOut_4_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_4_TDATA;
	wire _Allocator_io_export_closureOut_5_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_5_TDATA;
	wire _Allocator_io_export_closureOut_6_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_6_TDATA;
	wire _Allocator_io_export_closureOut_7_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_7_TDATA;
	wire _Allocator_io_export_closureOut_8_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_8_TDATA;
	wire _Allocator_io_export_closureOut_9_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_9_TDATA;
	wire _Allocator_io_export_closureOut_10_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_10_TDATA;
	wire _Allocator_io_export_closureOut_11_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_11_TDATA;
	wire _Allocator_io_export_closureOut_12_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_12_TDATA;
	wire _Allocator_io_export_closureOut_13_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_13_TDATA;
	wire _Allocator_io_export_closureOut_14_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_14_TDATA;
	wire _Allocator_io_export_closureOut_15_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_15_TDATA;
	wire _Allocator_io_export_closureOut_16_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_16_TDATA;
	wire _Allocator_io_export_closureOut_17_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_17_TDATA;
	wire _Allocator_io_export_closureOut_18_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_18_TDATA;
	wire _Allocator_io_export_closureOut_19_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_19_TDATA;
	wire _Allocator_io_export_closureOut_20_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_20_TDATA;
	wire _Allocator_io_export_closureOut_21_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_21_TDATA;
	wire _Allocator_io_export_closureOut_22_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_22_TDATA;
	wire _Allocator_io_export_closureOut_23_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_23_TDATA;
	wire _Allocator_io_export_closureOut_24_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_24_TDATA;
	wire _Allocator_io_export_closureOut_25_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_25_TDATA;
	wire _Allocator_io_export_closureOut_26_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_26_TDATA;
	wire _Allocator_io_export_closureOut_27_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_27_TDATA;
	wire _Allocator_io_export_closureOut_28_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_28_TDATA;
	wire _Allocator_io_export_closureOut_29_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_29_TDATA;
	wire _Allocator_io_export_closureOut_30_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_30_TDATA;
	wire _Allocator_io_export_closureOut_31_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_31_TDATA;
	wire _Allocator_io_export_closureOut_32_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_32_TDATA;
	wire _Allocator_io_export_closureOut_33_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_33_TDATA;
	wire _Allocator_io_export_closureOut_34_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_34_TDATA;
	wire _Allocator_io_export_closureOut_35_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_35_TDATA;
	wire _Allocator_io_export_closureOut_36_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_36_TDATA;
	wire _Allocator_io_export_closureOut_37_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_37_TDATA;
	wire _Allocator_io_export_closureOut_38_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_38_TDATA;
	wire _Allocator_io_export_closureOut_39_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_39_TDATA;
	wire _Allocator_io_export_closureOut_40_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_40_TDATA;
	wire _Allocator_io_export_closureOut_41_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_41_TDATA;
	wire _Allocator_io_export_closureOut_42_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_42_TDATA;
	wire _Allocator_io_export_closureOut_43_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_43_TDATA;
	wire _Allocator_io_export_closureOut_44_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_44_TDATA;
	wire _Allocator_io_export_closureOut_45_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_45_TDATA;
	wire _Allocator_io_export_closureOut_46_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_46_TDATA;
	wire _Allocator_io_export_closureOut_47_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_47_TDATA;
	wire _Allocator_io_export_closureOut_48_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_48_TDATA;
	wire _Allocator_io_export_closureOut_49_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_49_TDATA;
	wire _Allocator_io_export_closureOut_50_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_50_TDATA;
	wire _Allocator_io_export_closureOut_51_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_51_TDATA;
	wire _Allocator_io_export_closureOut_52_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_52_TDATA;
	wire _Allocator_io_export_closureOut_53_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_53_TDATA;
	wire _Allocator_io_export_closureOut_54_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_54_TDATA;
	wire _Allocator_io_export_closureOut_55_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_55_TDATA;
	wire _Allocator_io_export_closureOut_56_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_56_TDATA;
	wire _Allocator_io_export_closureOut_57_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_57_TDATA;
	wire _Allocator_io_export_closureOut_58_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_58_TDATA;
	wire _Allocator_io_export_closureOut_59_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_59_TDATA;
	wire _Allocator_io_export_closureOut_60_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_60_TDATA;
	wire _Allocator_io_export_closureOut_61_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_61_TDATA;
	wire _Allocator_io_export_closureOut_62_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_62_TDATA;
	wire _Allocator_io_export_closureOut_63_TVALID;
	wire [63:0] _Allocator_io_export_closureOut_63_TDATA;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_0_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_0_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_0_b_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_1_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_1_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_1_b_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_2_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_2_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_2_b_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_3_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_3_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_3_b_bits_resp;
	wire _Scheduler_1_io_export_taskOut_0_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_0_TDATA;
	wire _Scheduler_1_io_export_taskOut_1_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_1_TDATA;
	wire _Scheduler_1_io_export_taskOut_2_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_2_TDATA;
	wire _Scheduler_1_io_export_taskOut_3_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_3_TDATA;
	wire _Scheduler_1_io_export_taskOut_4_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_4_TDATA;
	wire _Scheduler_1_io_export_taskOut_5_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_5_TDATA;
	wire _Scheduler_1_io_export_taskOut_6_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_6_TDATA;
	wire _Scheduler_1_io_export_taskOut_7_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_7_TDATA;
	wire _Scheduler_1_io_export_taskOut_8_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_8_TDATA;
	wire _Scheduler_1_io_export_taskOut_9_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_9_TDATA;
	wire _Scheduler_1_io_export_taskOut_10_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_10_TDATA;
	wire _Scheduler_1_io_export_taskOut_11_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_11_TDATA;
	wire _Scheduler_1_io_export_taskOut_12_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_12_TDATA;
	wire _Scheduler_1_io_export_taskOut_13_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_13_TDATA;
	wire _Scheduler_1_io_export_taskOut_14_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_14_TDATA;
	wire _Scheduler_1_io_export_taskOut_15_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_15_TDATA;
	wire _Scheduler_1_io_export_taskOut_16_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_16_TDATA;
	wire _Scheduler_1_io_export_taskOut_17_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_17_TDATA;
	wire _Scheduler_1_io_export_taskOut_18_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_18_TDATA;
	wire _Scheduler_1_io_export_taskOut_19_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_19_TDATA;
	wire _Scheduler_1_io_export_taskOut_20_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_20_TDATA;
	wire _Scheduler_1_io_export_taskOut_21_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_21_TDATA;
	wire _Scheduler_1_io_export_taskOut_22_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_22_TDATA;
	wire _Scheduler_1_io_export_taskOut_23_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_23_TDATA;
	wire _Scheduler_1_io_export_taskOut_24_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_24_TDATA;
	wire _Scheduler_1_io_export_taskOut_25_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_25_TDATA;
	wire _Scheduler_1_io_export_taskOut_26_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_26_TDATA;
	wire _Scheduler_1_io_export_taskOut_27_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_27_TDATA;
	wire _Scheduler_1_io_export_taskOut_28_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_28_TDATA;
	wire _Scheduler_1_io_export_taskOut_29_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_29_TDATA;
	wire _Scheduler_1_io_export_taskOut_30_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_30_TDATA;
	wire _Scheduler_1_io_export_taskOut_31_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_31_TDATA;
	wire _Scheduler_1_io_export_taskOut_32_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_32_TDATA;
	wire _Scheduler_1_io_export_taskOut_33_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_33_TDATA;
	wire _Scheduler_1_io_export_taskOut_34_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_34_TDATA;
	wire _Scheduler_1_io_export_taskOut_35_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_35_TDATA;
	wire _Scheduler_1_io_export_taskOut_36_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_36_TDATA;
	wire _Scheduler_1_io_export_taskOut_37_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_37_TDATA;
	wire _Scheduler_1_io_export_taskOut_38_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_38_TDATA;
	wire _Scheduler_1_io_export_taskOut_39_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_39_TDATA;
	wire _Scheduler_1_io_export_taskOut_40_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_40_TDATA;
	wire _Scheduler_1_io_export_taskOut_41_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_41_TDATA;
	wire _Scheduler_1_io_export_taskOut_42_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_42_TDATA;
	wire _Scheduler_1_io_export_taskOut_43_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_43_TDATA;
	wire _Scheduler_1_io_export_taskOut_44_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_44_TDATA;
	wire _Scheduler_1_io_export_taskOut_45_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_45_TDATA;
	wire _Scheduler_1_io_export_taskOut_46_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_46_TDATA;
	wire _Scheduler_1_io_export_taskOut_47_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_47_TDATA;
	wire _Scheduler_1_io_export_taskOut_48_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_48_TDATA;
	wire _Scheduler_1_io_export_taskOut_49_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_49_TDATA;
	wire _Scheduler_1_io_export_taskOut_50_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_50_TDATA;
	wire _Scheduler_1_io_export_taskOut_51_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_51_TDATA;
	wire _Scheduler_1_io_export_taskOut_52_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_52_TDATA;
	wire _Scheduler_1_io_export_taskOut_53_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_53_TDATA;
	wire _Scheduler_1_io_export_taskOut_54_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_54_TDATA;
	wire _Scheduler_1_io_export_taskOut_55_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_55_TDATA;
	wire _Scheduler_1_io_export_taskOut_56_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_56_TDATA;
	wire _Scheduler_1_io_export_taskOut_57_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_57_TDATA;
	wire _Scheduler_1_io_export_taskOut_58_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_58_TDATA;
	wire _Scheduler_1_io_export_taskOut_59_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_59_TDATA;
	wire _Scheduler_1_io_export_taskOut_60_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_60_TDATA;
	wire _Scheduler_1_io_export_taskOut_61_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_61_TDATA;
	wire _Scheduler_1_io_export_taskOut_62_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_62_TDATA;
	wire _Scheduler_1_io_export_taskOut_63_TVALID;
	wire [255:0] _Scheduler_1_io_export_taskOut_63_TDATA;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_ar_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_r_valid;
	wire [63:0] _Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_data;
	wire [1:0] _Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_resp;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_aw_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_w_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_b_valid;
	wire [1:0] _Scheduler_1_io_internal_axi_mgmt_vss_0_b_bits_resp;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_1_ar_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_1_r_valid;
	wire [63:0] _Scheduler_1_io_internal_axi_mgmt_vss_1_r_bits_data;
	wire [1:0] _Scheduler_1_io_internal_axi_mgmt_vss_1_r_bits_resp;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_1_aw_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_1_w_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_1_b_valid;
	wire [1:0] _Scheduler_1_io_internal_axi_mgmt_vss_1_b_bits_resp;
	wire _Scheduler_1_connArgumentNotifier_0_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_0_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_1_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_1_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_2_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_2_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_3_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_3_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_4_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_4_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_5_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_5_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_6_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_6_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_7_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_7_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_8_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_8_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_9_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_9_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_10_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_10_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_11_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_11_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_12_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_12_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_13_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_13_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_14_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_14_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_15_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_15_data_qOutTask_ready;
	wire _peArray_63_1_argOut_TVALID;
	wire [63:0] _peArray_63_1_argOut_TDATA;
	wire _peArray_63_1_taskIn_TREADY;
	wire _peArray_62_1_argOut_TVALID;
	wire [63:0] _peArray_62_1_argOut_TDATA;
	wire _peArray_62_1_taskIn_TREADY;
	wire _peArray_61_1_argOut_TVALID;
	wire [63:0] _peArray_61_1_argOut_TDATA;
	wire _peArray_61_1_taskIn_TREADY;
	wire _peArray_60_1_argOut_TVALID;
	wire [63:0] _peArray_60_1_argOut_TDATA;
	wire _peArray_60_1_taskIn_TREADY;
	wire _peArray_59_1_argOut_TVALID;
	wire [63:0] _peArray_59_1_argOut_TDATA;
	wire _peArray_59_1_taskIn_TREADY;
	wire _peArray_58_1_argOut_TVALID;
	wire [63:0] _peArray_58_1_argOut_TDATA;
	wire _peArray_58_1_taskIn_TREADY;
	wire _peArray_57_1_argOut_TVALID;
	wire [63:0] _peArray_57_1_argOut_TDATA;
	wire _peArray_57_1_taskIn_TREADY;
	wire _peArray_56_1_argOut_TVALID;
	wire [63:0] _peArray_56_1_argOut_TDATA;
	wire _peArray_56_1_taskIn_TREADY;
	wire _peArray_55_1_argOut_TVALID;
	wire [63:0] _peArray_55_1_argOut_TDATA;
	wire _peArray_55_1_taskIn_TREADY;
	wire _peArray_54_1_argOut_TVALID;
	wire [63:0] _peArray_54_1_argOut_TDATA;
	wire _peArray_54_1_taskIn_TREADY;
	wire _peArray_53_1_argOut_TVALID;
	wire [63:0] _peArray_53_1_argOut_TDATA;
	wire _peArray_53_1_taskIn_TREADY;
	wire _peArray_52_1_argOut_TVALID;
	wire [63:0] _peArray_52_1_argOut_TDATA;
	wire _peArray_52_1_taskIn_TREADY;
	wire _peArray_51_1_argOut_TVALID;
	wire [63:0] _peArray_51_1_argOut_TDATA;
	wire _peArray_51_1_taskIn_TREADY;
	wire _peArray_50_1_argOut_TVALID;
	wire [63:0] _peArray_50_1_argOut_TDATA;
	wire _peArray_50_1_taskIn_TREADY;
	wire _peArray_49_1_argOut_TVALID;
	wire [63:0] _peArray_49_1_argOut_TDATA;
	wire _peArray_49_1_taskIn_TREADY;
	wire _peArray_48_1_argOut_TVALID;
	wire [63:0] _peArray_48_1_argOut_TDATA;
	wire _peArray_48_1_taskIn_TREADY;
	wire _peArray_47_1_argOut_TVALID;
	wire [63:0] _peArray_47_1_argOut_TDATA;
	wire _peArray_47_1_taskIn_TREADY;
	wire _peArray_46_1_argOut_TVALID;
	wire [63:0] _peArray_46_1_argOut_TDATA;
	wire _peArray_46_1_taskIn_TREADY;
	wire _peArray_45_1_argOut_TVALID;
	wire [63:0] _peArray_45_1_argOut_TDATA;
	wire _peArray_45_1_taskIn_TREADY;
	wire _peArray_44_1_argOut_TVALID;
	wire [63:0] _peArray_44_1_argOut_TDATA;
	wire _peArray_44_1_taskIn_TREADY;
	wire _peArray_43_1_argOut_TVALID;
	wire [63:0] _peArray_43_1_argOut_TDATA;
	wire _peArray_43_1_taskIn_TREADY;
	wire _peArray_42_1_argOut_TVALID;
	wire [63:0] _peArray_42_1_argOut_TDATA;
	wire _peArray_42_1_taskIn_TREADY;
	wire _peArray_41_1_argOut_TVALID;
	wire [63:0] _peArray_41_1_argOut_TDATA;
	wire _peArray_41_1_taskIn_TREADY;
	wire _peArray_40_1_argOut_TVALID;
	wire [63:0] _peArray_40_1_argOut_TDATA;
	wire _peArray_40_1_taskIn_TREADY;
	wire _peArray_39_1_argOut_TVALID;
	wire [63:0] _peArray_39_1_argOut_TDATA;
	wire _peArray_39_1_taskIn_TREADY;
	wire _peArray_38_1_argOut_TVALID;
	wire [63:0] _peArray_38_1_argOut_TDATA;
	wire _peArray_38_1_taskIn_TREADY;
	wire _peArray_37_1_argOut_TVALID;
	wire [63:0] _peArray_37_1_argOut_TDATA;
	wire _peArray_37_1_taskIn_TREADY;
	wire _peArray_36_1_argOut_TVALID;
	wire [63:0] _peArray_36_1_argOut_TDATA;
	wire _peArray_36_1_taskIn_TREADY;
	wire _peArray_35_1_argOut_TVALID;
	wire [63:0] _peArray_35_1_argOut_TDATA;
	wire _peArray_35_1_taskIn_TREADY;
	wire _peArray_34_1_argOut_TVALID;
	wire [63:0] _peArray_34_1_argOut_TDATA;
	wire _peArray_34_1_taskIn_TREADY;
	wire _peArray_33_1_argOut_TVALID;
	wire [63:0] _peArray_33_1_argOut_TDATA;
	wire _peArray_33_1_taskIn_TREADY;
	wire _peArray_32_1_argOut_TVALID;
	wire [63:0] _peArray_32_1_argOut_TDATA;
	wire _peArray_32_1_taskIn_TREADY;
	wire _peArray_31_1_argOut_TVALID;
	wire [63:0] _peArray_31_1_argOut_TDATA;
	wire _peArray_31_1_taskIn_TREADY;
	wire _peArray_30_1_argOut_TVALID;
	wire [63:0] _peArray_30_1_argOut_TDATA;
	wire _peArray_30_1_taskIn_TREADY;
	wire _peArray_29_1_argOut_TVALID;
	wire [63:0] _peArray_29_1_argOut_TDATA;
	wire _peArray_29_1_taskIn_TREADY;
	wire _peArray_28_1_argOut_TVALID;
	wire [63:0] _peArray_28_1_argOut_TDATA;
	wire _peArray_28_1_taskIn_TREADY;
	wire _peArray_27_1_argOut_TVALID;
	wire [63:0] _peArray_27_1_argOut_TDATA;
	wire _peArray_27_1_taskIn_TREADY;
	wire _peArray_26_1_argOut_TVALID;
	wire [63:0] _peArray_26_1_argOut_TDATA;
	wire _peArray_26_1_taskIn_TREADY;
	wire _peArray_25_1_argOut_TVALID;
	wire [63:0] _peArray_25_1_argOut_TDATA;
	wire _peArray_25_1_taskIn_TREADY;
	wire _peArray_24_1_argOut_TVALID;
	wire [63:0] _peArray_24_1_argOut_TDATA;
	wire _peArray_24_1_taskIn_TREADY;
	wire _peArray_23_1_argOut_TVALID;
	wire [63:0] _peArray_23_1_argOut_TDATA;
	wire _peArray_23_1_taskIn_TREADY;
	wire _peArray_22_1_argOut_TVALID;
	wire [63:0] _peArray_22_1_argOut_TDATA;
	wire _peArray_22_1_taskIn_TREADY;
	wire _peArray_21_1_argOut_TVALID;
	wire [63:0] _peArray_21_1_argOut_TDATA;
	wire _peArray_21_1_taskIn_TREADY;
	wire _peArray_20_1_argOut_TVALID;
	wire [63:0] _peArray_20_1_argOut_TDATA;
	wire _peArray_20_1_taskIn_TREADY;
	wire _peArray_19_1_argOut_TVALID;
	wire [63:0] _peArray_19_1_argOut_TDATA;
	wire _peArray_19_1_taskIn_TREADY;
	wire _peArray_18_1_argOut_TVALID;
	wire [63:0] _peArray_18_1_argOut_TDATA;
	wire _peArray_18_1_taskIn_TREADY;
	wire _peArray_17_1_argOut_TVALID;
	wire [63:0] _peArray_17_1_argOut_TDATA;
	wire _peArray_17_1_taskIn_TREADY;
	wire _peArray_16_1_argOut_TVALID;
	wire [63:0] _peArray_16_1_argOut_TDATA;
	wire _peArray_16_1_taskIn_TREADY;
	wire _peArray_15_1_argOut_TVALID;
	wire [63:0] _peArray_15_1_argOut_TDATA;
	wire _peArray_15_1_taskIn_TREADY;
	wire _peArray_14_1_argOut_TVALID;
	wire [63:0] _peArray_14_1_argOut_TDATA;
	wire _peArray_14_1_taskIn_TREADY;
	wire _peArray_13_1_argOut_TVALID;
	wire [63:0] _peArray_13_1_argOut_TDATA;
	wire _peArray_13_1_taskIn_TREADY;
	wire _peArray_12_1_argOut_TVALID;
	wire [63:0] _peArray_12_1_argOut_TDATA;
	wire _peArray_12_1_taskIn_TREADY;
	wire _peArray_11_1_argOut_TVALID;
	wire [63:0] _peArray_11_1_argOut_TDATA;
	wire _peArray_11_1_taskIn_TREADY;
	wire _peArray_10_1_argOut_TVALID;
	wire [63:0] _peArray_10_1_argOut_TDATA;
	wire _peArray_10_1_taskIn_TREADY;
	wire _peArray_9_1_argOut_TVALID;
	wire [63:0] _peArray_9_1_argOut_TDATA;
	wire _peArray_9_1_taskIn_TREADY;
	wire _peArray_8_1_argOut_TVALID;
	wire [63:0] _peArray_8_1_argOut_TDATA;
	wire _peArray_8_1_taskIn_TREADY;
	wire _peArray_7_1_argOut_TVALID;
	wire [63:0] _peArray_7_1_argOut_TDATA;
	wire _peArray_7_1_taskIn_TREADY;
	wire _peArray_6_1_argOut_TVALID;
	wire [63:0] _peArray_6_1_argOut_TDATA;
	wire _peArray_6_1_taskIn_TREADY;
	wire _peArray_5_1_argOut_TVALID;
	wire [63:0] _peArray_5_1_argOut_TDATA;
	wire _peArray_5_1_taskIn_TREADY;
	wire _peArray_4_1_argOut_TVALID;
	wire [63:0] _peArray_4_1_argOut_TDATA;
	wire _peArray_4_1_taskIn_TREADY;
	wire _peArray_3_1_argOut_TVALID;
	wire [63:0] _peArray_3_1_argOut_TDATA;
	wire _peArray_3_1_taskIn_TREADY;
	wire _peArray_2_1_argOut_TVALID;
	wire [63:0] _peArray_2_1_argOut_TDATA;
	wire _peArray_2_1_taskIn_TREADY;
	wire _peArray_1_1_argOut_TVALID;
	wire [63:0] _peArray_1_1_argOut_TDATA;
	wire _peArray_1_1_taskIn_TREADY;
	wire _peArray_0_1_argOut_TVALID;
	wire [63:0] _peArray_0_1_argOut_TDATA;
	wire _peArray_0_1_taskIn_TREADY;
	wire _Scheduler_io_export_taskOut_0_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_0_TDATA;
	wire _Scheduler_io_export_taskOut_1_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_1_TDATA;
	wire _Scheduler_io_export_taskOut_2_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_2_TDATA;
	wire _Scheduler_io_export_taskOut_3_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_3_TDATA;
	wire _Scheduler_io_export_taskOut_4_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_4_TDATA;
	wire _Scheduler_io_export_taskOut_5_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_5_TDATA;
	wire _Scheduler_io_export_taskOut_6_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_6_TDATA;
	wire _Scheduler_io_export_taskOut_7_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_7_TDATA;
	wire _Scheduler_io_export_taskOut_8_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_8_TDATA;
	wire _Scheduler_io_export_taskOut_9_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_9_TDATA;
	wire _Scheduler_io_export_taskOut_10_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_10_TDATA;
	wire _Scheduler_io_export_taskOut_11_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_11_TDATA;
	wire _Scheduler_io_export_taskOut_12_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_12_TDATA;
	wire _Scheduler_io_export_taskOut_13_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_13_TDATA;
	wire _Scheduler_io_export_taskOut_14_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_14_TDATA;
	wire _Scheduler_io_export_taskOut_15_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_15_TDATA;
	wire _Scheduler_io_export_taskOut_16_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_16_TDATA;
	wire _Scheduler_io_export_taskOut_17_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_17_TDATA;
	wire _Scheduler_io_export_taskOut_18_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_18_TDATA;
	wire _Scheduler_io_export_taskOut_19_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_19_TDATA;
	wire _Scheduler_io_export_taskOut_20_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_20_TDATA;
	wire _Scheduler_io_export_taskOut_21_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_21_TDATA;
	wire _Scheduler_io_export_taskOut_22_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_22_TDATA;
	wire _Scheduler_io_export_taskOut_23_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_23_TDATA;
	wire _Scheduler_io_export_taskOut_24_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_24_TDATA;
	wire _Scheduler_io_export_taskOut_25_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_25_TDATA;
	wire _Scheduler_io_export_taskOut_26_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_26_TDATA;
	wire _Scheduler_io_export_taskOut_27_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_27_TDATA;
	wire _Scheduler_io_export_taskOut_28_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_28_TDATA;
	wire _Scheduler_io_export_taskOut_29_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_29_TDATA;
	wire _Scheduler_io_export_taskOut_30_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_30_TDATA;
	wire _Scheduler_io_export_taskOut_31_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_31_TDATA;
	wire _Scheduler_io_export_taskOut_32_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_32_TDATA;
	wire _Scheduler_io_export_taskOut_33_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_33_TDATA;
	wire _Scheduler_io_export_taskOut_34_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_34_TDATA;
	wire _Scheduler_io_export_taskOut_35_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_35_TDATA;
	wire _Scheduler_io_export_taskOut_36_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_36_TDATA;
	wire _Scheduler_io_export_taskOut_37_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_37_TDATA;
	wire _Scheduler_io_export_taskOut_38_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_38_TDATA;
	wire _Scheduler_io_export_taskOut_39_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_39_TDATA;
	wire _Scheduler_io_export_taskOut_40_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_40_TDATA;
	wire _Scheduler_io_export_taskOut_41_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_41_TDATA;
	wire _Scheduler_io_export_taskOut_42_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_42_TDATA;
	wire _Scheduler_io_export_taskOut_43_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_43_TDATA;
	wire _Scheduler_io_export_taskOut_44_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_44_TDATA;
	wire _Scheduler_io_export_taskOut_45_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_45_TDATA;
	wire _Scheduler_io_export_taskOut_46_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_46_TDATA;
	wire _Scheduler_io_export_taskOut_47_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_47_TDATA;
	wire _Scheduler_io_export_taskOut_48_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_48_TDATA;
	wire _Scheduler_io_export_taskOut_49_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_49_TDATA;
	wire _Scheduler_io_export_taskOut_50_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_50_TDATA;
	wire _Scheduler_io_export_taskOut_51_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_51_TDATA;
	wire _Scheduler_io_export_taskOut_52_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_52_TDATA;
	wire _Scheduler_io_export_taskOut_53_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_53_TDATA;
	wire _Scheduler_io_export_taskOut_54_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_54_TDATA;
	wire _Scheduler_io_export_taskOut_55_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_55_TDATA;
	wire _Scheduler_io_export_taskOut_56_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_56_TDATA;
	wire _Scheduler_io_export_taskOut_57_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_57_TDATA;
	wire _Scheduler_io_export_taskOut_58_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_58_TDATA;
	wire _Scheduler_io_export_taskOut_59_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_59_TDATA;
	wire _Scheduler_io_export_taskOut_60_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_60_TDATA;
	wire _Scheduler_io_export_taskOut_61_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_61_TDATA;
	wire _Scheduler_io_export_taskOut_62_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_62_TDATA;
	wire _Scheduler_io_export_taskOut_63_TVALID;
	wire [127:0] _Scheduler_io_export_taskOut_63_TDATA;
	wire _Scheduler_io_export_taskIn_0_TREADY;
	wire _Scheduler_io_export_taskIn_1_TREADY;
	wire _Scheduler_io_export_taskIn_2_TREADY;
	wire _Scheduler_io_export_taskIn_3_TREADY;
	wire _Scheduler_io_export_taskIn_4_TREADY;
	wire _Scheduler_io_export_taskIn_5_TREADY;
	wire _Scheduler_io_export_taskIn_6_TREADY;
	wire _Scheduler_io_export_taskIn_7_TREADY;
	wire _Scheduler_io_export_taskIn_8_TREADY;
	wire _Scheduler_io_export_taskIn_9_TREADY;
	wire _Scheduler_io_export_taskIn_10_TREADY;
	wire _Scheduler_io_export_taskIn_11_TREADY;
	wire _Scheduler_io_export_taskIn_12_TREADY;
	wire _Scheduler_io_export_taskIn_13_TREADY;
	wire _Scheduler_io_export_taskIn_14_TREADY;
	wire _Scheduler_io_export_taskIn_15_TREADY;
	wire _Scheduler_io_export_taskIn_16_TREADY;
	wire _Scheduler_io_export_taskIn_17_TREADY;
	wire _Scheduler_io_export_taskIn_18_TREADY;
	wire _Scheduler_io_export_taskIn_19_TREADY;
	wire _Scheduler_io_export_taskIn_20_TREADY;
	wire _Scheduler_io_export_taskIn_21_TREADY;
	wire _Scheduler_io_export_taskIn_22_TREADY;
	wire _Scheduler_io_export_taskIn_23_TREADY;
	wire _Scheduler_io_export_taskIn_24_TREADY;
	wire _Scheduler_io_export_taskIn_25_TREADY;
	wire _Scheduler_io_export_taskIn_26_TREADY;
	wire _Scheduler_io_export_taskIn_27_TREADY;
	wire _Scheduler_io_export_taskIn_28_TREADY;
	wire _Scheduler_io_export_taskIn_29_TREADY;
	wire _Scheduler_io_export_taskIn_30_TREADY;
	wire _Scheduler_io_export_taskIn_31_TREADY;
	wire _Scheduler_io_export_taskIn_32_TREADY;
	wire _Scheduler_io_export_taskIn_33_TREADY;
	wire _Scheduler_io_export_taskIn_34_TREADY;
	wire _Scheduler_io_export_taskIn_35_TREADY;
	wire _Scheduler_io_export_taskIn_36_TREADY;
	wire _Scheduler_io_export_taskIn_37_TREADY;
	wire _Scheduler_io_export_taskIn_38_TREADY;
	wire _Scheduler_io_export_taskIn_39_TREADY;
	wire _Scheduler_io_export_taskIn_40_TREADY;
	wire _Scheduler_io_export_taskIn_41_TREADY;
	wire _Scheduler_io_export_taskIn_42_TREADY;
	wire _Scheduler_io_export_taskIn_43_TREADY;
	wire _Scheduler_io_export_taskIn_44_TREADY;
	wire _Scheduler_io_export_taskIn_45_TREADY;
	wire _Scheduler_io_export_taskIn_46_TREADY;
	wire _Scheduler_io_export_taskIn_47_TREADY;
	wire _Scheduler_io_export_taskIn_48_TREADY;
	wire _Scheduler_io_export_taskIn_49_TREADY;
	wire _Scheduler_io_export_taskIn_50_TREADY;
	wire _Scheduler_io_export_taskIn_51_TREADY;
	wire _Scheduler_io_export_taskIn_52_TREADY;
	wire _Scheduler_io_export_taskIn_53_TREADY;
	wire _Scheduler_io_export_taskIn_54_TREADY;
	wire _Scheduler_io_export_taskIn_55_TREADY;
	wire _Scheduler_io_export_taskIn_56_TREADY;
	wire _Scheduler_io_export_taskIn_57_TREADY;
	wire _Scheduler_io_export_taskIn_58_TREADY;
	wire _Scheduler_io_export_taskIn_59_TREADY;
	wire _Scheduler_io_export_taskIn_60_TREADY;
	wire _Scheduler_io_export_taskIn_61_TREADY;
	wire _Scheduler_io_export_taskIn_62_TREADY;
	wire _Scheduler_io_export_taskIn_63_TREADY;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_ar_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_r_valid;
	wire [63:0] _Scheduler_io_internal_axi_mgmt_vss_0_r_bits_data;
	wire [1:0] _Scheduler_io_internal_axi_mgmt_vss_0_r_bits_resp;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_aw_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_w_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_b_valid;
	wire [1:0] _Scheduler_io_internal_axi_mgmt_vss_0_b_bits_resp;
	wire _Scheduler_io_internal_axi_mgmt_vss_1_ar_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_1_r_valid;
	wire [63:0] _Scheduler_io_internal_axi_mgmt_vss_1_r_bits_data;
	wire [1:0] _Scheduler_io_internal_axi_mgmt_vss_1_r_bits_resp;
	wire _Scheduler_io_internal_axi_mgmt_vss_1_aw_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_1_w_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_1_b_valid;
	wire [1:0] _Scheduler_io_internal_axi_mgmt_vss_1_b_bits_resp;
	wire _peArray_63_closureIn_TREADY;
	wire _peArray_63_argOut_TVALID;
	wire [63:0] _peArray_63_argOut_TDATA;
	wire _peArray_63_taskOut_TVALID;
	wire [127:0] _peArray_63_taskOut_TDATA;
	wire _peArray_63_taskIn_TREADY;
	wire _peArray_62_closureIn_TREADY;
	wire _peArray_62_argOut_TVALID;
	wire [63:0] _peArray_62_argOut_TDATA;
	wire _peArray_62_taskOut_TVALID;
	wire [127:0] _peArray_62_taskOut_TDATA;
	wire _peArray_62_taskIn_TREADY;
	wire _peArray_61_closureIn_TREADY;
	wire _peArray_61_argOut_TVALID;
	wire [63:0] _peArray_61_argOut_TDATA;
	wire _peArray_61_taskOut_TVALID;
	wire [127:0] _peArray_61_taskOut_TDATA;
	wire _peArray_61_taskIn_TREADY;
	wire _peArray_60_closureIn_TREADY;
	wire _peArray_60_argOut_TVALID;
	wire [63:0] _peArray_60_argOut_TDATA;
	wire _peArray_60_taskOut_TVALID;
	wire [127:0] _peArray_60_taskOut_TDATA;
	wire _peArray_60_taskIn_TREADY;
	wire _peArray_59_closureIn_TREADY;
	wire _peArray_59_argOut_TVALID;
	wire [63:0] _peArray_59_argOut_TDATA;
	wire _peArray_59_taskOut_TVALID;
	wire [127:0] _peArray_59_taskOut_TDATA;
	wire _peArray_59_taskIn_TREADY;
	wire _peArray_58_closureIn_TREADY;
	wire _peArray_58_argOut_TVALID;
	wire [63:0] _peArray_58_argOut_TDATA;
	wire _peArray_58_taskOut_TVALID;
	wire [127:0] _peArray_58_taskOut_TDATA;
	wire _peArray_58_taskIn_TREADY;
	wire _peArray_57_closureIn_TREADY;
	wire _peArray_57_argOut_TVALID;
	wire [63:0] _peArray_57_argOut_TDATA;
	wire _peArray_57_taskOut_TVALID;
	wire [127:0] _peArray_57_taskOut_TDATA;
	wire _peArray_57_taskIn_TREADY;
	wire _peArray_56_closureIn_TREADY;
	wire _peArray_56_argOut_TVALID;
	wire [63:0] _peArray_56_argOut_TDATA;
	wire _peArray_56_taskOut_TVALID;
	wire [127:0] _peArray_56_taskOut_TDATA;
	wire _peArray_56_taskIn_TREADY;
	wire _peArray_55_closureIn_TREADY;
	wire _peArray_55_argOut_TVALID;
	wire [63:0] _peArray_55_argOut_TDATA;
	wire _peArray_55_taskOut_TVALID;
	wire [127:0] _peArray_55_taskOut_TDATA;
	wire _peArray_55_taskIn_TREADY;
	wire _peArray_54_closureIn_TREADY;
	wire _peArray_54_argOut_TVALID;
	wire [63:0] _peArray_54_argOut_TDATA;
	wire _peArray_54_taskOut_TVALID;
	wire [127:0] _peArray_54_taskOut_TDATA;
	wire _peArray_54_taskIn_TREADY;
	wire _peArray_53_closureIn_TREADY;
	wire _peArray_53_argOut_TVALID;
	wire [63:0] _peArray_53_argOut_TDATA;
	wire _peArray_53_taskOut_TVALID;
	wire [127:0] _peArray_53_taskOut_TDATA;
	wire _peArray_53_taskIn_TREADY;
	wire _peArray_52_closureIn_TREADY;
	wire _peArray_52_argOut_TVALID;
	wire [63:0] _peArray_52_argOut_TDATA;
	wire _peArray_52_taskOut_TVALID;
	wire [127:0] _peArray_52_taskOut_TDATA;
	wire _peArray_52_taskIn_TREADY;
	wire _peArray_51_closureIn_TREADY;
	wire _peArray_51_argOut_TVALID;
	wire [63:0] _peArray_51_argOut_TDATA;
	wire _peArray_51_taskOut_TVALID;
	wire [127:0] _peArray_51_taskOut_TDATA;
	wire _peArray_51_taskIn_TREADY;
	wire _peArray_50_closureIn_TREADY;
	wire _peArray_50_argOut_TVALID;
	wire [63:0] _peArray_50_argOut_TDATA;
	wire _peArray_50_taskOut_TVALID;
	wire [127:0] _peArray_50_taskOut_TDATA;
	wire _peArray_50_taskIn_TREADY;
	wire _peArray_49_closureIn_TREADY;
	wire _peArray_49_argOut_TVALID;
	wire [63:0] _peArray_49_argOut_TDATA;
	wire _peArray_49_taskOut_TVALID;
	wire [127:0] _peArray_49_taskOut_TDATA;
	wire _peArray_49_taskIn_TREADY;
	wire _peArray_48_closureIn_TREADY;
	wire _peArray_48_argOut_TVALID;
	wire [63:0] _peArray_48_argOut_TDATA;
	wire _peArray_48_taskOut_TVALID;
	wire [127:0] _peArray_48_taskOut_TDATA;
	wire _peArray_48_taskIn_TREADY;
	wire _peArray_47_closureIn_TREADY;
	wire _peArray_47_argOut_TVALID;
	wire [63:0] _peArray_47_argOut_TDATA;
	wire _peArray_47_taskOut_TVALID;
	wire [127:0] _peArray_47_taskOut_TDATA;
	wire _peArray_47_taskIn_TREADY;
	wire _peArray_46_closureIn_TREADY;
	wire _peArray_46_argOut_TVALID;
	wire [63:0] _peArray_46_argOut_TDATA;
	wire _peArray_46_taskOut_TVALID;
	wire [127:0] _peArray_46_taskOut_TDATA;
	wire _peArray_46_taskIn_TREADY;
	wire _peArray_45_closureIn_TREADY;
	wire _peArray_45_argOut_TVALID;
	wire [63:0] _peArray_45_argOut_TDATA;
	wire _peArray_45_taskOut_TVALID;
	wire [127:0] _peArray_45_taskOut_TDATA;
	wire _peArray_45_taskIn_TREADY;
	wire _peArray_44_closureIn_TREADY;
	wire _peArray_44_argOut_TVALID;
	wire [63:0] _peArray_44_argOut_TDATA;
	wire _peArray_44_taskOut_TVALID;
	wire [127:0] _peArray_44_taskOut_TDATA;
	wire _peArray_44_taskIn_TREADY;
	wire _peArray_43_closureIn_TREADY;
	wire _peArray_43_argOut_TVALID;
	wire [63:0] _peArray_43_argOut_TDATA;
	wire _peArray_43_taskOut_TVALID;
	wire [127:0] _peArray_43_taskOut_TDATA;
	wire _peArray_43_taskIn_TREADY;
	wire _peArray_42_closureIn_TREADY;
	wire _peArray_42_argOut_TVALID;
	wire [63:0] _peArray_42_argOut_TDATA;
	wire _peArray_42_taskOut_TVALID;
	wire [127:0] _peArray_42_taskOut_TDATA;
	wire _peArray_42_taskIn_TREADY;
	wire _peArray_41_closureIn_TREADY;
	wire _peArray_41_argOut_TVALID;
	wire [63:0] _peArray_41_argOut_TDATA;
	wire _peArray_41_taskOut_TVALID;
	wire [127:0] _peArray_41_taskOut_TDATA;
	wire _peArray_41_taskIn_TREADY;
	wire _peArray_40_closureIn_TREADY;
	wire _peArray_40_argOut_TVALID;
	wire [63:0] _peArray_40_argOut_TDATA;
	wire _peArray_40_taskOut_TVALID;
	wire [127:0] _peArray_40_taskOut_TDATA;
	wire _peArray_40_taskIn_TREADY;
	wire _peArray_39_closureIn_TREADY;
	wire _peArray_39_argOut_TVALID;
	wire [63:0] _peArray_39_argOut_TDATA;
	wire _peArray_39_taskOut_TVALID;
	wire [127:0] _peArray_39_taskOut_TDATA;
	wire _peArray_39_taskIn_TREADY;
	wire _peArray_38_closureIn_TREADY;
	wire _peArray_38_argOut_TVALID;
	wire [63:0] _peArray_38_argOut_TDATA;
	wire _peArray_38_taskOut_TVALID;
	wire [127:0] _peArray_38_taskOut_TDATA;
	wire _peArray_38_taskIn_TREADY;
	wire _peArray_37_closureIn_TREADY;
	wire _peArray_37_argOut_TVALID;
	wire [63:0] _peArray_37_argOut_TDATA;
	wire _peArray_37_taskOut_TVALID;
	wire [127:0] _peArray_37_taskOut_TDATA;
	wire _peArray_37_taskIn_TREADY;
	wire _peArray_36_closureIn_TREADY;
	wire _peArray_36_argOut_TVALID;
	wire [63:0] _peArray_36_argOut_TDATA;
	wire _peArray_36_taskOut_TVALID;
	wire [127:0] _peArray_36_taskOut_TDATA;
	wire _peArray_36_taskIn_TREADY;
	wire _peArray_35_closureIn_TREADY;
	wire _peArray_35_argOut_TVALID;
	wire [63:0] _peArray_35_argOut_TDATA;
	wire _peArray_35_taskOut_TVALID;
	wire [127:0] _peArray_35_taskOut_TDATA;
	wire _peArray_35_taskIn_TREADY;
	wire _peArray_34_closureIn_TREADY;
	wire _peArray_34_argOut_TVALID;
	wire [63:0] _peArray_34_argOut_TDATA;
	wire _peArray_34_taskOut_TVALID;
	wire [127:0] _peArray_34_taskOut_TDATA;
	wire _peArray_34_taskIn_TREADY;
	wire _peArray_33_closureIn_TREADY;
	wire _peArray_33_argOut_TVALID;
	wire [63:0] _peArray_33_argOut_TDATA;
	wire _peArray_33_taskOut_TVALID;
	wire [127:0] _peArray_33_taskOut_TDATA;
	wire _peArray_33_taskIn_TREADY;
	wire _peArray_32_closureIn_TREADY;
	wire _peArray_32_argOut_TVALID;
	wire [63:0] _peArray_32_argOut_TDATA;
	wire _peArray_32_taskOut_TVALID;
	wire [127:0] _peArray_32_taskOut_TDATA;
	wire _peArray_32_taskIn_TREADY;
	wire _peArray_31_closureIn_TREADY;
	wire _peArray_31_argOut_TVALID;
	wire [63:0] _peArray_31_argOut_TDATA;
	wire _peArray_31_taskOut_TVALID;
	wire [127:0] _peArray_31_taskOut_TDATA;
	wire _peArray_31_taskIn_TREADY;
	wire _peArray_30_closureIn_TREADY;
	wire _peArray_30_argOut_TVALID;
	wire [63:0] _peArray_30_argOut_TDATA;
	wire _peArray_30_taskOut_TVALID;
	wire [127:0] _peArray_30_taskOut_TDATA;
	wire _peArray_30_taskIn_TREADY;
	wire _peArray_29_closureIn_TREADY;
	wire _peArray_29_argOut_TVALID;
	wire [63:0] _peArray_29_argOut_TDATA;
	wire _peArray_29_taskOut_TVALID;
	wire [127:0] _peArray_29_taskOut_TDATA;
	wire _peArray_29_taskIn_TREADY;
	wire _peArray_28_closureIn_TREADY;
	wire _peArray_28_argOut_TVALID;
	wire [63:0] _peArray_28_argOut_TDATA;
	wire _peArray_28_taskOut_TVALID;
	wire [127:0] _peArray_28_taskOut_TDATA;
	wire _peArray_28_taskIn_TREADY;
	wire _peArray_27_closureIn_TREADY;
	wire _peArray_27_argOut_TVALID;
	wire [63:0] _peArray_27_argOut_TDATA;
	wire _peArray_27_taskOut_TVALID;
	wire [127:0] _peArray_27_taskOut_TDATA;
	wire _peArray_27_taskIn_TREADY;
	wire _peArray_26_closureIn_TREADY;
	wire _peArray_26_argOut_TVALID;
	wire [63:0] _peArray_26_argOut_TDATA;
	wire _peArray_26_taskOut_TVALID;
	wire [127:0] _peArray_26_taskOut_TDATA;
	wire _peArray_26_taskIn_TREADY;
	wire _peArray_25_closureIn_TREADY;
	wire _peArray_25_argOut_TVALID;
	wire [63:0] _peArray_25_argOut_TDATA;
	wire _peArray_25_taskOut_TVALID;
	wire [127:0] _peArray_25_taskOut_TDATA;
	wire _peArray_25_taskIn_TREADY;
	wire _peArray_24_closureIn_TREADY;
	wire _peArray_24_argOut_TVALID;
	wire [63:0] _peArray_24_argOut_TDATA;
	wire _peArray_24_taskOut_TVALID;
	wire [127:0] _peArray_24_taskOut_TDATA;
	wire _peArray_24_taskIn_TREADY;
	wire _peArray_23_closureIn_TREADY;
	wire _peArray_23_argOut_TVALID;
	wire [63:0] _peArray_23_argOut_TDATA;
	wire _peArray_23_taskOut_TVALID;
	wire [127:0] _peArray_23_taskOut_TDATA;
	wire _peArray_23_taskIn_TREADY;
	wire _peArray_22_closureIn_TREADY;
	wire _peArray_22_argOut_TVALID;
	wire [63:0] _peArray_22_argOut_TDATA;
	wire _peArray_22_taskOut_TVALID;
	wire [127:0] _peArray_22_taskOut_TDATA;
	wire _peArray_22_taskIn_TREADY;
	wire _peArray_21_closureIn_TREADY;
	wire _peArray_21_argOut_TVALID;
	wire [63:0] _peArray_21_argOut_TDATA;
	wire _peArray_21_taskOut_TVALID;
	wire [127:0] _peArray_21_taskOut_TDATA;
	wire _peArray_21_taskIn_TREADY;
	wire _peArray_20_closureIn_TREADY;
	wire _peArray_20_argOut_TVALID;
	wire [63:0] _peArray_20_argOut_TDATA;
	wire _peArray_20_taskOut_TVALID;
	wire [127:0] _peArray_20_taskOut_TDATA;
	wire _peArray_20_taskIn_TREADY;
	wire _peArray_19_closureIn_TREADY;
	wire _peArray_19_argOut_TVALID;
	wire [63:0] _peArray_19_argOut_TDATA;
	wire _peArray_19_taskOut_TVALID;
	wire [127:0] _peArray_19_taskOut_TDATA;
	wire _peArray_19_taskIn_TREADY;
	wire _peArray_18_closureIn_TREADY;
	wire _peArray_18_argOut_TVALID;
	wire [63:0] _peArray_18_argOut_TDATA;
	wire _peArray_18_taskOut_TVALID;
	wire [127:0] _peArray_18_taskOut_TDATA;
	wire _peArray_18_taskIn_TREADY;
	wire _peArray_17_closureIn_TREADY;
	wire _peArray_17_argOut_TVALID;
	wire [63:0] _peArray_17_argOut_TDATA;
	wire _peArray_17_taskOut_TVALID;
	wire [127:0] _peArray_17_taskOut_TDATA;
	wire _peArray_17_taskIn_TREADY;
	wire _peArray_16_closureIn_TREADY;
	wire _peArray_16_argOut_TVALID;
	wire [63:0] _peArray_16_argOut_TDATA;
	wire _peArray_16_taskOut_TVALID;
	wire [127:0] _peArray_16_taskOut_TDATA;
	wire _peArray_16_taskIn_TREADY;
	wire _peArray_15_closureIn_TREADY;
	wire _peArray_15_argOut_TVALID;
	wire [63:0] _peArray_15_argOut_TDATA;
	wire _peArray_15_taskOut_TVALID;
	wire [127:0] _peArray_15_taskOut_TDATA;
	wire _peArray_15_taskIn_TREADY;
	wire _peArray_14_closureIn_TREADY;
	wire _peArray_14_argOut_TVALID;
	wire [63:0] _peArray_14_argOut_TDATA;
	wire _peArray_14_taskOut_TVALID;
	wire [127:0] _peArray_14_taskOut_TDATA;
	wire _peArray_14_taskIn_TREADY;
	wire _peArray_13_closureIn_TREADY;
	wire _peArray_13_argOut_TVALID;
	wire [63:0] _peArray_13_argOut_TDATA;
	wire _peArray_13_taskOut_TVALID;
	wire [127:0] _peArray_13_taskOut_TDATA;
	wire _peArray_13_taskIn_TREADY;
	wire _peArray_12_closureIn_TREADY;
	wire _peArray_12_argOut_TVALID;
	wire [63:0] _peArray_12_argOut_TDATA;
	wire _peArray_12_taskOut_TVALID;
	wire [127:0] _peArray_12_taskOut_TDATA;
	wire _peArray_12_taskIn_TREADY;
	wire _peArray_11_closureIn_TREADY;
	wire _peArray_11_argOut_TVALID;
	wire [63:0] _peArray_11_argOut_TDATA;
	wire _peArray_11_taskOut_TVALID;
	wire [127:0] _peArray_11_taskOut_TDATA;
	wire _peArray_11_taskIn_TREADY;
	wire _peArray_10_closureIn_TREADY;
	wire _peArray_10_argOut_TVALID;
	wire [63:0] _peArray_10_argOut_TDATA;
	wire _peArray_10_taskOut_TVALID;
	wire [127:0] _peArray_10_taskOut_TDATA;
	wire _peArray_10_taskIn_TREADY;
	wire _peArray_9_closureIn_TREADY;
	wire _peArray_9_argOut_TVALID;
	wire [63:0] _peArray_9_argOut_TDATA;
	wire _peArray_9_taskOut_TVALID;
	wire [127:0] _peArray_9_taskOut_TDATA;
	wire _peArray_9_taskIn_TREADY;
	wire _peArray_8_closureIn_TREADY;
	wire _peArray_8_argOut_TVALID;
	wire [63:0] _peArray_8_argOut_TDATA;
	wire _peArray_8_taskOut_TVALID;
	wire [127:0] _peArray_8_taskOut_TDATA;
	wire _peArray_8_taskIn_TREADY;
	wire _peArray_7_closureIn_TREADY;
	wire _peArray_7_argOut_TVALID;
	wire [63:0] _peArray_7_argOut_TDATA;
	wire _peArray_7_taskOut_TVALID;
	wire [127:0] _peArray_7_taskOut_TDATA;
	wire _peArray_7_taskIn_TREADY;
	wire _peArray_6_closureIn_TREADY;
	wire _peArray_6_argOut_TVALID;
	wire [63:0] _peArray_6_argOut_TDATA;
	wire _peArray_6_taskOut_TVALID;
	wire [127:0] _peArray_6_taskOut_TDATA;
	wire _peArray_6_taskIn_TREADY;
	wire _peArray_5_closureIn_TREADY;
	wire _peArray_5_argOut_TVALID;
	wire [63:0] _peArray_5_argOut_TDATA;
	wire _peArray_5_taskOut_TVALID;
	wire [127:0] _peArray_5_taskOut_TDATA;
	wire _peArray_5_taskIn_TREADY;
	wire _peArray_4_closureIn_TREADY;
	wire _peArray_4_argOut_TVALID;
	wire [63:0] _peArray_4_argOut_TDATA;
	wire _peArray_4_taskOut_TVALID;
	wire [127:0] _peArray_4_taskOut_TDATA;
	wire _peArray_4_taskIn_TREADY;
	wire _peArray_3_closureIn_TREADY;
	wire _peArray_3_argOut_TVALID;
	wire [63:0] _peArray_3_argOut_TDATA;
	wire _peArray_3_taskOut_TVALID;
	wire [127:0] _peArray_3_taskOut_TDATA;
	wire _peArray_3_taskIn_TREADY;
	wire _peArray_2_closureIn_TREADY;
	wire _peArray_2_argOut_TVALID;
	wire [63:0] _peArray_2_argOut_TDATA;
	wire _peArray_2_taskOut_TVALID;
	wire [127:0] _peArray_2_taskOut_TDATA;
	wire _peArray_2_taskIn_TREADY;
	wire _peArray_1_closureIn_TREADY;
	wire _peArray_1_argOut_TVALID;
	wire [63:0] _peArray_1_argOut_TDATA;
	wire _peArray_1_taskOut_TVALID;
	wire [127:0] _peArray_1_taskOut_TDATA;
	wire _peArray_1_taskIn_TREADY;
	wire _peArray_0_closureIn_TREADY;
	wire _peArray_0_argOut_TVALID;
	wire [63:0] _peArray_0_argOut_TDATA;
	wire _peArray_0_taskOut_TVALID;
	wire [127:0] _peArray_0_taskOut_TDATA;
	wire _peArray_0_taskIn_TREADY;
	wire _demux_m_axil_0_ar_valid;
	wire [13:0] _demux_m_axil_0_ar_bits_addr;
	wire [2:0] _demux_m_axil_0_ar_bits_prot;
	wire _demux_m_axil_0_r_ready;
	wire _demux_m_axil_0_aw_valid;
	wire [13:0] _demux_m_axil_0_aw_bits_addr;
	wire [2:0] _demux_m_axil_0_aw_bits_prot;
	wire _demux_m_axil_0_w_valid;
	wire [63:0] _demux_m_axil_0_w_bits_data;
	wire [7:0] _demux_m_axil_0_w_bits_strb;
	wire _demux_m_axil_0_b_ready;
	wire _demux_m_axil_1_ar_valid;
	wire [13:0] _demux_m_axil_1_ar_bits_addr;
	wire [2:0] _demux_m_axil_1_ar_bits_prot;
	wire _demux_m_axil_1_r_ready;
	wire _demux_m_axil_1_aw_valid;
	wire [13:0] _demux_m_axil_1_aw_bits_addr;
	wire [2:0] _demux_m_axil_1_aw_bits_prot;
	wire _demux_m_axil_1_w_valid;
	wire [63:0] _demux_m_axil_1_w_bits_data;
	wire [7:0] _demux_m_axil_1_w_bits_strb;
	wire _demux_m_axil_1_b_ready;
	wire _demux_m_axil_2_ar_valid;
	wire [13:0] _demux_m_axil_2_ar_bits_addr;
	wire [2:0] _demux_m_axil_2_ar_bits_prot;
	wire _demux_m_axil_2_r_ready;
	wire _demux_m_axil_2_aw_valid;
	wire [13:0] _demux_m_axil_2_aw_bits_addr;
	wire [2:0] _demux_m_axil_2_aw_bits_prot;
	wire _demux_m_axil_2_w_valid;
	wire [63:0] _demux_m_axil_2_w_bits_data;
	wire [7:0] _demux_m_axil_2_w_bits_strb;
	wire _demux_m_axil_2_b_ready;
	wire _demux_m_axil_3_ar_valid;
	wire [13:0] _demux_m_axil_3_ar_bits_addr;
	wire [2:0] _demux_m_axil_3_ar_bits_prot;
	wire _demux_m_axil_3_r_ready;
	wire _demux_m_axil_3_aw_valid;
	wire [13:0] _demux_m_axil_3_aw_bits_addr;
	wire [2:0] _demux_m_axil_3_aw_bits_prot;
	wire _demux_m_axil_3_w_valid;
	wire [63:0] _demux_m_axil_3_w_bits_data;
	wire [7:0] _demux_m_axil_3_w_bits_strb;
	wire _demux_m_axil_3_b_ready;
	wire _demux_m_axil_4_ar_valid;
	wire [13:0] _demux_m_axil_4_ar_bits_addr;
	wire [2:0] _demux_m_axil_4_ar_bits_prot;
	wire _demux_m_axil_4_r_ready;
	wire _demux_m_axil_4_aw_valid;
	wire [13:0] _demux_m_axil_4_aw_bits_addr;
	wire [2:0] _demux_m_axil_4_aw_bits_prot;
	wire _demux_m_axil_4_w_valid;
	wire [63:0] _demux_m_axil_4_w_bits_data;
	wire [7:0] _demux_m_axil_4_w_bits_strb;
	wire _demux_m_axil_4_b_ready;
	wire _demux_m_axil_5_ar_valid;
	wire [13:0] _demux_m_axil_5_ar_bits_addr;
	wire [2:0] _demux_m_axil_5_ar_bits_prot;
	wire _demux_m_axil_5_r_ready;
	wire _demux_m_axil_5_aw_valid;
	wire [13:0] _demux_m_axil_5_aw_bits_addr;
	wire [2:0] _demux_m_axil_5_aw_bits_prot;
	wire _demux_m_axil_5_w_valid;
	wire [63:0] _demux_m_axil_5_w_bits_data;
	wire [7:0] _demux_m_axil_5_w_bits_strb;
	wire _demux_m_axil_5_b_ready;
	wire _demux_m_axil_6_ar_valid;
	wire [13:0] _demux_m_axil_6_ar_bits_addr;
	wire [2:0] _demux_m_axil_6_ar_bits_prot;
	wire _demux_m_axil_6_r_ready;
	wire _demux_m_axil_6_aw_valid;
	wire [13:0] _demux_m_axil_6_aw_bits_addr;
	wire [2:0] _demux_m_axil_6_aw_bits_prot;
	wire _demux_m_axil_6_w_valid;
	wire [63:0] _demux_m_axil_6_w_bits_data;
	wire [7:0] _demux_m_axil_6_w_bits_strb;
	wire _demux_m_axil_6_b_ready;
	wire _demux_m_axil_7_ar_valid;
	wire [13:0] _demux_m_axil_7_ar_bits_addr;
	wire [2:0] _demux_m_axil_7_ar_bits_prot;
	wire _demux_m_axil_7_r_ready;
	wire _demux_m_axil_7_aw_valid;
	wire [13:0] _demux_m_axil_7_aw_bits_addr;
	wire [2:0] _demux_m_axil_7_aw_bits_prot;
	wire _demux_m_axil_7_w_valid;
	wire [63:0] _demux_m_axil_7_w_bits_data;
	wire [7:0] _demux_m_axil_7_w_bits_strb;
	wire _demux_m_axil_7_b_ready;
	axi4LiteDemux demux(
		.clock(clock),
		.reset(reset),
		.s_axil_ar_ready(s_axil_mgmt_hardcilk_ARREADY),
		.s_axil_ar_valid(s_axil_mgmt_hardcilk_ARVALID),
		.s_axil_ar_bits_addr(s_axil_mgmt_hardcilk_ARADDR),
		.s_axil_ar_bits_prot(s_axil_mgmt_hardcilk_ARPROT),
		.s_axil_r_ready(s_axil_mgmt_hardcilk_RREADY),
		.s_axil_r_valid(s_axil_mgmt_hardcilk_RVALID),
		.s_axil_r_bits_data(s_axil_mgmt_hardcilk_RDATA),
		.s_axil_r_bits_resp(s_axil_mgmt_hardcilk_RRESP),
		.s_axil_aw_ready(s_axil_mgmt_hardcilk_AWREADY),
		.s_axil_aw_valid(s_axil_mgmt_hardcilk_AWVALID),
		.s_axil_aw_bits_addr(s_axil_mgmt_hardcilk_AWADDR),
		.s_axil_aw_bits_prot(s_axil_mgmt_hardcilk_AWPROT),
		.s_axil_w_ready(s_axil_mgmt_hardcilk_WREADY),
		.s_axil_w_valid(s_axil_mgmt_hardcilk_WVALID),
		.s_axil_w_bits_data(s_axil_mgmt_hardcilk_WDATA),
		.s_axil_w_bits_strb(s_axil_mgmt_hardcilk_WSTRB),
		.s_axil_b_ready(s_axil_mgmt_hardcilk_BREADY),
		.s_axil_b_valid(s_axil_mgmt_hardcilk_BVALID),
		.s_axil_b_bits_resp(s_axil_mgmt_hardcilk_BRESP),
		.m_axil_0_ar_ready(_Scheduler_io_internal_axi_mgmt_vss_0_ar_ready),
		.m_axil_0_ar_valid(_demux_m_axil_0_ar_valid),
		.m_axil_0_ar_bits_addr(_demux_m_axil_0_ar_bits_addr),
		.m_axil_0_ar_bits_prot(_demux_m_axil_0_ar_bits_prot),
		.m_axil_0_r_ready(_demux_m_axil_0_r_ready),
		.m_axil_0_r_valid(_Scheduler_io_internal_axi_mgmt_vss_0_r_valid),
		.m_axil_0_r_bits_data(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_data),
		.m_axil_0_r_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.m_axil_0_aw_ready(_Scheduler_io_internal_axi_mgmt_vss_0_aw_ready),
		.m_axil_0_aw_valid(_demux_m_axil_0_aw_valid),
		.m_axil_0_aw_bits_addr(_demux_m_axil_0_aw_bits_addr),
		.m_axil_0_aw_bits_prot(_demux_m_axil_0_aw_bits_prot),
		.m_axil_0_w_ready(_Scheduler_io_internal_axi_mgmt_vss_0_w_ready),
		.m_axil_0_w_valid(_demux_m_axil_0_w_valid),
		.m_axil_0_w_bits_data(_demux_m_axil_0_w_bits_data),
		.m_axil_0_w_bits_strb(_demux_m_axil_0_w_bits_strb),
		.m_axil_0_b_ready(_demux_m_axil_0_b_ready),
		.m_axil_0_b_valid(_Scheduler_io_internal_axi_mgmt_vss_0_b_valid),
		.m_axil_0_b_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.m_axil_1_ar_ready(_Scheduler_io_internal_axi_mgmt_vss_1_ar_ready),
		.m_axil_1_ar_valid(_demux_m_axil_1_ar_valid),
		.m_axil_1_ar_bits_addr(_demux_m_axil_1_ar_bits_addr),
		.m_axil_1_ar_bits_prot(_demux_m_axil_1_ar_bits_prot),
		.m_axil_1_r_ready(_demux_m_axil_1_r_ready),
		.m_axil_1_r_valid(_Scheduler_io_internal_axi_mgmt_vss_1_r_valid),
		.m_axil_1_r_bits_data(_Scheduler_io_internal_axi_mgmt_vss_1_r_bits_data),
		.m_axil_1_r_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_1_r_bits_resp),
		.m_axil_1_aw_ready(_Scheduler_io_internal_axi_mgmt_vss_1_aw_ready),
		.m_axil_1_aw_valid(_demux_m_axil_1_aw_valid),
		.m_axil_1_aw_bits_addr(_demux_m_axil_1_aw_bits_addr),
		.m_axil_1_aw_bits_prot(_demux_m_axil_1_aw_bits_prot),
		.m_axil_1_w_ready(_Scheduler_io_internal_axi_mgmt_vss_1_w_ready),
		.m_axil_1_w_valid(_demux_m_axil_1_w_valid),
		.m_axil_1_w_bits_data(_demux_m_axil_1_w_bits_data),
		.m_axil_1_w_bits_strb(_demux_m_axil_1_w_bits_strb),
		.m_axil_1_b_ready(_demux_m_axil_1_b_ready),
		.m_axil_1_b_valid(_Scheduler_io_internal_axi_mgmt_vss_1_b_valid),
		.m_axil_1_b_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_1_b_bits_resp),
		.m_axil_2_ar_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_ar_ready),
		.m_axil_2_ar_valid(_demux_m_axil_2_ar_valid),
		.m_axil_2_ar_bits_addr(_demux_m_axil_2_ar_bits_addr),
		.m_axil_2_ar_bits_prot(_demux_m_axil_2_ar_bits_prot),
		.m_axil_2_r_ready(_demux_m_axil_2_r_ready),
		.m_axil_2_r_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_valid),
		.m_axil_2_r_bits_data(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_data),
		.m_axil_2_r_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.m_axil_2_aw_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_aw_ready),
		.m_axil_2_aw_valid(_demux_m_axil_2_aw_valid),
		.m_axil_2_aw_bits_addr(_demux_m_axil_2_aw_bits_addr),
		.m_axil_2_aw_bits_prot(_demux_m_axil_2_aw_bits_prot),
		.m_axil_2_w_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_w_ready),
		.m_axil_2_w_valid(_demux_m_axil_2_w_valid),
		.m_axil_2_w_bits_data(_demux_m_axil_2_w_bits_data),
		.m_axil_2_w_bits_strb(_demux_m_axil_2_w_bits_strb),
		.m_axil_2_b_ready(_demux_m_axil_2_b_ready),
		.m_axil_2_b_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_valid),
		.m_axil_2_b_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.m_axil_3_ar_ready(_Scheduler_1_io_internal_axi_mgmt_vss_1_ar_ready),
		.m_axil_3_ar_valid(_demux_m_axil_3_ar_valid),
		.m_axil_3_ar_bits_addr(_demux_m_axil_3_ar_bits_addr),
		.m_axil_3_ar_bits_prot(_demux_m_axil_3_ar_bits_prot),
		.m_axil_3_r_ready(_demux_m_axil_3_r_ready),
		.m_axil_3_r_valid(_Scheduler_1_io_internal_axi_mgmt_vss_1_r_valid),
		.m_axil_3_r_bits_data(_Scheduler_1_io_internal_axi_mgmt_vss_1_r_bits_data),
		.m_axil_3_r_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_1_r_bits_resp),
		.m_axil_3_aw_ready(_Scheduler_1_io_internal_axi_mgmt_vss_1_aw_ready),
		.m_axil_3_aw_valid(_demux_m_axil_3_aw_valid),
		.m_axil_3_aw_bits_addr(_demux_m_axil_3_aw_bits_addr),
		.m_axil_3_aw_bits_prot(_demux_m_axil_3_aw_bits_prot),
		.m_axil_3_w_ready(_Scheduler_1_io_internal_axi_mgmt_vss_1_w_ready),
		.m_axil_3_w_valid(_demux_m_axil_3_w_valid),
		.m_axil_3_w_bits_data(_demux_m_axil_3_w_bits_data),
		.m_axil_3_w_bits_strb(_demux_m_axil_3_w_bits_strb),
		.m_axil_3_b_ready(_demux_m_axil_3_b_ready),
		.m_axil_3_b_valid(_Scheduler_1_io_internal_axi_mgmt_vss_1_b_valid),
		.m_axil_3_b_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_1_b_bits_resp),
		.m_axil_4_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_0_ar_ready),
		.m_axil_4_ar_valid(_demux_m_axil_4_ar_valid),
		.m_axil_4_ar_bits_addr(_demux_m_axil_4_ar_bits_addr),
		.m_axil_4_ar_bits_prot(_demux_m_axil_4_ar_bits_prot),
		.m_axil_4_r_ready(_demux_m_axil_4_r_ready),
		.m_axil_4_r_valid(_Allocator_io_internal_axi_mgmt_vcas_0_r_valid),
		.m_axil_4_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_data),
		.m_axil_4_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_resp),
		.m_axil_4_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_0_aw_ready),
		.m_axil_4_aw_valid(_demux_m_axil_4_aw_valid),
		.m_axil_4_aw_bits_addr(_demux_m_axil_4_aw_bits_addr),
		.m_axil_4_aw_bits_prot(_demux_m_axil_4_aw_bits_prot),
		.m_axil_4_w_ready(_Allocator_io_internal_axi_mgmt_vcas_0_w_ready),
		.m_axil_4_w_valid(_demux_m_axil_4_w_valid),
		.m_axil_4_w_bits_data(_demux_m_axil_4_w_bits_data),
		.m_axil_4_w_bits_strb(_demux_m_axil_4_w_bits_strb),
		.m_axil_4_b_ready(_demux_m_axil_4_b_ready),
		.m_axil_4_b_valid(_Allocator_io_internal_axi_mgmt_vcas_0_b_valid),
		.m_axil_4_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_b_bits_resp),
		.m_axil_5_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_1_ar_ready),
		.m_axil_5_ar_valid(_demux_m_axil_5_ar_valid),
		.m_axil_5_ar_bits_addr(_demux_m_axil_5_ar_bits_addr),
		.m_axil_5_ar_bits_prot(_demux_m_axil_5_ar_bits_prot),
		.m_axil_5_r_ready(_demux_m_axil_5_r_ready),
		.m_axil_5_r_valid(_Allocator_io_internal_axi_mgmt_vcas_1_r_valid),
		.m_axil_5_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_data),
		.m_axil_5_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_resp),
		.m_axil_5_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_1_aw_ready),
		.m_axil_5_aw_valid(_demux_m_axil_5_aw_valid),
		.m_axil_5_aw_bits_addr(_demux_m_axil_5_aw_bits_addr),
		.m_axil_5_aw_bits_prot(_demux_m_axil_5_aw_bits_prot),
		.m_axil_5_w_ready(_Allocator_io_internal_axi_mgmt_vcas_1_w_ready),
		.m_axil_5_w_valid(_demux_m_axil_5_w_valid),
		.m_axil_5_w_bits_data(_demux_m_axil_5_w_bits_data),
		.m_axil_5_w_bits_strb(_demux_m_axil_5_w_bits_strb),
		.m_axil_5_b_ready(_demux_m_axil_5_b_ready),
		.m_axil_5_b_valid(_Allocator_io_internal_axi_mgmt_vcas_1_b_valid),
		.m_axil_5_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_b_bits_resp),
		.m_axil_6_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_2_ar_ready),
		.m_axil_6_ar_valid(_demux_m_axil_6_ar_valid),
		.m_axil_6_ar_bits_addr(_demux_m_axil_6_ar_bits_addr),
		.m_axil_6_ar_bits_prot(_demux_m_axil_6_ar_bits_prot),
		.m_axil_6_r_ready(_demux_m_axil_6_r_ready),
		.m_axil_6_r_valid(_Allocator_io_internal_axi_mgmt_vcas_2_r_valid),
		.m_axil_6_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_data),
		.m_axil_6_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_resp),
		.m_axil_6_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_2_aw_ready),
		.m_axil_6_aw_valid(_demux_m_axil_6_aw_valid),
		.m_axil_6_aw_bits_addr(_demux_m_axil_6_aw_bits_addr),
		.m_axil_6_aw_bits_prot(_demux_m_axil_6_aw_bits_prot),
		.m_axil_6_w_ready(_Allocator_io_internal_axi_mgmt_vcas_2_w_ready),
		.m_axil_6_w_valid(_demux_m_axil_6_w_valid),
		.m_axil_6_w_bits_data(_demux_m_axil_6_w_bits_data),
		.m_axil_6_w_bits_strb(_demux_m_axil_6_w_bits_strb),
		.m_axil_6_b_ready(_demux_m_axil_6_b_ready),
		.m_axil_6_b_valid(_Allocator_io_internal_axi_mgmt_vcas_2_b_valid),
		.m_axil_6_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_b_bits_resp),
		.m_axil_7_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_3_ar_ready),
		.m_axil_7_ar_valid(_demux_m_axil_7_ar_valid),
		.m_axil_7_ar_bits_addr(_demux_m_axil_7_ar_bits_addr),
		.m_axil_7_ar_bits_prot(_demux_m_axil_7_ar_bits_prot),
		.m_axil_7_r_ready(_demux_m_axil_7_r_ready),
		.m_axil_7_r_valid(_Allocator_io_internal_axi_mgmt_vcas_3_r_valid),
		.m_axil_7_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_data),
		.m_axil_7_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_resp),
		.m_axil_7_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_3_aw_ready),
		.m_axil_7_aw_valid(_demux_m_axil_7_aw_valid),
		.m_axil_7_aw_bits_addr(_demux_m_axil_7_aw_bits_addr),
		.m_axil_7_aw_bits_prot(_demux_m_axil_7_aw_bits_prot),
		.m_axil_7_w_ready(_Allocator_io_internal_axi_mgmt_vcas_3_w_ready),
		.m_axil_7_w_valid(_demux_m_axil_7_w_valid),
		.m_axil_7_w_bits_data(_demux_m_axil_7_w_bits_data),
		.m_axil_7_w_bits_strb(_demux_m_axil_7_w_bits_strb),
		.m_axil_7_b_ready(_demux_m_axil_7_b_ready),
		.m_axil_7_b_valid(_Allocator_io_internal_axi_mgmt_vcas_3_b_valid),
		.m_axil_7_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_b_bits_resp)
	);
	fib peArray_0(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_0_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_0_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_0_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_0_TREADY),
		.argOut_TVALID(_peArray_0_argOut_TVALID),
		.argOut_TDATA(_peArray_0_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_0_TREADY),
		.taskOut_TVALID(_peArray_0_taskOut_TVALID),
		.taskOut_TDATA(_peArray_0_taskOut_TDATA),
		.taskIn_TREADY(_peArray_0_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_0_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_0_TDATA),
		.s_axi_control_ARREADY(fib_0_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_0_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_0_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_0_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_0_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_0_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_0_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_0_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_0_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_0_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_0_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_0_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_0_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_0_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_0_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_0_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_0_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_0_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_0_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_0_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_0_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_0_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_0_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_0_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_0_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_0_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_0_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_0_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_0_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_0_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_0_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_0_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_0_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_0_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_0_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_0_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_0_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_0_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_0_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_0_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_0_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_0_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_0_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_0_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_0_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_0_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_0_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_0_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_0_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_0_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_0_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_0_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_0_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_0_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_0_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_0_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_0_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_0_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_0_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_0_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_0_m_axi_gmem_BUSER)
	);
	fib peArray_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_1_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_1_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_1_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_1_TREADY),
		.argOut_TVALID(_peArray_1_argOut_TVALID),
		.argOut_TDATA(_peArray_1_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_1_TREADY),
		.taskOut_TVALID(_peArray_1_taskOut_TVALID),
		.taskOut_TDATA(_peArray_1_taskOut_TDATA),
		.taskIn_TREADY(_peArray_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_1_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_1_TDATA),
		.s_axi_control_ARREADY(fib_1_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_1_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_1_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_1_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_1_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_1_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_1_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_1_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_1_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_1_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_1_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_1_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_1_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_1_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_1_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_1_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_1_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_1_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_1_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_1_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_1_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_1_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_1_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_1_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_1_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_1_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_1_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_1_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_1_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_1_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_1_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_1_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_1_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_1_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_1_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_1_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_1_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_1_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_1_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_1_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_1_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_1_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_1_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_1_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_1_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_1_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_1_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_1_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_1_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_1_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_1_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_1_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_1_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_1_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_1_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_1_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_1_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_1_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_1_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_1_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_1_m_axi_gmem_BUSER)
	);
	fib peArray_2(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_2_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_2_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_2_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_2_TREADY),
		.argOut_TVALID(_peArray_2_argOut_TVALID),
		.argOut_TDATA(_peArray_2_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_2_TREADY),
		.taskOut_TVALID(_peArray_2_taskOut_TVALID),
		.taskOut_TDATA(_peArray_2_taskOut_TDATA),
		.taskIn_TREADY(_peArray_2_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_2_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_2_TDATA),
		.s_axi_control_ARREADY(fib_2_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_2_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_2_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_2_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_2_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_2_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_2_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_2_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_2_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_2_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_2_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_2_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_2_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_2_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_2_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_2_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_2_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_2_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_2_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_2_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_2_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_2_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_2_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_2_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_2_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_2_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_2_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_2_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_2_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_2_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_2_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_2_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_2_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_2_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_2_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_2_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_2_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_2_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_2_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_2_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_2_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_2_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_2_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_2_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_2_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_2_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_2_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_2_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_2_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_2_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_2_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_2_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_2_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_2_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_2_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_2_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_2_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_2_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_2_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_2_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_2_m_axi_gmem_BUSER)
	);
	fib peArray_3(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_3_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_3_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_3_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_3_TREADY),
		.argOut_TVALID(_peArray_3_argOut_TVALID),
		.argOut_TDATA(_peArray_3_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_3_TREADY),
		.taskOut_TVALID(_peArray_3_taskOut_TVALID),
		.taskOut_TDATA(_peArray_3_taskOut_TDATA),
		.taskIn_TREADY(_peArray_3_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_3_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_3_TDATA),
		.s_axi_control_ARREADY(fib_3_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_3_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_3_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_3_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_3_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_3_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_3_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_3_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_3_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_3_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_3_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_3_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_3_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_3_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_3_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_3_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_3_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_3_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_3_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_3_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_3_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_3_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_3_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_3_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_3_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_3_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_3_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_3_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_3_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_3_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_3_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_3_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_3_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_3_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_3_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_3_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_3_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_3_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_3_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_3_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_3_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_3_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_3_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_3_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_3_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_3_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_3_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_3_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_3_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_3_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_3_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_3_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_3_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_3_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_3_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_3_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_3_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_3_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_3_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_3_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_3_m_axi_gmem_BUSER)
	);
	fib peArray_4(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_4_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_4_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_4_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_4_TREADY),
		.argOut_TVALID(_peArray_4_argOut_TVALID),
		.argOut_TDATA(_peArray_4_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_4_TREADY),
		.taskOut_TVALID(_peArray_4_taskOut_TVALID),
		.taskOut_TDATA(_peArray_4_taskOut_TDATA),
		.taskIn_TREADY(_peArray_4_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_4_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_4_TDATA),
		.s_axi_control_ARREADY(fib_4_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_4_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_4_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_4_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_4_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_4_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_4_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_4_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_4_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_4_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_4_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_4_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_4_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_4_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_4_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_4_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_4_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_4_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_4_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_4_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_4_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_4_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_4_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_4_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_4_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_4_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_4_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_4_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_4_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_4_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_4_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_4_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_4_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_4_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_4_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_4_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_4_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_4_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_4_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_4_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_4_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_4_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_4_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_4_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_4_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_4_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_4_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_4_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_4_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_4_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_4_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_4_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_4_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_4_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_4_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_4_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_4_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_4_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_4_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_4_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_4_m_axi_gmem_BUSER)
	);
	fib peArray_5(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_5_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_5_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_5_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_5_TREADY),
		.argOut_TVALID(_peArray_5_argOut_TVALID),
		.argOut_TDATA(_peArray_5_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_5_TREADY),
		.taskOut_TVALID(_peArray_5_taskOut_TVALID),
		.taskOut_TDATA(_peArray_5_taskOut_TDATA),
		.taskIn_TREADY(_peArray_5_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_5_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_5_TDATA),
		.s_axi_control_ARREADY(fib_5_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_5_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_5_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_5_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_5_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_5_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_5_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_5_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_5_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_5_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_5_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_5_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_5_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_5_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_5_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_5_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_5_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_5_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_5_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_5_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_5_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_5_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_5_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_5_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_5_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_5_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_5_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_5_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_5_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_5_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_5_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_5_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_5_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_5_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_5_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_5_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_5_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_5_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_5_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_5_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_5_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_5_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_5_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_5_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_5_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_5_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_5_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_5_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_5_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_5_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_5_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_5_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_5_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_5_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_5_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_5_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_5_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_5_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_5_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_5_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_5_m_axi_gmem_BUSER)
	);
	fib peArray_6(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_6_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_6_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_6_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_6_TREADY),
		.argOut_TVALID(_peArray_6_argOut_TVALID),
		.argOut_TDATA(_peArray_6_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_6_TREADY),
		.taskOut_TVALID(_peArray_6_taskOut_TVALID),
		.taskOut_TDATA(_peArray_6_taskOut_TDATA),
		.taskIn_TREADY(_peArray_6_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_6_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_6_TDATA),
		.s_axi_control_ARREADY(fib_6_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_6_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_6_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_6_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_6_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_6_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_6_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_6_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_6_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_6_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_6_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_6_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_6_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_6_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_6_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_6_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_6_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_6_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_6_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_6_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_6_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_6_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_6_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_6_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_6_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_6_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_6_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_6_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_6_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_6_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_6_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_6_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_6_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_6_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_6_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_6_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_6_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_6_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_6_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_6_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_6_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_6_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_6_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_6_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_6_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_6_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_6_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_6_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_6_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_6_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_6_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_6_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_6_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_6_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_6_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_6_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_6_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_6_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_6_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_6_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_6_m_axi_gmem_BUSER)
	);
	fib peArray_7(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_7_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_7_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_7_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_7_TREADY),
		.argOut_TVALID(_peArray_7_argOut_TVALID),
		.argOut_TDATA(_peArray_7_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_7_TREADY),
		.taskOut_TVALID(_peArray_7_taskOut_TVALID),
		.taskOut_TDATA(_peArray_7_taskOut_TDATA),
		.taskIn_TREADY(_peArray_7_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_7_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_7_TDATA),
		.s_axi_control_ARREADY(fib_7_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_7_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_7_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_7_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_7_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_7_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_7_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_7_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_7_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_7_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_7_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_7_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_7_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_7_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_7_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_7_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_7_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_7_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_7_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_7_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_7_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_7_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_7_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_7_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_7_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_7_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_7_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_7_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_7_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_7_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_7_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_7_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_7_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_7_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_7_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_7_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_7_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_7_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_7_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_7_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_7_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_7_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_7_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_7_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_7_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_7_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_7_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_7_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_7_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_7_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_7_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_7_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_7_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_7_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_7_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_7_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_7_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_7_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_7_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_7_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_7_m_axi_gmem_BUSER)
	);
	fib peArray_8(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_8_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_8_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_8_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_8_TREADY),
		.argOut_TVALID(_peArray_8_argOut_TVALID),
		.argOut_TDATA(_peArray_8_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_8_TREADY),
		.taskOut_TVALID(_peArray_8_taskOut_TVALID),
		.taskOut_TDATA(_peArray_8_taskOut_TDATA),
		.taskIn_TREADY(_peArray_8_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_8_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_8_TDATA),
		.s_axi_control_ARREADY(fib_8_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_8_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_8_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_8_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_8_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_8_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_8_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_8_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_8_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_8_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_8_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_8_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_8_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_8_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_8_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_8_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_8_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_8_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_8_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_8_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_8_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_8_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_8_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_8_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_8_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_8_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_8_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_8_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_8_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_8_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_8_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_8_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_8_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_8_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_8_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_8_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_8_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_8_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_8_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_8_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_8_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_8_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_8_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_8_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_8_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_8_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_8_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_8_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_8_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_8_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_8_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_8_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_8_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_8_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_8_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_8_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_8_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_8_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_8_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_8_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_8_m_axi_gmem_BUSER)
	);
	fib peArray_9(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_9_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_9_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_9_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_9_TREADY),
		.argOut_TVALID(_peArray_9_argOut_TVALID),
		.argOut_TDATA(_peArray_9_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_9_TREADY),
		.taskOut_TVALID(_peArray_9_taskOut_TVALID),
		.taskOut_TDATA(_peArray_9_taskOut_TDATA),
		.taskIn_TREADY(_peArray_9_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_9_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_9_TDATA),
		.s_axi_control_ARREADY(fib_9_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_9_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_9_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_9_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_9_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_9_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_9_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_9_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_9_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_9_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_9_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_9_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_9_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_9_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_9_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_9_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_9_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_9_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_9_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_9_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_9_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_9_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_9_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_9_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_9_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_9_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_9_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_9_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_9_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_9_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_9_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_9_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_9_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_9_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_9_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_9_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_9_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_9_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_9_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_9_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_9_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_9_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_9_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_9_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_9_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_9_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_9_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_9_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_9_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_9_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_9_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_9_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_9_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_9_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_9_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_9_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_9_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_9_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_9_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_9_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_9_m_axi_gmem_BUSER)
	);
	fib peArray_10(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_10_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_10_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_10_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_10_TREADY),
		.argOut_TVALID(_peArray_10_argOut_TVALID),
		.argOut_TDATA(_peArray_10_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_10_TREADY),
		.taskOut_TVALID(_peArray_10_taskOut_TVALID),
		.taskOut_TDATA(_peArray_10_taskOut_TDATA),
		.taskIn_TREADY(_peArray_10_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_10_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_10_TDATA),
		.s_axi_control_ARREADY(fib_10_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_10_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_10_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_10_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_10_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_10_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_10_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_10_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_10_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_10_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_10_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_10_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_10_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_10_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_10_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_10_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_10_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_10_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_10_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_10_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_10_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_10_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_10_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_10_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_10_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_10_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_10_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_10_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_10_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_10_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_10_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_10_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_10_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_10_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_10_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_10_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_10_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_10_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_10_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_10_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_10_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_10_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_10_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_10_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_10_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_10_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_10_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_10_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_10_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_10_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_10_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_10_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_10_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_10_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_10_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_10_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_10_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_10_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_10_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_10_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_10_m_axi_gmem_BUSER)
	);
	fib peArray_11(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_11_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_11_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_11_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_11_TREADY),
		.argOut_TVALID(_peArray_11_argOut_TVALID),
		.argOut_TDATA(_peArray_11_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_11_TREADY),
		.taskOut_TVALID(_peArray_11_taskOut_TVALID),
		.taskOut_TDATA(_peArray_11_taskOut_TDATA),
		.taskIn_TREADY(_peArray_11_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_11_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_11_TDATA),
		.s_axi_control_ARREADY(fib_11_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_11_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_11_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_11_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_11_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_11_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_11_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_11_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_11_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_11_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_11_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_11_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_11_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_11_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_11_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_11_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_11_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_11_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_11_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_11_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_11_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_11_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_11_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_11_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_11_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_11_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_11_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_11_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_11_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_11_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_11_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_11_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_11_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_11_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_11_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_11_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_11_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_11_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_11_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_11_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_11_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_11_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_11_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_11_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_11_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_11_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_11_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_11_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_11_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_11_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_11_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_11_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_11_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_11_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_11_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_11_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_11_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_11_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_11_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_11_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_11_m_axi_gmem_BUSER)
	);
	fib peArray_12(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_12_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_12_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_12_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_12_TREADY),
		.argOut_TVALID(_peArray_12_argOut_TVALID),
		.argOut_TDATA(_peArray_12_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_12_TREADY),
		.taskOut_TVALID(_peArray_12_taskOut_TVALID),
		.taskOut_TDATA(_peArray_12_taskOut_TDATA),
		.taskIn_TREADY(_peArray_12_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_12_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_12_TDATA),
		.s_axi_control_ARREADY(fib_12_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_12_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_12_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_12_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_12_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_12_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_12_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_12_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_12_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_12_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_12_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_12_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_12_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_12_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_12_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_12_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_12_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_12_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_12_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_12_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_12_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_12_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_12_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_12_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_12_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_12_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_12_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_12_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_12_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_12_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_12_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_12_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_12_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_12_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_12_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_12_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_12_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_12_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_12_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_12_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_12_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_12_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_12_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_12_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_12_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_12_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_12_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_12_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_12_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_12_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_12_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_12_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_12_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_12_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_12_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_12_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_12_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_12_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_12_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_12_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_12_m_axi_gmem_BUSER)
	);
	fib peArray_13(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_13_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_13_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_13_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_13_TREADY),
		.argOut_TVALID(_peArray_13_argOut_TVALID),
		.argOut_TDATA(_peArray_13_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_13_TREADY),
		.taskOut_TVALID(_peArray_13_taskOut_TVALID),
		.taskOut_TDATA(_peArray_13_taskOut_TDATA),
		.taskIn_TREADY(_peArray_13_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_13_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_13_TDATA),
		.s_axi_control_ARREADY(fib_13_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_13_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_13_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_13_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_13_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_13_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_13_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_13_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_13_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_13_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_13_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_13_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_13_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_13_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_13_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_13_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_13_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_13_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_13_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_13_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_13_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_13_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_13_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_13_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_13_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_13_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_13_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_13_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_13_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_13_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_13_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_13_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_13_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_13_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_13_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_13_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_13_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_13_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_13_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_13_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_13_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_13_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_13_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_13_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_13_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_13_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_13_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_13_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_13_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_13_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_13_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_13_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_13_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_13_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_13_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_13_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_13_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_13_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_13_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_13_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_13_m_axi_gmem_BUSER)
	);
	fib peArray_14(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_14_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_14_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_14_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_14_TREADY),
		.argOut_TVALID(_peArray_14_argOut_TVALID),
		.argOut_TDATA(_peArray_14_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_14_TREADY),
		.taskOut_TVALID(_peArray_14_taskOut_TVALID),
		.taskOut_TDATA(_peArray_14_taskOut_TDATA),
		.taskIn_TREADY(_peArray_14_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_14_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_14_TDATA),
		.s_axi_control_ARREADY(fib_14_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_14_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_14_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_14_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_14_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_14_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_14_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_14_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_14_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_14_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_14_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_14_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_14_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_14_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_14_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_14_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_14_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_14_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_14_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_14_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_14_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_14_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_14_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_14_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_14_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_14_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_14_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_14_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_14_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_14_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_14_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_14_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_14_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_14_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_14_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_14_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_14_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_14_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_14_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_14_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_14_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_14_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_14_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_14_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_14_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_14_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_14_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_14_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_14_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_14_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_14_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_14_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_14_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_14_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_14_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_14_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_14_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_14_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_14_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_14_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_14_m_axi_gmem_BUSER)
	);
	fib peArray_15(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_15_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_15_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_15_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_15_TREADY),
		.argOut_TVALID(_peArray_15_argOut_TVALID),
		.argOut_TDATA(_peArray_15_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_15_TREADY),
		.taskOut_TVALID(_peArray_15_taskOut_TVALID),
		.taskOut_TDATA(_peArray_15_taskOut_TDATA),
		.taskIn_TREADY(_peArray_15_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_15_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_15_TDATA),
		.s_axi_control_ARREADY(fib_15_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_15_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_15_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_15_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_15_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_15_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_15_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_15_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_15_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_15_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_15_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_15_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_15_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_15_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_15_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_15_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_15_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_15_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_15_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_15_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_15_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_15_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_15_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_15_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_15_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_15_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_15_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_15_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_15_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_15_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_15_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_15_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_15_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_15_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_15_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_15_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_15_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_15_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_15_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_15_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_15_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_15_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_15_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_15_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_15_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_15_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_15_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_15_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_15_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_15_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_15_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_15_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_15_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_15_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_15_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_15_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_15_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_15_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_15_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_15_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_15_m_axi_gmem_BUSER)
	);
	fib peArray_16(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_16_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_16_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_16_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_16_TREADY),
		.argOut_TVALID(_peArray_16_argOut_TVALID),
		.argOut_TDATA(_peArray_16_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_16_TREADY),
		.taskOut_TVALID(_peArray_16_taskOut_TVALID),
		.taskOut_TDATA(_peArray_16_taskOut_TDATA),
		.taskIn_TREADY(_peArray_16_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_16_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_16_TDATA),
		.s_axi_control_ARREADY(fib_16_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_16_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_16_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_16_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_16_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_16_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_16_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_16_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_16_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_16_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_16_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_16_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_16_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_16_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_16_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_16_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_16_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_16_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_16_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_16_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_16_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_16_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_16_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_16_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_16_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_16_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_16_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_16_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_16_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_16_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_16_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_16_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_16_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_16_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_16_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_16_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_16_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_16_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_16_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_16_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_16_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_16_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_16_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_16_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_16_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_16_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_16_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_16_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_16_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_16_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_16_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_16_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_16_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_16_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_16_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_16_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_16_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_16_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_16_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_16_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_16_m_axi_gmem_BUSER)
	);
	fib peArray_17(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_17_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_17_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_17_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_17_TREADY),
		.argOut_TVALID(_peArray_17_argOut_TVALID),
		.argOut_TDATA(_peArray_17_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_17_TREADY),
		.taskOut_TVALID(_peArray_17_taskOut_TVALID),
		.taskOut_TDATA(_peArray_17_taskOut_TDATA),
		.taskIn_TREADY(_peArray_17_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_17_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_17_TDATA),
		.s_axi_control_ARREADY(fib_17_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_17_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_17_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_17_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_17_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_17_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_17_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_17_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_17_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_17_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_17_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_17_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_17_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_17_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_17_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_17_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_17_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_17_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_17_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_17_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_17_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_17_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_17_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_17_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_17_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_17_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_17_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_17_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_17_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_17_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_17_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_17_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_17_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_17_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_17_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_17_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_17_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_17_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_17_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_17_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_17_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_17_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_17_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_17_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_17_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_17_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_17_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_17_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_17_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_17_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_17_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_17_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_17_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_17_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_17_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_17_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_17_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_17_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_17_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_17_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_17_m_axi_gmem_BUSER)
	);
	fib peArray_18(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_18_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_18_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_18_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_18_TREADY),
		.argOut_TVALID(_peArray_18_argOut_TVALID),
		.argOut_TDATA(_peArray_18_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_18_TREADY),
		.taskOut_TVALID(_peArray_18_taskOut_TVALID),
		.taskOut_TDATA(_peArray_18_taskOut_TDATA),
		.taskIn_TREADY(_peArray_18_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_18_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_18_TDATA),
		.s_axi_control_ARREADY(fib_18_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_18_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_18_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_18_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_18_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_18_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_18_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_18_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_18_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_18_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_18_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_18_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_18_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_18_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_18_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_18_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_18_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_18_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_18_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_18_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_18_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_18_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_18_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_18_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_18_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_18_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_18_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_18_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_18_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_18_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_18_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_18_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_18_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_18_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_18_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_18_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_18_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_18_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_18_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_18_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_18_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_18_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_18_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_18_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_18_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_18_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_18_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_18_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_18_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_18_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_18_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_18_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_18_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_18_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_18_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_18_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_18_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_18_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_18_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_18_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_18_m_axi_gmem_BUSER)
	);
	fib peArray_19(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_19_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_19_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_19_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_19_TREADY),
		.argOut_TVALID(_peArray_19_argOut_TVALID),
		.argOut_TDATA(_peArray_19_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_19_TREADY),
		.taskOut_TVALID(_peArray_19_taskOut_TVALID),
		.taskOut_TDATA(_peArray_19_taskOut_TDATA),
		.taskIn_TREADY(_peArray_19_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_19_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_19_TDATA),
		.s_axi_control_ARREADY(fib_19_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_19_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_19_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_19_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_19_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_19_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_19_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_19_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_19_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_19_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_19_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_19_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_19_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_19_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_19_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_19_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_19_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_19_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_19_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_19_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_19_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_19_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_19_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_19_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_19_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_19_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_19_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_19_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_19_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_19_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_19_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_19_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_19_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_19_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_19_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_19_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_19_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_19_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_19_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_19_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_19_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_19_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_19_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_19_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_19_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_19_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_19_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_19_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_19_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_19_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_19_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_19_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_19_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_19_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_19_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_19_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_19_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_19_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_19_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_19_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_19_m_axi_gmem_BUSER)
	);
	fib peArray_20(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_20_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_20_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_20_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_20_TREADY),
		.argOut_TVALID(_peArray_20_argOut_TVALID),
		.argOut_TDATA(_peArray_20_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_20_TREADY),
		.taskOut_TVALID(_peArray_20_taskOut_TVALID),
		.taskOut_TDATA(_peArray_20_taskOut_TDATA),
		.taskIn_TREADY(_peArray_20_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_20_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_20_TDATA),
		.s_axi_control_ARREADY(fib_20_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_20_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_20_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_20_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_20_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_20_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_20_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_20_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_20_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_20_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_20_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_20_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_20_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_20_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_20_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_20_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_20_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_20_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_20_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_20_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_20_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_20_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_20_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_20_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_20_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_20_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_20_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_20_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_20_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_20_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_20_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_20_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_20_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_20_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_20_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_20_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_20_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_20_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_20_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_20_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_20_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_20_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_20_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_20_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_20_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_20_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_20_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_20_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_20_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_20_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_20_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_20_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_20_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_20_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_20_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_20_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_20_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_20_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_20_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_20_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_20_m_axi_gmem_BUSER)
	);
	fib peArray_21(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_21_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_21_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_21_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_21_TREADY),
		.argOut_TVALID(_peArray_21_argOut_TVALID),
		.argOut_TDATA(_peArray_21_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_21_TREADY),
		.taskOut_TVALID(_peArray_21_taskOut_TVALID),
		.taskOut_TDATA(_peArray_21_taskOut_TDATA),
		.taskIn_TREADY(_peArray_21_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_21_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_21_TDATA),
		.s_axi_control_ARREADY(fib_21_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_21_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_21_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_21_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_21_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_21_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_21_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_21_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_21_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_21_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_21_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_21_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_21_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_21_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_21_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_21_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_21_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_21_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_21_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_21_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_21_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_21_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_21_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_21_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_21_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_21_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_21_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_21_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_21_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_21_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_21_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_21_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_21_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_21_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_21_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_21_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_21_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_21_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_21_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_21_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_21_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_21_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_21_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_21_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_21_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_21_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_21_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_21_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_21_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_21_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_21_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_21_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_21_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_21_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_21_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_21_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_21_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_21_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_21_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_21_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_21_m_axi_gmem_BUSER)
	);
	fib peArray_22(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_22_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_22_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_22_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_22_TREADY),
		.argOut_TVALID(_peArray_22_argOut_TVALID),
		.argOut_TDATA(_peArray_22_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_22_TREADY),
		.taskOut_TVALID(_peArray_22_taskOut_TVALID),
		.taskOut_TDATA(_peArray_22_taskOut_TDATA),
		.taskIn_TREADY(_peArray_22_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_22_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_22_TDATA),
		.s_axi_control_ARREADY(fib_22_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_22_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_22_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_22_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_22_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_22_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_22_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_22_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_22_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_22_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_22_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_22_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_22_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_22_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_22_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_22_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_22_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_22_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_22_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_22_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_22_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_22_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_22_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_22_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_22_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_22_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_22_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_22_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_22_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_22_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_22_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_22_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_22_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_22_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_22_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_22_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_22_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_22_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_22_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_22_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_22_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_22_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_22_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_22_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_22_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_22_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_22_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_22_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_22_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_22_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_22_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_22_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_22_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_22_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_22_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_22_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_22_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_22_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_22_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_22_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_22_m_axi_gmem_BUSER)
	);
	fib peArray_23(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_23_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_23_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_23_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_23_TREADY),
		.argOut_TVALID(_peArray_23_argOut_TVALID),
		.argOut_TDATA(_peArray_23_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_23_TREADY),
		.taskOut_TVALID(_peArray_23_taskOut_TVALID),
		.taskOut_TDATA(_peArray_23_taskOut_TDATA),
		.taskIn_TREADY(_peArray_23_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_23_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_23_TDATA),
		.s_axi_control_ARREADY(fib_23_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_23_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_23_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_23_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_23_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_23_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_23_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_23_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_23_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_23_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_23_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_23_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_23_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_23_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_23_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_23_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_23_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_23_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_23_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_23_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_23_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_23_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_23_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_23_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_23_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_23_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_23_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_23_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_23_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_23_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_23_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_23_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_23_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_23_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_23_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_23_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_23_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_23_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_23_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_23_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_23_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_23_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_23_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_23_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_23_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_23_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_23_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_23_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_23_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_23_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_23_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_23_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_23_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_23_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_23_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_23_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_23_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_23_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_23_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_23_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_23_m_axi_gmem_BUSER)
	);
	fib peArray_24(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_24_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_24_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_24_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_24_TREADY),
		.argOut_TVALID(_peArray_24_argOut_TVALID),
		.argOut_TDATA(_peArray_24_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_24_TREADY),
		.taskOut_TVALID(_peArray_24_taskOut_TVALID),
		.taskOut_TDATA(_peArray_24_taskOut_TDATA),
		.taskIn_TREADY(_peArray_24_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_24_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_24_TDATA),
		.s_axi_control_ARREADY(fib_24_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_24_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_24_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_24_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_24_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_24_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_24_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_24_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_24_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_24_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_24_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_24_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_24_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_24_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_24_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_24_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_24_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_24_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_24_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_24_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_24_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_24_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_24_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_24_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_24_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_24_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_24_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_24_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_24_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_24_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_24_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_24_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_24_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_24_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_24_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_24_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_24_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_24_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_24_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_24_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_24_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_24_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_24_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_24_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_24_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_24_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_24_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_24_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_24_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_24_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_24_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_24_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_24_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_24_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_24_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_24_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_24_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_24_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_24_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_24_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_24_m_axi_gmem_BUSER)
	);
	fib peArray_25(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_25_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_25_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_25_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_25_TREADY),
		.argOut_TVALID(_peArray_25_argOut_TVALID),
		.argOut_TDATA(_peArray_25_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_25_TREADY),
		.taskOut_TVALID(_peArray_25_taskOut_TVALID),
		.taskOut_TDATA(_peArray_25_taskOut_TDATA),
		.taskIn_TREADY(_peArray_25_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_25_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_25_TDATA),
		.s_axi_control_ARREADY(fib_25_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_25_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_25_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_25_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_25_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_25_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_25_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_25_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_25_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_25_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_25_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_25_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_25_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_25_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_25_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_25_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_25_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_25_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_25_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_25_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_25_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_25_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_25_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_25_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_25_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_25_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_25_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_25_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_25_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_25_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_25_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_25_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_25_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_25_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_25_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_25_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_25_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_25_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_25_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_25_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_25_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_25_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_25_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_25_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_25_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_25_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_25_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_25_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_25_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_25_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_25_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_25_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_25_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_25_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_25_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_25_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_25_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_25_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_25_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_25_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_25_m_axi_gmem_BUSER)
	);
	fib peArray_26(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_26_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_26_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_26_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_26_TREADY),
		.argOut_TVALID(_peArray_26_argOut_TVALID),
		.argOut_TDATA(_peArray_26_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_26_TREADY),
		.taskOut_TVALID(_peArray_26_taskOut_TVALID),
		.taskOut_TDATA(_peArray_26_taskOut_TDATA),
		.taskIn_TREADY(_peArray_26_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_26_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_26_TDATA),
		.s_axi_control_ARREADY(fib_26_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_26_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_26_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_26_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_26_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_26_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_26_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_26_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_26_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_26_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_26_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_26_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_26_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_26_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_26_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_26_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_26_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_26_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_26_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_26_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_26_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_26_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_26_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_26_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_26_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_26_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_26_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_26_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_26_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_26_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_26_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_26_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_26_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_26_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_26_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_26_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_26_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_26_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_26_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_26_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_26_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_26_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_26_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_26_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_26_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_26_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_26_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_26_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_26_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_26_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_26_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_26_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_26_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_26_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_26_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_26_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_26_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_26_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_26_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_26_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_26_m_axi_gmem_BUSER)
	);
	fib peArray_27(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_27_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_27_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_27_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_27_TREADY),
		.argOut_TVALID(_peArray_27_argOut_TVALID),
		.argOut_TDATA(_peArray_27_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_27_TREADY),
		.taskOut_TVALID(_peArray_27_taskOut_TVALID),
		.taskOut_TDATA(_peArray_27_taskOut_TDATA),
		.taskIn_TREADY(_peArray_27_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_27_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_27_TDATA),
		.s_axi_control_ARREADY(fib_27_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_27_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_27_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_27_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_27_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_27_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_27_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_27_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_27_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_27_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_27_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_27_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_27_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_27_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_27_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_27_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_27_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_27_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_27_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_27_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_27_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_27_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_27_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_27_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_27_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_27_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_27_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_27_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_27_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_27_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_27_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_27_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_27_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_27_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_27_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_27_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_27_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_27_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_27_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_27_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_27_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_27_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_27_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_27_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_27_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_27_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_27_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_27_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_27_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_27_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_27_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_27_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_27_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_27_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_27_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_27_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_27_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_27_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_27_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_27_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_27_m_axi_gmem_BUSER)
	);
	fib peArray_28(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_28_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_28_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_28_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_28_TREADY),
		.argOut_TVALID(_peArray_28_argOut_TVALID),
		.argOut_TDATA(_peArray_28_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_28_TREADY),
		.taskOut_TVALID(_peArray_28_taskOut_TVALID),
		.taskOut_TDATA(_peArray_28_taskOut_TDATA),
		.taskIn_TREADY(_peArray_28_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_28_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_28_TDATA),
		.s_axi_control_ARREADY(fib_28_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_28_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_28_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_28_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_28_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_28_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_28_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_28_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_28_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_28_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_28_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_28_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_28_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_28_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_28_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_28_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_28_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_28_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_28_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_28_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_28_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_28_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_28_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_28_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_28_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_28_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_28_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_28_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_28_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_28_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_28_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_28_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_28_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_28_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_28_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_28_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_28_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_28_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_28_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_28_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_28_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_28_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_28_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_28_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_28_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_28_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_28_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_28_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_28_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_28_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_28_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_28_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_28_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_28_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_28_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_28_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_28_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_28_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_28_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_28_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_28_m_axi_gmem_BUSER)
	);
	fib peArray_29(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_29_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_29_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_29_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_29_TREADY),
		.argOut_TVALID(_peArray_29_argOut_TVALID),
		.argOut_TDATA(_peArray_29_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_29_TREADY),
		.taskOut_TVALID(_peArray_29_taskOut_TVALID),
		.taskOut_TDATA(_peArray_29_taskOut_TDATA),
		.taskIn_TREADY(_peArray_29_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_29_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_29_TDATA),
		.s_axi_control_ARREADY(fib_29_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_29_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_29_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_29_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_29_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_29_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_29_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_29_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_29_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_29_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_29_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_29_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_29_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_29_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_29_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_29_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_29_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_29_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_29_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_29_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_29_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_29_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_29_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_29_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_29_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_29_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_29_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_29_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_29_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_29_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_29_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_29_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_29_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_29_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_29_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_29_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_29_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_29_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_29_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_29_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_29_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_29_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_29_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_29_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_29_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_29_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_29_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_29_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_29_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_29_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_29_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_29_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_29_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_29_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_29_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_29_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_29_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_29_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_29_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_29_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_29_m_axi_gmem_BUSER)
	);
	fib peArray_30(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_30_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_30_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_30_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_30_TREADY),
		.argOut_TVALID(_peArray_30_argOut_TVALID),
		.argOut_TDATA(_peArray_30_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_30_TREADY),
		.taskOut_TVALID(_peArray_30_taskOut_TVALID),
		.taskOut_TDATA(_peArray_30_taskOut_TDATA),
		.taskIn_TREADY(_peArray_30_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_30_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_30_TDATA),
		.s_axi_control_ARREADY(fib_30_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_30_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_30_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_30_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_30_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_30_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_30_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_30_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_30_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_30_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_30_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_30_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_30_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_30_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_30_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_30_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_30_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_30_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_30_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_30_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_30_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_30_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_30_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_30_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_30_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_30_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_30_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_30_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_30_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_30_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_30_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_30_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_30_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_30_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_30_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_30_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_30_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_30_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_30_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_30_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_30_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_30_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_30_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_30_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_30_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_30_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_30_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_30_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_30_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_30_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_30_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_30_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_30_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_30_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_30_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_30_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_30_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_30_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_30_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_30_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_30_m_axi_gmem_BUSER)
	);
	fib peArray_31(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_31_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_31_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_31_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_31_TREADY),
		.argOut_TVALID(_peArray_31_argOut_TVALID),
		.argOut_TDATA(_peArray_31_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_31_TREADY),
		.taskOut_TVALID(_peArray_31_taskOut_TVALID),
		.taskOut_TDATA(_peArray_31_taskOut_TDATA),
		.taskIn_TREADY(_peArray_31_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_31_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_31_TDATA),
		.s_axi_control_ARREADY(fib_31_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_31_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_31_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_31_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_31_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_31_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_31_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_31_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_31_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_31_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_31_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_31_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_31_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_31_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_31_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_31_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_31_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_31_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_31_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_31_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_31_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_31_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_31_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_31_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_31_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_31_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_31_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_31_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_31_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_31_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_31_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_31_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_31_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_31_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_31_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_31_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_31_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_31_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_31_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_31_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_31_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_31_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_31_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_31_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_31_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_31_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_31_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_31_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_31_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_31_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_31_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_31_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_31_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_31_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_31_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_31_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_31_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_31_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_31_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_31_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_31_m_axi_gmem_BUSER)
	);
	fib peArray_32(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_32_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_32_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_32_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_32_TREADY),
		.argOut_TVALID(_peArray_32_argOut_TVALID),
		.argOut_TDATA(_peArray_32_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_32_TREADY),
		.taskOut_TVALID(_peArray_32_taskOut_TVALID),
		.taskOut_TDATA(_peArray_32_taskOut_TDATA),
		.taskIn_TREADY(_peArray_32_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_32_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_32_TDATA),
		.s_axi_control_ARREADY(fib_32_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_32_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_32_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_32_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_32_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_32_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_32_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_32_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_32_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_32_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_32_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_32_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_32_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_32_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_32_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_32_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_32_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_32_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_32_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_32_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_32_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_32_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_32_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_32_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_32_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_32_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_32_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_32_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_32_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_32_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_32_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_32_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_32_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_32_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_32_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_32_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_32_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_32_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_32_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_32_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_32_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_32_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_32_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_32_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_32_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_32_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_32_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_32_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_32_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_32_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_32_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_32_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_32_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_32_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_32_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_32_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_32_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_32_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_32_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_32_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_32_m_axi_gmem_BUSER)
	);
	fib peArray_33(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_33_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_33_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_33_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_33_TREADY),
		.argOut_TVALID(_peArray_33_argOut_TVALID),
		.argOut_TDATA(_peArray_33_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_33_TREADY),
		.taskOut_TVALID(_peArray_33_taskOut_TVALID),
		.taskOut_TDATA(_peArray_33_taskOut_TDATA),
		.taskIn_TREADY(_peArray_33_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_33_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_33_TDATA),
		.s_axi_control_ARREADY(fib_33_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_33_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_33_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_33_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_33_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_33_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_33_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_33_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_33_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_33_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_33_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_33_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_33_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_33_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_33_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_33_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_33_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_33_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_33_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_33_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_33_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_33_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_33_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_33_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_33_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_33_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_33_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_33_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_33_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_33_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_33_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_33_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_33_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_33_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_33_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_33_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_33_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_33_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_33_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_33_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_33_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_33_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_33_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_33_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_33_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_33_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_33_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_33_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_33_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_33_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_33_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_33_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_33_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_33_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_33_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_33_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_33_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_33_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_33_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_33_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_33_m_axi_gmem_BUSER)
	);
	fib peArray_34(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_34_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_34_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_34_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_34_TREADY),
		.argOut_TVALID(_peArray_34_argOut_TVALID),
		.argOut_TDATA(_peArray_34_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_34_TREADY),
		.taskOut_TVALID(_peArray_34_taskOut_TVALID),
		.taskOut_TDATA(_peArray_34_taskOut_TDATA),
		.taskIn_TREADY(_peArray_34_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_34_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_34_TDATA),
		.s_axi_control_ARREADY(fib_34_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_34_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_34_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_34_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_34_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_34_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_34_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_34_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_34_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_34_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_34_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_34_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_34_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_34_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_34_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_34_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_34_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_34_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_34_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_34_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_34_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_34_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_34_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_34_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_34_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_34_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_34_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_34_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_34_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_34_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_34_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_34_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_34_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_34_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_34_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_34_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_34_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_34_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_34_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_34_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_34_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_34_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_34_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_34_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_34_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_34_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_34_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_34_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_34_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_34_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_34_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_34_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_34_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_34_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_34_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_34_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_34_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_34_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_34_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_34_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_34_m_axi_gmem_BUSER)
	);
	fib peArray_35(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_35_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_35_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_35_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_35_TREADY),
		.argOut_TVALID(_peArray_35_argOut_TVALID),
		.argOut_TDATA(_peArray_35_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_35_TREADY),
		.taskOut_TVALID(_peArray_35_taskOut_TVALID),
		.taskOut_TDATA(_peArray_35_taskOut_TDATA),
		.taskIn_TREADY(_peArray_35_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_35_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_35_TDATA),
		.s_axi_control_ARREADY(fib_35_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_35_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_35_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_35_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_35_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_35_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_35_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_35_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_35_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_35_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_35_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_35_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_35_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_35_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_35_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_35_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_35_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_35_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_35_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_35_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_35_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_35_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_35_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_35_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_35_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_35_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_35_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_35_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_35_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_35_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_35_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_35_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_35_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_35_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_35_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_35_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_35_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_35_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_35_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_35_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_35_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_35_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_35_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_35_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_35_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_35_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_35_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_35_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_35_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_35_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_35_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_35_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_35_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_35_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_35_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_35_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_35_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_35_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_35_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_35_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_35_m_axi_gmem_BUSER)
	);
	fib peArray_36(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_36_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_36_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_36_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_36_TREADY),
		.argOut_TVALID(_peArray_36_argOut_TVALID),
		.argOut_TDATA(_peArray_36_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_36_TREADY),
		.taskOut_TVALID(_peArray_36_taskOut_TVALID),
		.taskOut_TDATA(_peArray_36_taskOut_TDATA),
		.taskIn_TREADY(_peArray_36_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_36_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_36_TDATA),
		.s_axi_control_ARREADY(fib_36_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_36_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_36_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_36_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_36_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_36_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_36_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_36_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_36_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_36_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_36_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_36_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_36_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_36_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_36_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_36_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_36_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_36_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_36_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_36_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_36_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_36_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_36_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_36_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_36_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_36_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_36_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_36_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_36_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_36_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_36_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_36_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_36_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_36_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_36_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_36_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_36_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_36_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_36_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_36_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_36_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_36_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_36_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_36_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_36_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_36_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_36_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_36_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_36_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_36_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_36_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_36_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_36_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_36_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_36_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_36_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_36_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_36_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_36_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_36_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_36_m_axi_gmem_BUSER)
	);
	fib peArray_37(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_37_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_37_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_37_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_37_TREADY),
		.argOut_TVALID(_peArray_37_argOut_TVALID),
		.argOut_TDATA(_peArray_37_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_37_TREADY),
		.taskOut_TVALID(_peArray_37_taskOut_TVALID),
		.taskOut_TDATA(_peArray_37_taskOut_TDATA),
		.taskIn_TREADY(_peArray_37_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_37_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_37_TDATA),
		.s_axi_control_ARREADY(fib_37_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_37_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_37_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_37_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_37_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_37_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_37_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_37_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_37_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_37_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_37_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_37_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_37_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_37_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_37_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_37_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_37_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_37_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_37_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_37_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_37_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_37_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_37_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_37_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_37_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_37_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_37_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_37_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_37_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_37_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_37_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_37_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_37_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_37_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_37_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_37_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_37_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_37_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_37_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_37_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_37_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_37_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_37_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_37_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_37_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_37_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_37_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_37_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_37_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_37_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_37_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_37_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_37_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_37_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_37_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_37_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_37_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_37_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_37_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_37_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_37_m_axi_gmem_BUSER)
	);
	fib peArray_38(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_38_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_38_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_38_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_38_TREADY),
		.argOut_TVALID(_peArray_38_argOut_TVALID),
		.argOut_TDATA(_peArray_38_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_38_TREADY),
		.taskOut_TVALID(_peArray_38_taskOut_TVALID),
		.taskOut_TDATA(_peArray_38_taskOut_TDATA),
		.taskIn_TREADY(_peArray_38_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_38_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_38_TDATA),
		.s_axi_control_ARREADY(fib_38_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_38_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_38_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_38_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_38_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_38_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_38_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_38_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_38_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_38_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_38_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_38_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_38_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_38_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_38_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_38_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_38_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_38_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_38_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_38_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_38_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_38_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_38_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_38_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_38_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_38_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_38_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_38_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_38_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_38_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_38_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_38_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_38_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_38_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_38_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_38_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_38_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_38_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_38_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_38_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_38_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_38_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_38_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_38_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_38_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_38_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_38_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_38_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_38_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_38_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_38_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_38_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_38_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_38_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_38_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_38_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_38_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_38_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_38_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_38_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_38_m_axi_gmem_BUSER)
	);
	fib peArray_39(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_39_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_39_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_39_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_39_TREADY),
		.argOut_TVALID(_peArray_39_argOut_TVALID),
		.argOut_TDATA(_peArray_39_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_39_TREADY),
		.taskOut_TVALID(_peArray_39_taskOut_TVALID),
		.taskOut_TDATA(_peArray_39_taskOut_TDATA),
		.taskIn_TREADY(_peArray_39_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_39_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_39_TDATA),
		.s_axi_control_ARREADY(fib_39_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_39_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_39_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_39_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_39_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_39_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_39_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_39_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_39_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_39_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_39_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_39_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_39_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_39_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_39_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_39_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_39_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_39_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_39_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_39_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_39_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_39_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_39_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_39_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_39_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_39_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_39_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_39_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_39_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_39_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_39_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_39_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_39_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_39_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_39_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_39_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_39_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_39_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_39_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_39_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_39_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_39_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_39_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_39_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_39_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_39_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_39_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_39_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_39_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_39_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_39_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_39_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_39_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_39_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_39_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_39_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_39_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_39_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_39_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_39_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_39_m_axi_gmem_BUSER)
	);
	fib peArray_40(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_40_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_40_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_40_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_40_TREADY),
		.argOut_TVALID(_peArray_40_argOut_TVALID),
		.argOut_TDATA(_peArray_40_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_40_TREADY),
		.taskOut_TVALID(_peArray_40_taskOut_TVALID),
		.taskOut_TDATA(_peArray_40_taskOut_TDATA),
		.taskIn_TREADY(_peArray_40_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_40_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_40_TDATA),
		.s_axi_control_ARREADY(fib_40_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_40_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_40_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_40_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_40_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_40_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_40_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_40_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_40_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_40_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_40_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_40_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_40_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_40_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_40_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_40_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_40_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_40_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_40_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_40_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_40_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_40_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_40_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_40_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_40_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_40_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_40_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_40_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_40_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_40_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_40_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_40_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_40_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_40_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_40_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_40_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_40_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_40_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_40_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_40_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_40_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_40_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_40_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_40_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_40_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_40_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_40_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_40_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_40_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_40_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_40_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_40_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_40_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_40_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_40_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_40_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_40_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_40_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_40_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_40_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_40_m_axi_gmem_BUSER)
	);
	fib peArray_41(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_41_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_41_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_41_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_41_TREADY),
		.argOut_TVALID(_peArray_41_argOut_TVALID),
		.argOut_TDATA(_peArray_41_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_41_TREADY),
		.taskOut_TVALID(_peArray_41_taskOut_TVALID),
		.taskOut_TDATA(_peArray_41_taskOut_TDATA),
		.taskIn_TREADY(_peArray_41_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_41_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_41_TDATA),
		.s_axi_control_ARREADY(fib_41_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_41_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_41_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_41_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_41_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_41_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_41_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_41_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_41_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_41_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_41_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_41_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_41_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_41_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_41_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_41_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_41_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_41_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_41_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_41_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_41_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_41_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_41_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_41_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_41_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_41_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_41_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_41_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_41_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_41_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_41_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_41_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_41_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_41_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_41_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_41_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_41_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_41_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_41_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_41_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_41_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_41_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_41_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_41_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_41_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_41_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_41_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_41_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_41_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_41_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_41_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_41_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_41_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_41_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_41_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_41_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_41_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_41_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_41_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_41_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_41_m_axi_gmem_BUSER)
	);
	fib peArray_42(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_42_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_42_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_42_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_42_TREADY),
		.argOut_TVALID(_peArray_42_argOut_TVALID),
		.argOut_TDATA(_peArray_42_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_42_TREADY),
		.taskOut_TVALID(_peArray_42_taskOut_TVALID),
		.taskOut_TDATA(_peArray_42_taskOut_TDATA),
		.taskIn_TREADY(_peArray_42_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_42_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_42_TDATA),
		.s_axi_control_ARREADY(fib_42_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_42_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_42_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_42_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_42_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_42_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_42_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_42_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_42_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_42_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_42_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_42_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_42_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_42_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_42_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_42_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_42_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_42_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_42_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_42_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_42_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_42_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_42_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_42_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_42_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_42_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_42_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_42_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_42_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_42_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_42_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_42_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_42_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_42_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_42_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_42_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_42_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_42_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_42_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_42_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_42_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_42_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_42_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_42_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_42_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_42_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_42_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_42_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_42_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_42_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_42_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_42_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_42_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_42_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_42_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_42_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_42_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_42_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_42_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_42_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_42_m_axi_gmem_BUSER)
	);
	fib peArray_43(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_43_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_43_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_43_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_43_TREADY),
		.argOut_TVALID(_peArray_43_argOut_TVALID),
		.argOut_TDATA(_peArray_43_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_43_TREADY),
		.taskOut_TVALID(_peArray_43_taskOut_TVALID),
		.taskOut_TDATA(_peArray_43_taskOut_TDATA),
		.taskIn_TREADY(_peArray_43_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_43_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_43_TDATA),
		.s_axi_control_ARREADY(fib_43_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_43_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_43_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_43_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_43_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_43_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_43_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_43_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_43_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_43_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_43_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_43_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_43_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_43_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_43_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_43_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_43_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_43_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_43_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_43_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_43_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_43_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_43_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_43_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_43_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_43_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_43_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_43_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_43_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_43_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_43_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_43_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_43_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_43_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_43_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_43_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_43_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_43_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_43_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_43_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_43_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_43_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_43_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_43_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_43_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_43_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_43_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_43_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_43_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_43_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_43_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_43_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_43_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_43_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_43_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_43_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_43_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_43_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_43_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_43_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_43_m_axi_gmem_BUSER)
	);
	fib peArray_44(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_44_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_44_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_44_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_44_TREADY),
		.argOut_TVALID(_peArray_44_argOut_TVALID),
		.argOut_TDATA(_peArray_44_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_44_TREADY),
		.taskOut_TVALID(_peArray_44_taskOut_TVALID),
		.taskOut_TDATA(_peArray_44_taskOut_TDATA),
		.taskIn_TREADY(_peArray_44_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_44_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_44_TDATA),
		.s_axi_control_ARREADY(fib_44_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_44_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_44_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_44_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_44_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_44_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_44_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_44_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_44_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_44_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_44_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_44_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_44_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_44_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_44_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_44_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_44_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_44_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_44_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_44_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_44_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_44_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_44_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_44_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_44_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_44_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_44_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_44_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_44_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_44_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_44_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_44_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_44_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_44_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_44_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_44_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_44_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_44_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_44_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_44_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_44_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_44_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_44_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_44_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_44_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_44_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_44_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_44_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_44_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_44_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_44_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_44_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_44_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_44_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_44_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_44_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_44_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_44_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_44_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_44_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_44_m_axi_gmem_BUSER)
	);
	fib peArray_45(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_45_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_45_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_45_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_45_TREADY),
		.argOut_TVALID(_peArray_45_argOut_TVALID),
		.argOut_TDATA(_peArray_45_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_45_TREADY),
		.taskOut_TVALID(_peArray_45_taskOut_TVALID),
		.taskOut_TDATA(_peArray_45_taskOut_TDATA),
		.taskIn_TREADY(_peArray_45_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_45_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_45_TDATA),
		.s_axi_control_ARREADY(fib_45_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_45_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_45_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_45_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_45_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_45_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_45_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_45_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_45_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_45_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_45_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_45_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_45_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_45_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_45_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_45_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_45_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_45_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_45_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_45_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_45_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_45_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_45_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_45_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_45_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_45_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_45_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_45_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_45_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_45_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_45_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_45_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_45_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_45_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_45_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_45_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_45_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_45_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_45_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_45_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_45_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_45_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_45_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_45_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_45_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_45_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_45_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_45_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_45_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_45_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_45_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_45_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_45_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_45_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_45_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_45_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_45_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_45_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_45_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_45_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_45_m_axi_gmem_BUSER)
	);
	fib peArray_46(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_46_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_46_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_46_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_46_TREADY),
		.argOut_TVALID(_peArray_46_argOut_TVALID),
		.argOut_TDATA(_peArray_46_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_46_TREADY),
		.taskOut_TVALID(_peArray_46_taskOut_TVALID),
		.taskOut_TDATA(_peArray_46_taskOut_TDATA),
		.taskIn_TREADY(_peArray_46_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_46_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_46_TDATA),
		.s_axi_control_ARREADY(fib_46_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_46_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_46_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_46_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_46_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_46_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_46_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_46_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_46_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_46_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_46_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_46_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_46_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_46_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_46_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_46_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_46_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_46_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_46_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_46_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_46_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_46_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_46_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_46_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_46_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_46_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_46_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_46_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_46_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_46_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_46_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_46_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_46_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_46_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_46_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_46_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_46_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_46_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_46_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_46_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_46_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_46_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_46_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_46_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_46_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_46_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_46_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_46_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_46_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_46_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_46_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_46_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_46_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_46_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_46_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_46_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_46_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_46_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_46_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_46_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_46_m_axi_gmem_BUSER)
	);
	fib peArray_47(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_47_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_47_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_47_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_47_TREADY),
		.argOut_TVALID(_peArray_47_argOut_TVALID),
		.argOut_TDATA(_peArray_47_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_47_TREADY),
		.taskOut_TVALID(_peArray_47_taskOut_TVALID),
		.taskOut_TDATA(_peArray_47_taskOut_TDATA),
		.taskIn_TREADY(_peArray_47_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_47_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_47_TDATA),
		.s_axi_control_ARREADY(fib_47_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_47_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_47_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_47_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_47_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_47_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_47_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_47_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_47_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_47_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_47_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_47_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_47_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_47_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_47_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_47_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_47_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_47_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_47_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_47_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_47_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_47_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_47_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_47_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_47_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_47_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_47_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_47_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_47_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_47_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_47_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_47_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_47_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_47_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_47_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_47_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_47_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_47_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_47_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_47_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_47_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_47_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_47_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_47_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_47_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_47_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_47_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_47_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_47_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_47_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_47_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_47_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_47_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_47_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_47_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_47_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_47_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_47_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_47_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_47_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_47_m_axi_gmem_BUSER)
	);
	fib peArray_48(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_48_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_48_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_48_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_48_TREADY),
		.argOut_TVALID(_peArray_48_argOut_TVALID),
		.argOut_TDATA(_peArray_48_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_48_TREADY),
		.taskOut_TVALID(_peArray_48_taskOut_TVALID),
		.taskOut_TDATA(_peArray_48_taskOut_TDATA),
		.taskIn_TREADY(_peArray_48_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_48_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_48_TDATA),
		.s_axi_control_ARREADY(fib_48_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_48_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_48_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_48_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_48_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_48_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_48_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_48_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_48_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_48_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_48_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_48_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_48_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_48_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_48_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_48_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_48_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_48_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_48_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_48_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_48_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_48_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_48_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_48_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_48_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_48_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_48_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_48_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_48_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_48_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_48_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_48_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_48_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_48_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_48_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_48_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_48_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_48_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_48_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_48_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_48_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_48_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_48_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_48_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_48_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_48_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_48_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_48_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_48_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_48_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_48_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_48_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_48_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_48_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_48_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_48_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_48_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_48_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_48_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_48_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_48_m_axi_gmem_BUSER)
	);
	fib peArray_49(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_49_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_49_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_49_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_49_TREADY),
		.argOut_TVALID(_peArray_49_argOut_TVALID),
		.argOut_TDATA(_peArray_49_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_49_TREADY),
		.taskOut_TVALID(_peArray_49_taskOut_TVALID),
		.taskOut_TDATA(_peArray_49_taskOut_TDATA),
		.taskIn_TREADY(_peArray_49_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_49_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_49_TDATA),
		.s_axi_control_ARREADY(fib_49_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_49_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_49_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_49_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_49_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_49_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_49_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_49_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_49_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_49_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_49_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_49_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_49_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_49_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_49_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_49_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_49_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_49_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_49_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_49_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_49_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_49_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_49_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_49_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_49_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_49_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_49_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_49_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_49_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_49_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_49_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_49_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_49_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_49_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_49_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_49_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_49_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_49_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_49_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_49_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_49_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_49_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_49_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_49_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_49_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_49_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_49_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_49_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_49_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_49_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_49_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_49_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_49_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_49_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_49_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_49_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_49_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_49_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_49_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_49_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_49_m_axi_gmem_BUSER)
	);
	fib peArray_50(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_50_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_50_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_50_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_50_TREADY),
		.argOut_TVALID(_peArray_50_argOut_TVALID),
		.argOut_TDATA(_peArray_50_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_50_TREADY),
		.taskOut_TVALID(_peArray_50_taskOut_TVALID),
		.taskOut_TDATA(_peArray_50_taskOut_TDATA),
		.taskIn_TREADY(_peArray_50_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_50_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_50_TDATA),
		.s_axi_control_ARREADY(fib_50_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_50_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_50_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_50_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_50_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_50_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_50_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_50_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_50_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_50_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_50_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_50_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_50_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_50_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_50_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_50_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_50_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_50_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_50_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_50_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_50_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_50_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_50_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_50_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_50_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_50_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_50_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_50_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_50_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_50_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_50_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_50_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_50_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_50_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_50_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_50_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_50_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_50_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_50_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_50_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_50_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_50_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_50_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_50_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_50_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_50_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_50_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_50_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_50_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_50_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_50_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_50_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_50_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_50_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_50_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_50_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_50_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_50_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_50_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_50_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_50_m_axi_gmem_BUSER)
	);
	fib peArray_51(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_51_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_51_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_51_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_51_TREADY),
		.argOut_TVALID(_peArray_51_argOut_TVALID),
		.argOut_TDATA(_peArray_51_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_51_TREADY),
		.taskOut_TVALID(_peArray_51_taskOut_TVALID),
		.taskOut_TDATA(_peArray_51_taskOut_TDATA),
		.taskIn_TREADY(_peArray_51_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_51_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_51_TDATA),
		.s_axi_control_ARREADY(fib_51_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_51_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_51_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_51_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_51_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_51_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_51_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_51_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_51_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_51_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_51_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_51_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_51_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_51_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_51_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_51_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_51_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_51_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_51_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_51_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_51_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_51_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_51_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_51_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_51_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_51_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_51_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_51_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_51_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_51_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_51_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_51_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_51_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_51_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_51_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_51_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_51_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_51_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_51_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_51_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_51_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_51_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_51_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_51_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_51_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_51_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_51_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_51_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_51_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_51_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_51_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_51_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_51_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_51_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_51_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_51_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_51_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_51_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_51_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_51_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_51_m_axi_gmem_BUSER)
	);
	fib peArray_52(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_52_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_52_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_52_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_52_TREADY),
		.argOut_TVALID(_peArray_52_argOut_TVALID),
		.argOut_TDATA(_peArray_52_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_52_TREADY),
		.taskOut_TVALID(_peArray_52_taskOut_TVALID),
		.taskOut_TDATA(_peArray_52_taskOut_TDATA),
		.taskIn_TREADY(_peArray_52_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_52_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_52_TDATA),
		.s_axi_control_ARREADY(fib_52_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_52_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_52_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_52_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_52_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_52_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_52_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_52_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_52_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_52_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_52_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_52_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_52_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_52_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_52_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_52_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_52_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_52_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_52_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_52_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_52_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_52_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_52_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_52_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_52_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_52_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_52_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_52_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_52_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_52_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_52_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_52_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_52_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_52_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_52_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_52_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_52_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_52_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_52_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_52_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_52_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_52_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_52_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_52_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_52_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_52_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_52_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_52_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_52_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_52_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_52_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_52_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_52_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_52_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_52_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_52_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_52_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_52_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_52_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_52_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_52_m_axi_gmem_BUSER)
	);
	fib peArray_53(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_53_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_53_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_53_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_53_TREADY),
		.argOut_TVALID(_peArray_53_argOut_TVALID),
		.argOut_TDATA(_peArray_53_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_53_TREADY),
		.taskOut_TVALID(_peArray_53_taskOut_TVALID),
		.taskOut_TDATA(_peArray_53_taskOut_TDATA),
		.taskIn_TREADY(_peArray_53_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_53_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_53_TDATA),
		.s_axi_control_ARREADY(fib_53_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_53_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_53_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_53_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_53_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_53_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_53_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_53_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_53_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_53_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_53_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_53_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_53_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_53_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_53_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_53_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_53_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_53_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_53_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_53_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_53_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_53_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_53_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_53_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_53_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_53_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_53_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_53_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_53_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_53_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_53_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_53_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_53_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_53_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_53_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_53_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_53_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_53_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_53_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_53_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_53_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_53_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_53_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_53_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_53_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_53_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_53_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_53_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_53_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_53_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_53_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_53_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_53_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_53_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_53_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_53_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_53_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_53_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_53_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_53_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_53_m_axi_gmem_BUSER)
	);
	fib peArray_54(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_54_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_54_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_54_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_54_TREADY),
		.argOut_TVALID(_peArray_54_argOut_TVALID),
		.argOut_TDATA(_peArray_54_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_54_TREADY),
		.taskOut_TVALID(_peArray_54_taskOut_TVALID),
		.taskOut_TDATA(_peArray_54_taskOut_TDATA),
		.taskIn_TREADY(_peArray_54_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_54_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_54_TDATA),
		.s_axi_control_ARREADY(fib_54_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_54_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_54_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_54_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_54_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_54_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_54_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_54_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_54_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_54_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_54_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_54_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_54_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_54_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_54_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_54_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_54_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_54_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_54_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_54_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_54_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_54_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_54_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_54_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_54_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_54_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_54_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_54_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_54_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_54_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_54_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_54_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_54_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_54_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_54_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_54_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_54_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_54_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_54_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_54_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_54_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_54_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_54_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_54_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_54_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_54_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_54_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_54_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_54_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_54_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_54_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_54_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_54_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_54_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_54_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_54_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_54_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_54_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_54_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_54_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_54_m_axi_gmem_BUSER)
	);
	fib peArray_55(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_55_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_55_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_55_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_55_TREADY),
		.argOut_TVALID(_peArray_55_argOut_TVALID),
		.argOut_TDATA(_peArray_55_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_55_TREADY),
		.taskOut_TVALID(_peArray_55_taskOut_TVALID),
		.taskOut_TDATA(_peArray_55_taskOut_TDATA),
		.taskIn_TREADY(_peArray_55_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_55_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_55_TDATA),
		.s_axi_control_ARREADY(fib_55_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_55_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_55_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_55_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_55_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_55_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_55_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_55_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_55_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_55_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_55_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_55_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_55_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_55_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_55_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_55_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_55_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_55_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_55_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_55_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_55_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_55_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_55_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_55_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_55_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_55_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_55_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_55_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_55_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_55_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_55_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_55_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_55_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_55_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_55_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_55_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_55_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_55_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_55_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_55_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_55_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_55_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_55_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_55_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_55_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_55_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_55_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_55_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_55_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_55_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_55_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_55_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_55_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_55_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_55_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_55_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_55_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_55_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_55_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_55_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_55_m_axi_gmem_BUSER)
	);
	fib peArray_56(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_56_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_56_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_56_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_56_TREADY),
		.argOut_TVALID(_peArray_56_argOut_TVALID),
		.argOut_TDATA(_peArray_56_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_56_TREADY),
		.taskOut_TVALID(_peArray_56_taskOut_TVALID),
		.taskOut_TDATA(_peArray_56_taskOut_TDATA),
		.taskIn_TREADY(_peArray_56_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_56_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_56_TDATA),
		.s_axi_control_ARREADY(fib_56_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_56_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_56_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_56_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_56_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_56_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_56_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_56_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_56_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_56_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_56_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_56_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_56_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_56_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_56_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_56_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_56_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_56_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_56_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_56_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_56_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_56_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_56_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_56_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_56_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_56_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_56_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_56_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_56_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_56_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_56_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_56_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_56_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_56_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_56_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_56_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_56_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_56_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_56_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_56_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_56_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_56_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_56_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_56_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_56_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_56_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_56_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_56_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_56_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_56_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_56_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_56_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_56_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_56_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_56_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_56_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_56_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_56_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_56_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_56_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_56_m_axi_gmem_BUSER)
	);
	fib peArray_57(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_57_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_57_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_57_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_57_TREADY),
		.argOut_TVALID(_peArray_57_argOut_TVALID),
		.argOut_TDATA(_peArray_57_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_57_TREADY),
		.taskOut_TVALID(_peArray_57_taskOut_TVALID),
		.taskOut_TDATA(_peArray_57_taskOut_TDATA),
		.taskIn_TREADY(_peArray_57_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_57_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_57_TDATA),
		.s_axi_control_ARREADY(fib_57_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_57_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_57_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_57_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_57_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_57_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_57_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_57_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_57_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_57_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_57_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_57_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_57_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_57_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_57_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_57_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_57_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_57_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_57_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_57_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_57_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_57_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_57_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_57_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_57_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_57_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_57_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_57_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_57_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_57_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_57_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_57_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_57_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_57_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_57_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_57_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_57_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_57_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_57_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_57_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_57_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_57_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_57_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_57_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_57_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_57_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_57_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_57_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_57_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_57_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_57_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_57_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_57_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_57_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_57_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_57_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_57_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_57_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_57_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_57_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_57_m_axi_gmem_BUSER)
	);
	fib peArray_58(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_58_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_58_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_58_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_58_TREADY),
		.argOut_TVALID(_peArray_58_argOut_TVALID),
		.argOut_TDATA(_peArray_58_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_58_TREADY),
		.taskOut_TVALID(_peArray_58_taskOut_TVALID),
		.taskOut_TDATA(_peArray_58_taskOut_TDATA),
		.taskIn_TREADY(_peArray_58_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_58_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_58_TDATA),
		.s_axi_control_ARREADY(fib_58_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_58_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_58_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_58_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_58_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_58_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_58_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_58_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_58_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_58_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_58_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_58_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_58_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_58_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_58_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_58_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_58_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_58_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_58_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_58_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_58_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_58_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_58_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_58_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_58_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_58_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_58_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_58_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_58_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_58_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_58_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_58_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_58_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_58_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_58_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_58_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_58_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_58_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_58_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_58_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_58_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_58_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_58_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_58_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_58_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_58_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_58_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_58_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_58_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_58_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_58_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_58_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_58_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_58_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_58_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_58_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_58_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_58_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_58_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_58_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_58_m_axi_gmem_BUSER)
	);
	fib peArray_59(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_59_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_59_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_59_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_59_TREADY),
		.argOut_TVALID(_peArray_59_argOut_TVALID),
		.argOut_TDATA(_peArray_59_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_59_TREADY),
		.taskOut_TVALID(_peArray_59_taskOut_TVALID),
		.taskOut_TDATA(_peArray_59_taskOut_TDATA),
		.taskIn_TREADY(_peArray_59_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_59_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_59_TDATA),
		.s_axi_control_ARREADY(fib_59_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_59_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_59_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_59_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_59_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_59_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_59_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_59_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_59_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_59_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_59_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_59_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_59_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_59_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_59_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_59_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_59_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_59_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_59_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_59_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_59_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_59_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_59_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_59_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_59_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_59_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_59_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_59_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_59_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_59_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_59_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_59_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_59_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_59_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_59_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_59_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_59_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_59_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_59_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_59_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_59_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_59_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_59_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_59_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_59_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_59_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_59_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_59_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_59_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_59_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_59_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_59_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_59_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_59_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_59_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_59_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_59_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_59_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_59_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_59_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_59_m_axi_gmem_BUSER)
	);
	fib peArray_60(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_60_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_60_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_60_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_60_TREADY),
		.argOut_TVALID(_peArray_60_argOut_TVALID),
		.argOut_TDATA(_peArray_60_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_60_TREADY),
		.taskOut_TVALID(_peArray_60_taskOut_TVALID),
		.taskOut_TDATA(_peArray_60_taskOut_TDATA),
		.taskIn_TREADY(_peArray_60_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_60_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_60_TDATA),
		.s_axi_control_ARREADY(fib_60_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_60_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_60_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_60_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_60_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_60_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_60_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_60_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_60_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_60_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_60_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_60_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_60_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_60_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_60_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_60_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_60_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_60_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_60_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_60_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_60_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_60_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_60_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_60_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_60_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_60_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_60_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_60_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_60_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_60_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_60_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_60_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_60_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_60_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_60_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_60_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_60_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_60_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_60_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_60_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_60_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_60_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_60_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_60_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_60_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_60_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_60_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_60_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_60_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_60_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_60_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_60_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_60_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_60_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_60_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_60_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_60_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_60_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_60_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_60_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_60_m_axi_gmem_BUSER)
	);
	fib peArray_61(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_61_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_61_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_61_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_61_TREADY),
		.argOut_TVALID(_peArray_61_argOut_TVALID),
		.argOut_TDATA(_peArray_61_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_61_TREADY),
		.taskOut_TVALID(_peArray_61_taskOut_TVALID),
		.taskOut_TDATA(_peArray_61_taskOut_TDATA),
		.taskIn_TREADY(_peArray_61_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_61_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_61_TDATA),
		.s_axi_control_ARREADY(fib_61_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_61_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_61_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_61_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_61_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_61_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_61_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_61_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_61_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_61_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_61_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_61_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_61_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_61_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_61_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_61_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_61_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_61_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_61_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_61_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_61_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_61_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_61_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_61_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_61_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_61_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_61_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_61_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_61_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_61_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_61_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_61_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_61_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_61_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_61_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_61_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_61_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_61_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_61_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_61_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_61_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_61_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_61_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_61_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_61_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_61_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_61_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_61_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_61_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_61_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_61_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_61_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_61_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_61_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_61_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_61_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_61_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_61_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_61_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_61_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_61_m_axi_gmem_BUSER)
	);
	fib peArray_62(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_62_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_62_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_62_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_62_TREADY),
		.argOut_TVALID(_peArray_62_argOut_TVALID),
		.argOut_TDATA(_peArray_62_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_62_TREADY),
		.taskOut_TVALID(_peArray_62_taskOut_TVALID),
		.taskOut_TDATA(_peArray_62_taskOut_TDATA),
		.taskIn_TREADY(_peArray_62_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_62_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_62_TDATA),
		.s_axi_control_ARREADY(fib_62_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_62_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_62_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_62_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_62_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_62_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_62_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_62_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_62_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_62_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_62_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_62_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_62_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_62_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_62_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_62_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_62_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_62_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_62_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_62_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_62_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_62_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_62_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_62_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_62_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_62_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_62_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_62_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_62_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_62_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_62_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_62_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_62_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_62_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_62_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_62_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_62_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_62_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_62_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_62_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_62_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_62_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_62_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_62_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_62_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_62_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_62_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_62_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_62_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_62_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_62_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_62_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_62_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_62_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_62_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_62_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_62_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_62_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_62_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_62_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_62_m_axi_gmem_BUSER)
	);
	fib peArray_63(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_63_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_63_TVALID),
		.closureIn_TDATA(_Allocator_io_export_closureOut_63_TDATA),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_63_TREADY),
		.argOut_TVALID(_peArray_63_argOut_TVALID),
		.argOut_TDATA(_peArray_63_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_63_TREADY),
		.taskOut_TVALID(_peArray_63_taskOut_TVALID),
		.taskOut_TDATA(_peArray_63_taskOut_TDATA),
		.taskIn_TREADY(_peArray_63_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_63_TVALID),
		.taskIn_TDATA(_Scheduler_io_export_taskOut_63_TDATA),
		.s_axi_control_ARREADY(fib_63_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(fib_63_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(fib_63_s_axi_control_ARADDR),
		.s_axi_control_RREADY(fib_63_s_axi_control_RREADY),
		.s_axi_control_RVALID(fib_63_s_axi_control_RVALID),
		.s_axi_control_RDATA(fib_63_s_axi_control_RDATA),
		.s_axi_control_RRESP(fib_63_s_axi_control_RRESP),
		.s_axi_control_AWREADY(fib_63_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(fib_63_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(fib_63_s_axi_control_AWADDR),
		.s_axi_control_WREADY(fib_63_s_axi_control_WREADY),
		.s_axi_control_WVALID(fib_63_s_axi_control_WVALID),
		.s_axi_control_WDATA(fib_63_s_axi_control_WDATA),
		.s_axi_control_WSTRB(fib_63_s_axi_control_WSTRB),
		.s_axi_control_BREADY(fib_63_s_axi_control_BREADY),
		.s_axi_control_BVALID(fib_63_s_axi_control_BVALID),
		.s_axi_control_BRESP(fib_63_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(fib_63_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(fib_63_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(fib_63_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(fib_63_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(fib_63_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(fib_63_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(fib_63_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(fib_63_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(fib_63_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(fib_63_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(fib_63_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(fib_63_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(fib_63_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(fib_63_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(fib_63_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(fib_63_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(fib_63_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(fib_63_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(fib_63_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(fib_63_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(fib_63_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(fib_63_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(fib_63_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(fib_63_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(fib_63_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(fib_63_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(fib_63_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(fib_63_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(fib_63_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(fib_63_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(fib_63_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(fib_63_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(fib_63_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(fib_63_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(fib_63_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(fib_63_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(fib_63_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(fib_63_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(fib_63_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(fib_63_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(fib_63_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(fib_63_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(fib_63_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(fib_63_m_axi_gmem_BUSER)
	);
	Scheduler Scheduler(
		.clock(clock),
		.reset(reset),
		.io_export_taskOut_0_TREADY(_peArray_0_taskIn_TREADY),
		.io_export_taskOut_0_TVALID(_Scheduler_io_export_taskOut_0_TVALID),
		.io_export_taskOut_0_TDATA(_Scheduler_io_export_taskOut_0_TDATA),
		.io_export_taskOut_1_TREADY(_peArray_1_taskIn_TREADY),
		.io_export_taskOut_1_TVALID(_Scheduler_io_export_taskOut_1_TVALID),
		.io_export_taskOut_1_TDATA(_Scheduler_io_export_taskOut_1_TDATA),
		.io_export_taskOut_2_TREADY(_peArray_2_taskIn_TREADY),
		.io_export_taskOut_2_TVALID(_Scheduler_io_export_taskOut_2_TVALID),
		.io_export_taskOut_2_TDATA(_Scheduler_io_export_taskOut_2_TDATA),
		.io_export_taskOut_3_TREADY(_peArray_3_taskIn_TREADY),
		.io_export_taskOut_3_TVALID(_Scheduler_io_export_taskOut_3_TVALID),
		.io_export_taskOut_3_TDATA(_Scheduler_io_export_taskOut_3_TDATA),
		.io_export_taskOut_4_TREADY(_peArray_4_taskIn_TREADY),
		.io_export_taskOut_4_TVALID(_Scheduler_io_export_taskOut_4_TVALID),
		.io_export_taskOut_4_TDATA(_Scheduler_io_export_taskOut_4_TDATA),
		.io_export_taskOut_5_TREADY(_peArray_5_taskIn_TREADY),
		.io_export_taskOut_5_TVALID(_Scheduler_io_export_taskOut_5_TVALID),
		.io_export_taskOut_5_TDATA(_Scheduler_io_export_taskOut_5_TDATA),
		.io_export_taskOut_6_TREADY(_peArray_6_taskIn_TREADY),
		.io_export_taskOut_6_TVALID(_Scheduler_io_export_taskOut_6_TVALID),
		.io_export_taskOut_6_TDATA(_Scheduler_io_export_taskOut_6_TDATA),
		.io_export_taskOut_7_TREADY(_peArray_7_taskIn_TREADY),
		.io_export_taskOut_7_TVALID(_Scheduler_io_export_taskOut_7_TVALID),
		.io_export_taskOut_7_TDATA(_Scheduler_io_export_taskOut_7_TDATA),
		.io_export_taskOut_8_TREADY(_peArray_8_taskIn_TREADY),
		.io_export_taskOut_8_TVALID(_Scheduler_io_export_taskOut_8_TVALID),
		.io_export_taskOut_8_TDATA(_Scheduler_io_export_taskOut_8_TDATA),
		.io_export_taskOut_9_TREADY(_peArray_9_taskIn_TREADY),
		.io_export_taskOut_9_TVALID(_Scheduler_io_export_taskOut_9_TVALID),
		.io_export_taskOut_9_TDATA(_Scheduler_io_export_taskOut_9_TDATA),
		.io_export_taskOut_10_TREADY(_peArray_10_taskIn_TREADY),
		.io_export_taskOut_10_TVALID(_Scheduler_io_export_taskOut_10_TVALID),
		.io_export_taskOut_10_TDATA(_Scheduler_io_export_taskOut_10_TDATA),
		.io_export_taskOut_11_TREADY(_peArray_11_taskIn_TREADY),
		.io_export_taskOut_11_TVALID(_Scheduler_io_export_taskOut_11_TVALID),
		.io_export_taskOut_11_TDATA(_Scheduler_io_export_taskOut_11_TDATA),
		.io_export_taskOut_12_TREADY(_peArray_12_taskIn_TREADY),
		.io_export_taskOut_12_TVALID(_Scheduler_io_export_taskOut_12_TVALID),
		.io_export_taskOut_12_TDATA(_Scheduler_io_export_taskOut_12_TDATA),
		.io_export_taskOut_13_TREADY(_peArray_13_taskIn_TREADY),
		.io_export_taskOut_13_TVALID(_Scheduler_io_export_taskOut_13_TVALID),
		.io_export_taskOut_13_TDATA(_Scheduler_io_export_taskOut_13_TDATA),
		.io_export_taskOut_14_TREADY(_peArray_14_taskIn_TREADY),
		.io_export_taskOut_14_TVALID(_Scheduler_io_export_taskOut_14_TVALID),
		.io_export_taskOut_14_TDATA(_Scheduler_io_export_taskOut_14_TDATA),
		.io_export_taskOut_15_TREADY(_peArray_15_taskIn_TREADY),
		.io_export_taskOut_15_TVALID(_Scheduler_io_export_taskOut_15_TVALID),
		.io_export_taskOut_15_TDATA(_Scheduler_io_export_taskOut_15_TDATA),
		.io_export_taskOut_16_TREADY(_peArray_16_taskIn_TREADY),
		.io_export_taskOut_16_TVALID(_Scheduler_io_export_taskOut_16_TVALID),
		.io_export_taskOut_16_TDATA(_Scheduler_io_export_taskOut_16_TDATA),
		.io_export_taskOut_17_TREADY(_peArray_17_taskIn_TREADY),
		.io_export_taskOut_17_TVALID(_Scheduler_io_export_taskOut_17_TVALID),
		.io_export_taskOut_17_TDATA(_Scheduler_io_export_taskOut_17_TDATA),
		.io_export_taskOut_18_TREADY(_peArray_18_taskIn_TREADY),
		.io_export_taskOut_18_TVALID(_Scheduler_io_export_taskOut_18_TVALID),
		.io_export_taskOut_18_TDATA(_Scheduler_io_export_taskOut_18_TDATA),
		.io_export_taskOut_19_TREADY(_peArray_19_taskIn_TREADY),
		.io_export_taskOut_19_TVALID(_Scheduler_io_export_taskOut_19_TVALID),
		.io_export_taskOut_19_TDATA(_Scheduler_io_export_taskOut_19_TDATA),
		.io_export_taskOut_20_TREADY(_peArray_20_taskIn_TREADY),
		.io_export_taskOut_20_TVALID(_Scheduler_io_export_taskOut_20_TVALID),
		.io_export_taskOut_20_TDATA(_Scheduler_io_export_taskOut_20_TDATA),
		.io_export_taskOut_21_TREADY(_peArray_21_taskIn_TREADY),
		.io_export_taskOut_21_TVALID(_Scheduler_io_export_taskOut_21_TVALID),
		.io_export_taskOut_21_TDATA(_Scheduler_io_export_taskOut_21_TDATA),
		.io_export_taskOut_22_TREADY(_peArray_22_taskIn_TREADY),
		.io_export_taskOut_22_TVALID(_Scheduler_io_export_taskOut_22_TVALID),
		.io_export_taskOut_22_TDATA(_Scheduler_io_export_taskOut_22_TDATA),
		.io_export_taskOut_23_TREADY(_peArray_23_taskIn_TREADY),
		.io_export_taskOut_23_TVALID(_Scheduler_io_export_taskOut_23_TVALID),
		.io_export_taskOut_23_TDATA(_Scheduler_io_export_taskOut_23_TDATA),
		.io_export_taskOut_24_TREADY(_peArray_24_taskIn_TREADY),
		.io_export_taskOut_24_TVALID(_Scheduler_io_export_taskOut_24_TVALID),
		.io_export_taskOut_24_TDATA(_Scheduler_io_export_taskOut_24_TDATA),
		.io_export_taskOut_25_TREADY(_peArray_25_taskIn_TREADY),
		.io_export_taskOut_25_TVALID(_Scheduler_io_export_taskOut_25_TVALID),
		.io_export_taskOut_25_TDATA(_Scheduler_io_export_taskOut_25_TDATA),
		.io_export_taskOut_26_TREADY(_peArray_26_taskIn_TREADY),
		.io_export_taskOut_26_TVALID(_Scheduler_io_export_taskOut_26_TVALID),
		.io_export_taskOut_26_TDATA(_Scheduler_io_export_taskOut_26_TDATA),
		.io_export_taskOut_27_TREADY(_peArray_27_taskIn_TREADY),
		.io_export_taskOut_27_TVALID(_Scheduler_io_export_taskOut_27_TVALID),
		.io_export_taskOut_27_TDATA(_Scheduler_io_export_taskOut_27_TDATA),
		.io_export_taskOut_28_TREADY(_peArray_28_taskIn_TREADY),
		.io_export_taskOut_28_TVALID(_Scheduler_io_export_taskOut_28_TVALID),
		.io_export_taskOut_28_TDATA(_Scheduler_io_export_taskOut_28_TDATA),
		.io_export_taskOut_29_TREADY(_peArray_29_taskIn_TREADY),
		.io_export_taskOut_29_TVALID(_Scheduler_io_export_taskOut_29_TVALID),
		.io_export_taskOut_29_TDATA(_Scheduler_io_export_taskOut_29_TDATA),
		.io_export_taskOut_30_TREADY(_peArray_30_taskIn_TREADY),
		.io_export_taskOut_30_TVALID(_Scheduler_io_export_taskOut_30_TVALID),
		.io_export_taskOut_30_TDATA(_Scheduler_io_export_taskOut_30_TDATA),
		.io_export_taskOut_31_TREADY(_peArray_31_taskIn_TREADY),
		.io_export_taskOut_31_TVALID(_Scheduler_io_export_taskOut_31_TVALID),
		.io_export_taskOut_31_TDATA(_Scheduler_io_export_taskOut_31_TDATA),
		.io_export_taskOut_32_TREADY(_peArray_32_taskIn_TREADY),
		.io_export_taskOut_32_TVALID(_Scheduler_io_export_taskOut_32_TVALID),
		.io_export_taskOut_32_TDATA(_Scheduler_io_export_taskOut_32_TDATA),
		.io_export_taskOut_33_TREADY(_peArray_33_taskIn_TREADY),
		.io_export_taskOut_33_TVALID(_Scheduler_io_export_taskOut_33_TVALID),
		.io_export_taskOut_33_TDATA(_Scheduler_io_export_taskOut_33_TDATA),
		.io_export_taskOut_34_TREADY(_peArray_34_taskIn_TREADY),
		.io_export_taskOut_34_TVALID(_Scheduler_io_export_taskOut_34_TVALID),
		.io_export_taskOut_34_TDATA(_Scheduler_io_export_taskOut_34_TDATA),
		.io_export_taskOut_35_TREADY(_peArray_35_taskIn_TREADY),
		.io_export_taskOut_35_TVALID(_Scheduler_io_export_taskOut_35_TVALID),
		.io_export_taskOut_35_TDATA(_Scheduler_io_export_taskOut_35_TDATA),
		.io_export_taskOut_36_TREADY(_peArray_36_taskIn_TREADY),
		.io_export_taskOut_36_TVALID(_Scheduler_io_export_taskOut_36_TVALID),
		.io_export_taskOut_36_TDATA(_Scheduler_io_export_taskOut_36_TDATA),
		.io_export_taskOut_37_TREADY(_peArray_37_taskIn_TREADY),
		.io_export_taskOut_37_TVALID(_Scheduler_io_export_taskOut_37_TVALID),
		.io_export_taskOut_37_TDATA(_Scheduler_io_export_taskOut_37_TDATA),
		.io_export_taskOut_38_TREADY(_peArray_38_taskIn_TREADY),
		.io_export_taskOut_38_TVALID(_Scheduler_io_export_taskOut_38_TVALID),
		.io_export_taskOut_38_TDATA(_Scheduler_io_export_taskOut_38_TDATA),
		.io_export_taskOut_39_TREADY(_peArray_39_taskIn_TREADY),
		.io_export_taskOut_39_TVALID(_Scheduler_io_export_taskOut_39_TVALID),
		.io_export_taskOut_39_TDATA(_Scheduler_io_export_taskOut_39_TDATA),
		.io_export_taskOut_40_TREADY(_peArray_40_taskIn_TREADY),
		.io_export_taskOut_40_TVALID(_Scheduler_io_export_taskOut_40_TVALID),
		.io_export_taskOut_40_TDATA(_Scheduler_io_export_taskOut_40_TDATA),
		.io_export_taskOut_41_TREADY(_peArray_41_taskIn_TREADY),
		.io_export_taskOut_41_TVALID(_Scheduler_io_export_taskOut_41_TVALID),
		.io_export_taskOut_41_TDATA(_Scheduler_io_export_taskOut_41_TDATA),
		.io_export_taskOut_42_TREADY(_peArray_42_taskIn_TREADY),
		.io_export_taskOut_42_TVALID(_Scheduler_io_export_taskOut_42_TVALID),
		.io_export_taskOut_42_TDATA(_Scheduler_io_export_taskOut_42_TDATA),
		.io_export_taskOut_43_TREADY(_peArray_43_taskIn_TREADY),
		.io_export_taskOut_43_TVALID(_Scheduler_io_export_taskOut_43_TVALID),
		.io_export_taskOut_43_TDATA(_Scheduler_io_export_taskOut_43_TDATA),
		.io_export_taskOut_44_TREADY(_peArray_44_taskIn_TREADY),
		.io_export_taskOut_44_TVALID(_Scheduler_io_export_taskOut_44_TVALID),
		.io_export_taskOut_44_TDATA(_Scheduler_io_export_taskOut_44_TDATA),
		.io_export_taskOut_45_TREADY(_peArray_45_taskIn_TREADY),
		.io_export_taskOut_45_TVALID(_Scheduler_io_export_taskOut_45_TVALID),
		.io_export_taskOut_45_TDATA(_Scheduler_io_export_taskOut_45_TDATA),
		.io_export_taskOut_46_TREADY(_peArray_46_taskIn_TREADY),
		.io_export_taskOut_46_TVALID(_Scheduler_io_export_taskOut_46_TVALID),
		.io_export_taskOut_46_TDATA(_Scheduler_io_export_taskOut_46_TDATA),
		.io_export_taskOut_47_TREADY(_peArray_47_taskIn_TREADY),
		.io_export_taskOut_47_TVALID(_Scheduler_io_export_taskOut_47_TVALID),
		.io_export_taskOut_47_TDATA(_Scheduler_io_export_taskOut_47_TDATA),
		.io_export_taskOut_48_TREADY(_peArray_48_taskIn_TREADY),
		.io_export_taskOut_48_TVALID(_Scheduler_io_export_taskOut_48_TVALID),
		.io_export_taskOut_48_TDATA(_Scheduler_io_export_taskOut_48_TDATA),
		.io_export_taskOut_49_TREADY(_peArray_49_taskIn_TREADY),
		.io_export_taskOut_49_TVALID(_Scheduler_io_export_taskOut_49_TVALID),
		.io_export_taskOut_49_TDATA(_Scheduler_io_export_taskOut_49_TDATA),
		.io_export_taskOut_50_TREADY(_peArray_50_taskIn_TREADY),
		.io_export_taskOut_50_TVALID(_Scheduler_io_export_taskOut_50_TVALID),
		.io_export_taskOut_50_TDATA(_Scheduler_io_export_taskOut_50_TDATA),
		.io_export_taskOut_51_TREADY(_peArray_51_taskIn_TREADY),
		.io_export_taskOut_51_TVALID(_Scheduler_io_export_taskOut_51_TVALID),
		.io_export_taskOut_51_TDATA(_Scheduler_io_export_taskOut_51_TDATA),
		.io_export_taskOut_52_TREADY(_peArray_52_taskIn_TREADY),
		.io_export_taskOut_52_TVALID(_Scheduler_io_export_taskOut_52_TVALID),
		.io_export_taskOut_52_TDATA(_Scheduler_io_export_taskOut_52_TDATA),
		.io_export_taskOut_53_TREADY(_peArray_53_taskIn_TREADY),
		.io_export_taskOut_53_TVALID(_Scheduler_io_export_taskOut_53_TVALID),
		.io_export_taskOut_53_TDATA(_Scheduler_io_export_taskOut_53_TDATA),
		.io_export_taskOut_54_TREADY(_peArray_54_taskIn_TREADY),
		.io_export_taskOut_54_TVALID(_Scheduler_io_export_taskOut_54_TVALID),
		.io_export_taskOut_54_TDATA(_Scheduler_io_export_taskOut_54_TDATA),
		.io_export_taskOut_55_TREADY(_peArray_55_taskIn_TREADY),
		.io_export_taskOut_55_TVALID(_Scheduler_io_export_taskOut_55_TVALID),
		.io_export_taskOut_55_TDATA(_Scheduler_io_export_taskOut_55_TDATA),
		.io_export_taskOut_56_TREADY(_peArray_56_taskIn_TREADY),
		.io_export_taskOut_56_TVALID(_Scheduler_io_export_taskOut_56_TVALID),
		.io_export_taskOut_56_TDATA(_Scheduler_io_export_taskOut_56_TDATA),
		.io_export_taskOut_57_TREADY(_peArray_57_taskIn_TREADY),
		.io_export_taskOut_57_TVALID(_Scheduler_io_export_taskOut_57_TVALID),
		.io_export_taskOut_57_TDATA(_Scheduler_io_export_taskOut_57_TDATA),
		.io_export_taskOut_58_TREADY(_peArray_58_taskIn_TREADY),
		.io_export_taskOut_58_TVALID(_Scheduler_io_export_taskOut_58_TVALID),
		.io_export_taskOut_58_TDATA(_Scheduler_io_export_taskOut_58_TDATA),
		.io_export_taskOut_59_TREADY(_peArray_59_taskIn_TREADY),
		.io_export_taskOut_59_TVALID(_Scheduler_io_export_taskOut_59_TVALID),
		.io_export_taskOut_59_TDATA(_Scheduler_io_export_taskOut_59_TDATA),
		.io_export_taskOut_60_TREADY(_peArray_60_taskIn_TREADY),
		.io_export_taskOut_60_TVALID(_Scheduler_io_export_taskOut_60_TVALID),
		.io_export_taskOut_60_TDATA(_Scheduler_io_export_taskOut_60_TDATA),
		.io_export_taskOut_61_TREADY(_peArray_61_taskIn_TREADY),
		.io_export_taskOut_61_TVALID(_Scheduler_io_export_taskOut_61_TVALID),
		.io_export_taskOut_61_TDATA(_Scheduler_io_export_taskOut_61_TDATA),
		.io_export_taskOut_62_TREADY(_peArray_62_taskIn_TREADY),
		.io_export_taskOut_62_TVALID(_Scheduler_io_export_taskOut_62_TVALID),
		.io_export_taskOut_62_TDATA(_Scheduler_io_export_taskOut_62_TDATA),
		.io_export_taskOut_63_TREADY(_peArray_63_taskIn_TREADY),
		.io_export_taskOut_63_TVALID(_Scheduler_io_export_taskOut_63_TVALID),
		.io_export_taskOut_63_TDATA(_Scheduler_io_export_taskOut_63_TDATA),
		.io_export_taskIn_0_TREADY(_Scheduler_io_export_taskIn_0_TREADY),
		.io_export_taskIn_0_TVALID(_peArray_0_taskOut_TVALID),
		.io_export_taskIn_0_TDATA(_peArray_0_taskOut_TDATA),
		.io_export_taskIn_1_TREADY(_Scheduler_io_export_taskIn_1_TREADY),
		.io_export_taskIn_1_TVALID(_peArray_1_taskOut_TVALID),
		.io_export_taskIn_1_TDATA(_peArray_1_taskOut_TDATA),
		.io_export_taskIn_2_TREADY(_Scheduler_io_export_taskIn_2_TREADY),
		.io_export_taskIn_2_TVALID(_peArray_2_taskOut_TVALID),
		.io_export_taskIn_2_TDATA(_peArray_2_taskOut_TDATA),
		.io_export_taskIn_3_TREADY(_Scheduler_io_export_taskIn_3_TREADY),
		.io_export_taskIn_3_TVALID(_peArray_3_taskOut_TVALID),
		.io_export_taskIn_3_TDATA(_peArray_3_taskOut_TDATA),
		.io_export_taskIn_4_TREADY(_Scheduler_io_export_taskIn_4_TREADY),
		.io_export_taskIn_4_TVALID(_peArray_4_taskOut_TVALID),
		.io_export_taskIn_4_TDATA(_peArray_4_taskOut_TDATA),
		.io_export_taskIn_5_TREADY(_Scheduler_io_export_taskIn_5_TREADY),
		.io_export_taskIn_5_TVALID(_peArray_5_taskOut_TVALID),
		.io_export_taskIn_5_TDATA(_peArray_5_taskOut_TDATA),
		.io_export_taskIn_6_TREADY(_Scheduler_io_export_taskIn_6_TREADY),
		.io_export_taskIn_6_TVALID(_peArray_6_taskOut_TVALID),
		.io_export_taskIn_6_TDATA(_peArray_6_taskOut_TDATA),
		.io_export_taskIn_7_TREADY(_Scheduler_io_export_taskIn_7_TREADY),
		.io_export_taskIn_7_TVALID(_peArray_7_taskOut_TVALID),
		.io_export_taskIn_7_TDATA(_peArray_7_taskOut_TDATA),
		.io_export_taskIn_8_TREADY(_Scheduler_io_export_taskIn_8_TREADY),
		.io_export_taskIn_8_TVALID(_peArray_8_taskOut_TVALID),
		.io_export_taskIn_8_TDATA(_peArray_8_taskOut_TDATA),
		.io_export_taskIn_9_TREADY(_Scheduler_io_export_taskIn_9_TREADY),
		.io_export_taskIn_9_TVALID(_peArray_9_taskOut_TVALID),
		.io_export_taskIn_9_TDATA(_peArray_9_taskOut_TDATA),
		.io_export_taskIn_10_TREADY(_Scheduler_io_export_taskIn_10_TREADY),
		.io_export_taskIn_10_TVALID(_peArray_10_taskOut_TVALID),
		.io_export_taskIn_10_TDATA(_peArray_10_taskOut_TDATA),
		.io_export_taskIn_11_TREADY(_Scheduler_io_export_taskIn_11_TREADY),
		.io_export_taskIn_11_TVALID(_peArray_11_taskOut_TVALID),
		.io_export_taskIn_11_TDATA(_peArray_11_taskOut_TDATA),
		.io_export_taskIn_12_TREADY(_Scheduler_io_export_taskIn_12_TREADY),
		.io_export_taskIn_12_TVALID(_peArray_12_taskOut_TVALID),
		.io_export_taskIn_12_TDATA(_peArray_12_taskOut_TDATA),
		.io_export_taskIn_13_TREADY(_Scheduler_io_export_taskIn_13_TREADY),
		.io_export_taskIn_13_TVALID(_peArray_13_taskOut_TVALID),
		.io_export_taskIn_13_TDATA(_peArray_13_taskOut_TDATA),
		.io_export_taskIn_14_TREADY(_Scheduler_io_export_taskIn_14_TREADY),
		.io_export_taskIn_14_TVALID(_peArray_14_taskOut_TVALID),
		.io_export_taskIn_14_TDATA(_peArray_14_taskOut_TDATA),
		.io_export_taskIn_15_TREADY(_Scheduler_io_export_taskIn_15_TREADY),
		.io_export_taskIn_15_TVALID(_peArray_15_taskOut_TVALID),
		.io_export_taskIn_15_TDATA(_peArray_15_taskOut_TDATA),
		.io_export_taskIn_16_TREADY(_Scheduler_io_export_taskIn_16_TREADY),
		.io_export_taskIn_16_TVALID(_peArray_16_taskOut_TVALID),
		.io_export_taskIn_16_TDATA(_peArray_16_taskOut_TDATA),
		.io_export_taskIn_17_TREADY(_Scheduler_io_export_taskIn_17_TREADY),
		.io_export_taskIn_17_TVALID(_peArray_17_taskOut_TVALID),
		.io_export_taskIn_17_TDATA(_peArray_17_taskOut_TDATA),
		.io_export_taskIn_18_TREADY(_Scheduler_io_export_taskIn_18_TREADY),
		.io_export_taskIn_18_TVALID(_peArray_18_taskOut_TVALID),
		.io_export_taskIn_18_TDATA(_peArray_18_taskOut_TDATA),
		.io_export_taskIn_19_TREADY(_Scheduler_io_export_taskIn_19_TREADY),
		.io_export_taskIn_19_TVALID(_peArray_19_taskOut_TVALID),
		.io_export_taskIn_19_TDATA(_peArray_19_taskOut_TDATA),
		.io_export_taskIn_20_TREADY(_Scheduler_io_export_taskIn_20_TREADY),
		.io_export_taskIn_20_TVALID(_peArray_20_taskOut_TVALID),
		.io_export_taskIn_20_TDATA(_peArray_20_taskOut_TDATA),
		.io_export_taskIn_21_TREADY(_Scheduler_io_export_taskIn_21_TREADY),
		.io_export_taskIn_21_TVALID(_peArray_21_taskOut_TVALID),
		.io_export_taskIn_21_TDATA(_peArray_21_taskOut_TDATA),
		.io_export_taskIn_22_TREADY(_Scheduler_io_export_taskIn_22_TREADY),
		.io_export_taskIn_22_TVALID(_peArray_22_taskOut_TVALID),
		.io_export_taskIn_22_TDATA(_peArray_22_taskOut_TDATA),
		.io_export_taskIn_23_TREADY(_Scheduler_io_export_taskIn_23_TREADY),
		.io_export_taskIn_23_TVALID(_peArray_23_taskOut_TVALID),
		.io_export_taskIn_23_TDATA(_peArray_23_taskOut_TDATA),
		.io_export_taskIn_24_TREADY(_Scheduler_io_export_taskIn_24_TREADY),
		.io_export_taskIn_24_TVALID(_peArray_24_taskOut_TVALID),
		.io_export_taskIn_24_TDATA(_peArray_24_taskOut_TDATA),
		.io_export_taskIn_25_TREADY(_Scheduler_io_export_taskIn_25_TREADY),
		.io_export_taskIn_25_TVALID(_peArray_25_taskOut_TVALID),
		.io_export_taskIn_25_TDATA(_peArray_25_taskOut_TDATA),
		.io_export_taskIn_26_TREADY(_Scheduler_io_export_taskIn_26_TREADY),
		.io_export_taskIn_26_TVALID(_peArray_26_taskOut_TVALID),
		.io_export_taskIn_26_TDATA(_peArray_26_taskOut_TDATA),
		.io_export_taskIn_27_TREADY(_Scheduler_io_export_taskIn_27_TREADY),
		.io_export_taskIn_27_TVALID(_peArray_27_taskOut_TVALID),
		.io_export_taskIn_27_TDATA(_peArray_27_taskOut_TDATA),
		.io_export_taskIn_28_TREADY(_Scheduler_io_export_taskIn_28_TREADY),
		.io_export_taskIn_28_TVALID(_peArray_28_taskOut_TVALID),
		.io_export_taskIn_28_TDATA(_peArray_28_taskOut_TDATA),
		.io_export_taskIn_29_TREADY(_Scheduler_io_export_taskIn_29_TREADY),
		.io_export_taskIn_29_TVALID(_peArray_29_taskOut_TVALID),
		.io_export_taskIn_29_TDATA(_peArray_29_taskOut_TDATA),
		.io_export_taskIn_30_TREADY(_Scheduler_io_export_taskIn_30_TREADY),
		.io_export_taskIn_30_TVALID(_peArray_30_taskOut_TVALID),
		.io_export_taskIn_30_TDATA(_peArray_30_taskOut_TDATA),
		.io_export_taskIn_31_TREADY(_Scheduler_io_export_taskIn_31_TREADY),
		.io_export_taskIn_31_TVALID(_peArray_31_taskOut_TVALID),
		.io_export_taskIn_31_TDATA(_peArray_31_taskOut_TDATA),
		.io_export_taskIn_32_TREADY(_Scheduler_io_export_taskIn_32_TREADY),
		.io_export_taskIn_32_TVALID(_peArray_32_taskOut_TVALID),
		.io_export_taskIn_32_TDATA(_peArray_32_taskOut_TDATA),
		.io_export_taskIn_33_TREADY(_Scheduler_io_export_taskIn_33_TREADY),
		.io_export_taskIn_33_TVALID(_peArray_33_taskOut_TVALID),
		.io_export_taskIn_33_TDATA(_peArray_33_taskOut_TDATA),
		.io_export_taskIn_34_TREADY(_Scheduler_io_export_taskIn_34_TREADY),
		.io_export_taskIn_34_TVALID(_peArray_34_taskOut_TVALID),
		.io_export_taskIn_34_TDATA(_peArray_34_taskOut_TDATA),
		.io_export_taskIn_35_TREADY(_Scheduler_io_export_taskIn_35_TREADY),
		.io_export_taskIn_35_TVALID(_peArray_35_taskOut_TVALID),
		.io_export_taskIn_35_TDATA(_peArray_35_taskOut_TDATA),
		.io_export_taskIn_36_TREADY(_Scheduler_io_export_taskIn_36_TREADY),
		.io_export_taskIn_36_TVALID(_peArray_36_taskOut_TVALID),
		.io_export_taskIn_36_TDATA(_peArray_36_taskOut_TDATA),
		.io_export_taskIn_37_TREADY(_Scheduler_io_export_taskIn_37_TREADY),
		.io_export_taskIn_37_TVALID(_peArray_37_taskOut_TVALID),
		.io_export_taskIn_37_TDATA(_peArray_37_taskOut_TDATA),
		.io_export_taskIn_38_TREADY(_Scheduler_io_export_taskIn_38_TREADY),
		.io_export_taskIn_38_TVALID(_peArray_38_taskOut_TVALID),
		.io_export_taskIn_38_TDATA(_peArray_38_taskOut_TDATA),
		.io_export_taskIn_39_TREADY(_Scheduler_io_export_taskIn_39_TREADY),
		.io_export_taskIn_39_TVALID(_peArray_39_taskOut_TVALID),
		.io_export_taskIn_39_TDATA(_peArray_39_taskOut_TDATA),
		.io_export_taskIn_40_TREADY(_Scheduler_io_export_taskIn_40_TREADY),
		.io_export_taskIn_40_TVALID(_peArray_40_taskOut_TVALID),
		.io_export_taskIn_40_TDATA(_peArray_40_taskOut_TDATA),
		.io_export_taskIn_41_TREADY(_Scheduler_io_export_taskIn_41_TREADY),
		.io_export_taskIn_41_TVALID(_peArray_41_taskOut_TVALID),
		.io_export_taskIn_41_TDATA(_peArray_41_taskOut_TDATA),
		.io_export_taskIn_42_TREADY(_Scheduler_io_export_taskIn_42_TREADY),
		.io_export_taskIn_42_TVALID(_peArray_42_taskOut_TVALID),
		.io_export_taskIn_42_TDATA(_peArray_42_taskOut_TDATA),
		.io_export_taskIn_43_TREADY(_Scheduler_io_export_taskIn_43_TREADY),
		.io_export_taskIn_43_TVALID(_peArray_43_taskOut_TVALID),
		.io_export_taskIn_43_TDATA(_peArray_43_taskOut_TDATA),
		.io_export_taskIn_44_TREADY(_Scheduler_io_export_taskIn_44_TREADY),
		.io_export_taskIn_44_TVALID(_peArray_44_taskOut_TVALID),
		.io_export_taskIn_44_TDATA(_peArray_44_taskOut_TDATA),
		.io_export_taskIn_45_TREADY(_Scheduler_io_export_taskIn_45_TREADY),
		.io_export_taskIn_45_TVALID(_peArray_45_taskOut_TVALID),
		.io_export_taskIn_45_TDATA(_peArray_45_taskOut_TDATA),
		.io_export_taskIn_46_TREADY(_Scheduler_io_export_taskIn_46_TREADY),
		.io_export_taskIn_46_TVALID(_peArray_46_taskOut_TVALID),
		.io_export_taskIn_46_TDATA(_peArray_46_taskOut_TDATA),
		.io_export_taskIn_47_TREADY(_Scheduler_io_export_taskIn_47_TREADY),
		.io_export_taskIn_47_TVALID(_peArray_47_taskOut_TVALID),
		.io_export_taskIn_47_TDATA(_peArray_47_taskOut_TDATA),
		.io_export_taskIn_48_TREADY(_Scheduler_io_export_taskIn_48_TREADY),
		.io_export_taskIn_48_TVALID(_peArray_48_taskOut_TVALID),
		.io_export_taskIn_48_TDATA(_peArray_48_taskOut_TDATA),
		.io_export_taskIn_49_TREADY(_Scheduler_io_export_taskIn_49_TREADY),
		.io_export_taskIn_49_TVALID(_peArray_49_taskOut_TVALID),
		.io_export_taskIn_49_TDATA(_peArray_49_taskOut_TDATA),
		.io_export_taskIn_50_TREADY(_Scheduler_io_export_taskIn_50_TREADY),
		.io_export_taskIn_50_TVALID(_peArray_50_taskOut_TVALID),
		.io_export_taskIn_50_TDATA(_peArray_50_taskOut_TDATA),
		.io_export_taskIn_51_TREADY(_Scheduler_io_export_taskIn_51_TREADY),
		.io_export_taskIn_51_TVALID(_peArray_51_taskOut_TVALID),
		.io_export_taskIn_51_TDATA(_peArray_51_taskOut_TDATA),
		.io_export_taskIn_52_TREADY(_Scheduler_io_export_taskIn_52_TREADY),
		.io_export_taskIn_52_TVALID(_peArray_52_taskOut_TVALID),
		.io_export_taskIn_52_TDATA(_peArray_52_taskOut_TDATA),
		.io_export_taskIn_53_TREADY(_Scheduler_io_export_taskIn_53_TREADY),
		.io_export_taskIn_53_TVALID(_peArray_53_taskOut_TVALID),
		.io_export_taskIn_53_TDATA(_peArray_53_taskOut_TDATA),
		.io_export_taskIn_54_TREADY(_Scheduler_io_export_taskIn_54_TREADY),
		.io_export_taskIn_54_TVALID(_peArray_54_taskOut_TVALID),
		.io_export_taskIn_54_TDATA(_peArray_54_taskOut_TDATA),
		.io_export_taskIn_55_TREADY(_Scheduler_io_export_taskIn_55_TREADY),
		.io_export_taskIn_55_TVALID(_peArray_55_taskOut_TVALID),
		.io_export_taskIn_55_TDATA(_peArray_55_taskOut_TDATA),
		.io_export_taskIn_56_TREADY(_Scheduler_io_export_taskIn_56_TREADY),
		.io_export_taskIn_56_TVALID(_peArray_56_taskOut_TVALID),
		.io_export_taskIn_56_TDATA(_peArray_56_taskOut_TDATA),
		.io_export_taskIn_57_TREADY(_Scheduler_io_export_taskIn_57_TREADY),
		.io_export_taskIn_57_TVALID(_peArray_57_taskOut_TVALID),
		.io_export_taskIn_57_TDATA(_peArray_57_taskOut_TDATA),
		.io_export_taskIn_58_TREADY(_Scheduler_io_export_taskIn_58_TREADY),
		.io_export_taskIn_58_TVALID(_peArray_58_taskOut_TVALID),
		.io_export_taskIn_58_TDATA(_peArray_58_taskOut_TDATA),
		.io_export_taskIn_59_TREADY(_Scheduler_io_export_taskIn_59_TREADY),
		.io_export_taskIn_59_TVALID(_peArray_59_taskOut_TVALID),
		.io_export_taskIn_59_TDATA(_peArray_59_taskOut_TDATA),
		.io_export_taskIn_60_TREADY(_Scheduler_io_export_taskIn_60_TREADY),
		.io_export_taskIn_60_TVALID(_peArray_60_taskOut_TVALID),
		.io_export_taskIn_60_TDATA(_peArray_60_taskOut_TDATA),
		.io_export_taskIn_61_TREADY(_Scheduler_io_export_taskIn_61_TREADY),
		.io_export_taskIn_61_TVALID(_peArray_61_taskOut_TVALID),
		.io_export_taskIn_61_TDATA(_peArray_61_taskOut_TDATA),
		.io_export_taskIn_62_TREADY(_Scheduler_io_export_taskIn_62_TREADY),
		.io_export_taskIn_62_TVALID(_peArray_62_taskOut_TVALID),
		.io_export_taskIn_62_TDATA(_peArray_62_taskOut_TDATA),
		.io_export_taskIn_63_TREADY(_Scheduler_io_export_taskIn_63_TREADY),
		.io_export_taskIn_63_TVALID(_peArray_63_taskOut_TVALID),
		.io_export_taskIn_63_TDATA(_peArray_63_taskOut_TDATA),
		.io_internal_vss_axi_full_0_ar_ready(fib_schedulerAXI_0_ARREADY),
		.io_internal_vss_axi_full_0_ar_valid(fib_schedulerAXI_0_ARVALID),
		.io_internal_vss_axi_full_0_ar_bits_id(fib_schedulerAXI_0_ARID),
		.io_internal_vss_axi_full_0_ar_bits_addr(fib_schedulerAXI_0_ARADDR),
		.io_internal_vss_axi_full_0_ar_bits_len(fib_schedulerAXI_0_ARLEN),
		.io_internal_vss_axi_full_0_ar_bits_size(fib_schedulerAXI_0_ARSIZE),
		.io_internal_vss_axi_full_0_ar_bits_burst(fib_schedulerAXI_0_ARBURST),
		.io_internal_vss_axi_full_0_ar_bits_lock(fib_schedulerAXI_0_ARLOCK),
		.io_internal_vss_axi_full_0_ar_bits_cache(fib_schedulerAXI_0_ARCACHE),
		.io_internal_vss_axi_full_0_ar_bits_prot(fib_schedulerAXI_0_ARPROT),
		.io_internal_vss_axi_full_0_ar_bits_qos(fib_schedulerAXI_0_ARQOS),
		.io_internal_vss_axi_full_0_ar_bits_region(fib_schedulerAXI_0_ARREGION),
		.io_internal_vss_axi_full_0_r_ready(fib_schedulerAXI_0_RREADY),
		.io_internal_vss_axi_full_0_r_valid(fib_schedulerAXI_0_RVALID),
		.io_internal_vss_axi_full_0_r_bits_id(fib_schedulerAXI_0_RID),
		.io_internal_vss_axi_full_0_r_bits_data(fib_schedulerAXI_0_RDATA),
		.io_internal_vss_axi_full_0_r_bits_resp(fib_schedulerAXI_0_RRESP),
		.io_internal_vss_axi_full_0_r_bits_last(fib_schedulerAXI_0_RLAST),
		.io_internal_vss_axi_full_0_aw_ready(fib_schedulerAXI_0_AWREADY),
		.io_internal_vss_axi_full_0_aw_valid(fib_schedulerAXI_0_AWVALID),
		.io_internal_vss_axi_full_0_aw_bits_id(fib_schedulerAXI_0_AWID),
		.io_internal_vss_axi_full_0_aw_bits_addr(fib_schedulerAXI_0_AWADDR),
		.io_internal_vss_axi_full_0_aw_bits_len(fib_schedulerAXI_0_AWLEN),
		.io_internal_vss_axi_full_0_aw_bits_size(fib_schedulerAXI_0_AWSIZE),
		.io_internal_vss_axi_full_0_aw_bits_burst(fib_schedulerAXI_0_AWBURST),
		.io_internal_vss_axi_full_0_aw_bits_lock(fib_schedulerAXI_0_AWLOCK),
		.io_internal_vss_axi_full_0_aw_bits_cache(fib_schedulerAXI_0_AWCACHE),
		.io_internal_vss_axi_full_0_aw_bits_prot(fib_schedulerAXI_0_AWPROT),
		.io_internal_vss_axi_full_0_aw_bits_qos(fib_schedulerAXI_0_AWQOS),
		.io_internal_vss_axi_full_0_aw_bits_region(fib_schedulerAXI_0_AWREGION),
		.io_internal_vss_axi_full_0_w_ready(fib_schedulerAXI_0_WREADY),
		.io_internal_vss_axi_full_0_w_valid(fib_schedulerAXI_0_WVALID),
		.io_internal_vss_axi_full_0_w_bits_data(fib_schedulerAXI_0_WDATA),
		.io_internal_vss_axi_full_0_w_bits_strb(fib_schedulerAXI_0_WSTRB),
		.io_internal_vss_axi_full_0_w_bits_last(fib_schedulerAXI_0_WLAST),
		.io_internal_vss_axi_full_0_b_ready(fib_schedulerAXI_0_BREADY),
		.io_internal_vss_axi_full_0_b_valid(fib_schedulerAXI_0_BVALID),
		.io_internal_vss_axi_full_0_b_bits_id(fib_schedulerAXI_0_BID),
		.io_internal_vss_axi_full_0_b_bits_resp(fib_schedulerAXI_0_BRESP),
		.io_internal_axi_mgmt_vss_0_ar_ready(_Scheduler_io_internal_axi_mgmt_vss_0_ar_ready),
		.io_internal_axi_mgmt_vss_0_ar_valid(_demux_m_axil_0_ar_valid),
		.io_internal_axi_mgmt_vss_0_ar_bits_addr(_demux_m_axil_0_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_ar_bits_prot(_demux_m_axil_0_ar_bits_prot),
		.io_internal_axi_mgmt_vss_0_r_ready(_demux_m_axil_0_r_ready),
		.io_internal_axi_mgmt_vss_0_r_valid(_Scheduler_io_internal_axi_mgmt_vss_0_r_valid),
		.io_internal_axi_mgmt_vss_0_r_bits_data(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_internal_axi_mgmt_vss_0_r_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_internal_axi_mgmt_vss_0_aw_ready(_Scheduler_io_internal_axi_mgmt_vss_0_aw_ready),
		.io_internal_axi_mgmt_vss_0_aw_valid(_demux_m_axil_0_aw_valid),
		.io_internal_axi_mgmt_vss_0_aw_bits_addr(_demux_m_axil_0_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_aw_bits_prot(_demux_m_axil_0_aw_bits_prot),
		.io_internal_axi_mgmt_vss_0_w_ready(_Scheduler_io_internal_axi_mgmt_vss_0_w_ready),
		.io_internal_axi_mgmt_vss_0_w_valid(_demux_m_axil_0_w_valid),
		.io_internal_axi_mgmt_vss_0_w_bits_data(_demux_m_axil_0_w_bits_data),
		.io_internal_axi_mgmt_vss_0_w_bits_strb(_demux_m_axil_0_w_bits_strb),
		.io_internal_axi_mgmt_vss_0_b_ready(_demux_m_axil_0_b_ready),
		.io_internal_axi_mgmt_vss_0_b_valid(_Scheduler_io_internal_axi_mgmt_vss_0_b_valid),
		.io_internal_axi_mgmt_vss_0_b_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.io_internal_axi_mgmt_vss_1_ar_ready(_Scheduler_io_internal_axi_mgmt_vss_1_ar_ready),
		.io_internal_axi_mgmt_vss_1_ar_valid(_demux_m_axil_1_ar_valid),
		.io_internal_axi_mgmt_vss_1_ar_bits_addr(_demux_m_axil_1_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_1_ar_bits_prot(_demux_m_axil_1_ar_bits_prot),
		.io_internal_axi_mgmt_vss_1_r_ready(_demux_m_axil_1_r_ready),
		.io_internal_axi_mgmt_vss_1_r_valid(_Scheduler_io_internal_axi_mgmt_vss_1_r_valid),
		.io_internal_axi_mgmt_vss_1_r_bits_data(_Scheduler_io_internal_axi_mgmt_vss_1_r_bits_data),
		.io_internal_axi_mgmt_vss_1_r_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_1_r_bits_resp),
		.io_internal_axi_mgmt_vss_1_aw_ready(_Scheduler_io_internal_axi_mgmt_vss_1_aw_ready),
		.io_internal_axi_mgmt_vss_1_aw_valid(_demux_m_axil_1_aw_valid),
		.io_internal_axi_mgmt_vss_1_aw_bits_addr(_demux_m_axil_1_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_1_aw_bits_prot(_demux_m_axil_1_aw_bits_prot),
		.io_internal_axi_mgmt_vss_1_w_ready(_Scheduler_io_internal_axi_mgmt_vss_1_w_ready),
		.io_internal_axi_mgmt_vss_1_w_valid(_demux_m_axil_1_w_valid),
		.io_internal_axi_mgmt_vss_1_w_bits_data(_demux_m_axil_1_w_bits_data),
		.io_internal_axi_mgmt_vss_1_w_bits_strb(_demux_m_axil_1_w_bits_strb),
		.io_internal_axi_mgmt_vss_1_b_ready(_demux_m_axil_1_b_ready),
		.io_internal_axi_mgmt_vss_1_b_valid(_Scheduler_io_internal_axi_mgmt_vss_1_b_valid),
		.io_internal_axi_mgmt_vss_1_b_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_1_b_bits_resp)
	);
	sum peArray_0_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_64_TREADY),
		.argOut_TVALID(_peArray_0_1_argOut_TVALID),
		.argOut_TDATA(_peArray_0_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_0_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_0_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_0_TDATA),
		.s_axi_control_ARREADY(sum_0_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_0_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_0_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_0_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_0_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_0_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_0_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_0_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_0_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_0_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_0_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_0_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_0_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_0_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_0_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_0_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_0_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_0_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_0_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_0_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_0_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_0_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_0_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_0_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_0_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_0_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_0_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_0_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_0_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_0_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_0_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_0_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_0_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_0_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_0_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_0_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_0_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_0_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_0_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_0_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_0_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_0_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_0_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_0_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_0_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_0_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_0_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_0_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_0_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_0_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_0_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_0_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_0_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_0_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_0_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_0_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_0_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_0_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_0_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_0_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_0_m_axi_gmem_BUSER)
	);
	sum peArray_1_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_65_TREADY),
		.argOut_TVALID(_peArray_1_1_argOut_TVALID),
		.argOut_TDATA(_peArray_1_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_1_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_1_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_1_TDATA),
		.s_axi_control_ARREADY(sum_1_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_1_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_1_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_1_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_1_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_1_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_1_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_1_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_1_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_1_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_1_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_1_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_1_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_1_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_1_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_1_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_1_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_1_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_1_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_1_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_1_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_1_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_1_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_1_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_1_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_1_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_1_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_1_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_1_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_1_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_1_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_1_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_1_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_1_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_1_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_1_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_1_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_1_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_1_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_1_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_1_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_1_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_1_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_1_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_1_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_1_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_1_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_1_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_1_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_1_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_1_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_1_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_1_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_1_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_1_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_1_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_1_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_1_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_1_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_1_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_1_m_axi_gmem_BUSER)
	);
	sum peArray_2_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_66_TREADY),
		.argOut_TVALID(_peArray_2_1_argOut_TVALID),
		.argOut_TDATA(_peArray_2_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_2_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_2_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_2_TDATA),
		.s_axi_control_ARREADY(sum_2_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_2_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_2_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_2_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_2_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_2_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_2_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_2_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_2_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_2_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_2_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_2_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_2_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_2_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_2_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_2_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_2_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_2_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_2_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_2_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_2_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_2_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_2_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_2_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_2_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_2_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_2_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_2_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_2_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_2_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_2_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_2_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_2_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_2_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_2_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_2_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_2_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_2_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_2_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_2_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_2_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_2_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_2_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_2_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_2_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_2_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_2_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_2_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_2_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_2_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_2_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_2_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_2_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_2_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_2_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_2_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_2_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_2_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_2_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_2_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_2_m_axi_gmem_BUSER)
	);
	sum peArray_3_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_67_TREADY),
		.argOut_TVALID(_peArray_3_1_argOut_TVALID),
		.argOut_TDATA(_peArray_3_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_3_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_3_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_3_TDATA),
		.s_axi_control_ARREADY(sum_3_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_3_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_3_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_3_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_3_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_3_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_3_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_3_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_3_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_3_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_3_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_3_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_3_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_3_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_3_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_3_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_3_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_3_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_3_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_3_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_3_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_3_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_3_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_3_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_3_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_3_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_3_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_3_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_3_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_3_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_3_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_3_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_3_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_3_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_3_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_3_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_3_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_3_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_3_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_3_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_3_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_3_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_3_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_3_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_3_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_3_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_3_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_3_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_3_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_3_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_3_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_3_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_3_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_3_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_3_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_3_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_3_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_3_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_3_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_3_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_3_m_axi_gmem_BUSER)
	);
	sum peArray_4_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_68_TREADY),
		.argOut_TVALID(_peArray_4_1_argOut_TVALID),
		.argOut_TDATA(_peArray_4_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_4_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_4_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_4_TDATA),
		.s_axi_control_ARREADY(sum_4_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_4_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_4_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_4_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_4_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_4_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_4_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_4_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_4_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_4_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_4_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_4_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_4_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_4_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_4_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_4_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_4_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_4_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_4_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_4_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_4_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_4_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_4_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_4_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_4_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_4_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_4_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_4_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_4_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_4_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_4_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_4_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_4_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_4_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_4_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_4_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_4_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_4_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_4_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_4_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_4_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_4_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_4_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_4_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_4_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_4_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_4_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_4_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_4_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_4_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_4_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_4_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_4_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_4_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_4_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_4_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_4_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_4_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_4_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_4_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_4_m_axi_gmem_BUSER)
	);
	sum peArray_5_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_69_TREADY),
		.argOut_TVALID(_peArray_5_1_argOut_TVALID),
		.argOut_TDATA(_peArray_5_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_5_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_5_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_5_TDATA),
		.s_axi_control_ARREADY(sum_5_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_5_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_5_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_5_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_5_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_5_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_5_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_5_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_5_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_5_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_5_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_5_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_5_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_5_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_5_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_5_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_5_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_5_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_5_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_5_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_5_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_5_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_5_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_5_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_5_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_5_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_5_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_5_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_5_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_5_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_5_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_5_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_5_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_5_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_5_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_5_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_5_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_5_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_5_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_5_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_5_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_5_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_5_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_5_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_5_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_5_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_5_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_5_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_5_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_5_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_5_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_5_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_5_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_5_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_5_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_5_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_5_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_5_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_5_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_5_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_5_m_axi_gmem_BUSER)
	);
	sum peArray_6_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_70_TREADY),
		.argOut_TVALID(_peArray_6_1_argOut_TVALID),
		.argOut_TDATA(_peArray_6_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_6_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_6_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_6_TDATA),
		.s_axi_control_ARREADY(sum_6_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_6_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_6_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_6_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_6_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_6_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_6_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_6_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_6_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_6_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_6_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_6_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_6_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_6_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_6_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_6_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_6_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_6_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_6_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_6_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_6_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_6_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_6_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_6_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_6_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_6_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_6_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_6_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_6_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_6_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_6_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_6_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_6_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_6_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_6_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_6_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_6_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_6_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_6_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_6_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_6_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_6_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_6_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_6_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_6_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_6_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_6_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_6_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_6_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_6_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_6_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_6_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_6_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_6_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_6_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_6_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_6_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_6_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_6_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_6_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_6_m_axi_gmem_BUSER)
	);
	sum peArray_7_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_71_TREADY),
		.argOut_TVALID(_peArray_7_1_argOut_TVALID),
		.argOut_TDATA(_peArray_7_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_7_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_7_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_7_TDATA),
		.s_axi_control_ARREADY(sum_7_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_7_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_7_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_7_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_7_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_7_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_7_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_7_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_7_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_7_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_7_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_7_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_7_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_7_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_7_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_7_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_7_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_7_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_7_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_7_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_7_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_7_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_7_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_7_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_7_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_7_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_7_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_7_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_7_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_7_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_7_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_7_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_7_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_7_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_7_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_7_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_7_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_7_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_7_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_7_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_7_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_7_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_7_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_7_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_7_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_7_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_7_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_7_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_7_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_7_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_7_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_7_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_7_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_7_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_7_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_7_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_7_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_7_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_7_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_7_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_7_m_axi_gmem_BUSER)
	);
	sum peArray_8_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_72_TREADY),
		.argOut_TVALID(_peArray_8_1_argOut_TVALID),
		.argOut_TDATA(_peArray_8_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_8_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_8_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_8_TDATA),
		.s_axi_control_ARREADY(sum_8_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_8_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_8_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_8_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_8_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_8_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_8_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_8_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_8_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_8_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_8_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_8_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_8_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_8_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_8_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_8_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_8_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_8_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_8_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_8_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_8_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_8_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_8_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_8_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_8_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_8_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_8_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_8_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_8_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_8_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_8_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_8_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_8_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_8_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_8_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_8_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_8_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_8_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_8_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_8_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_8_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_8_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_8_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_8_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_8_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_8_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_8_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_8_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_8_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_8_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_8_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_8_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_8_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_8_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_8_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_8_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_8_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_8_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_8_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_8_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_8_m_axi_gmem_BUSER)
	);
	sum peArray_9_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_73_TREADY),
		.argOut_TVALID(_peArray_9_1_argOut_TVALID),
		.argOut_TDATA(_peArray_9_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_9_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_9_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_9_TDATA),
		.s_axi_control_ARREADY(sum_9_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_9_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_9_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_9_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_9_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_9_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_9_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_9_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_9_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_9_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_9_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_9_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_9_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_9_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_9_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_9_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_9_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_9_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_9_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_9_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_9_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_9_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_9_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_9_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_9_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_9_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_9_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_9_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_9_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_9_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_9_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_9_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_9_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_9_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_9_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_9_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_9_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_9_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_9_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_9_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_9_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_9_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_9_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_9_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_9_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_9_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_9_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_9_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_9_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_9_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_9_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_9_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_9_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_9_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_9_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_9_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_9_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_9_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_9_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_9_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_9_m_axi_gmem_BUSER)
	);
	sum peArray_10_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_74_TREADY),
		.argOut_TVALID(_peArray_10_1_argOut_TVALID),
		.argOut_TDATA(_peArray_10_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_10_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_10_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_10_TDATA),
		.s_axi_control_ARREADY(sum_10_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_10_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_10_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_10_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_10_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_10_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_10_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_10_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_10_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_10_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_10_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_10_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_10_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_10_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_10_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_10_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_10_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_10_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_10_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_10_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_10_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_10_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_10_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_10_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_10_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_10_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_10_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_10_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_10_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_10_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_10_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_10_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_10_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_10_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_10_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_10_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_10_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_10_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_10_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_10_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_10_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_10_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_10_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_10_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_10_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_10_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_10_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_10_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_10_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_10_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_10_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_10_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_10_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_10_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_10_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_10_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_10_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_10_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_10_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_10_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_10_m_axi_gmem_BUSER)
	);
	sum peArray_11_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_75_TREADY),
		.argOut_TVALID(_peArray_11_1_argOut_TVALID),
		.argOut_TDATA(_peArray_11_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_11_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_11_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_11_TDATA),
		.s_axi_control_ARREADY(sum_11_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_11_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_11_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_11_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_11_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_11_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_11_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_11_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_11_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_11_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_11_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_11_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_11_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_11_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_11_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_11_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_11_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_11_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_11_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_11_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_11_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_11_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_11_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_11_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_11_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_11_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_11_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_11_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_11_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_11_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_11_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_11_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_11_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_11_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_11_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_11_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_11_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_11_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_11_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_11_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_11_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_11_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_11_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_11_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_11_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_11_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_11_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_11_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_11_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_11_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_11_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_11_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_11_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_11_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_11_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_11_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_11_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_11_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_11_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_11_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_11_m_axi_gmem_BUSER)
	);
	sum peArray_12_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_76_TREADY),
		.argOut_TVALID(_peArray_12_1_argOut_TVALID),
		.argOut_TDATA(_peArray_12_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_12_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_12_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_12_TDATA),
		.s_axi_control_ARREADY(sum_12_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_12_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_12_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_12_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_12_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_12_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_12_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_12_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_12_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_12_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_12_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_12_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_12_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_12_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_12_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_12_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_12_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_12_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_12_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_12_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_12_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_12_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_12_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_12_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_12_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_12_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_12_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_12_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_12_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_12_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_12_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_12_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_12_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_12_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_12_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_12_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_12_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_12_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_12_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_12_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_12_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_12_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_12_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_12_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_12_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_12_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_12_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_12_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_12_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_12_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_12_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_12_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_12_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_12_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_12_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_12_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_12_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_12_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_12_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_12_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_12_m_axi_gmem_BUSER)
	);
	sum peArray_13_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_77_TREADY),
		.argOut_TVALID(_peArray_13_1_argOut_TVALID),
		.argOut_TDATA(_peArray_13_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_13_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_13_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_13_TDATA),
		.s_axi_control_ARREADY(sum_13_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_13_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_13_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_13_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_13_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_13_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_13_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_13_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_13_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_13_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_13_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_13_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_13_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_13_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_13_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_13_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_13_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_13_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_13_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_13_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_13_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_13_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_13_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_13_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_13_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_13_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_13_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_13_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_13_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_13_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_13_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_13_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_13_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_13_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_13_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_13_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_13_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_13_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_13_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_13_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_13_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_13_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_13_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_13_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_13_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_13_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_13_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_13_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_13_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_13_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_13_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_13_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_13_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_13_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_13_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_13_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_13_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_13_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_13_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_13_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_13_m_axi_gmem_BUSER)
	);
	sum peArray_14_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_78_TREADY),
		.argOut_TVALID(_peArray_14_1_argOut_TVALID),
		.argOut_TDATA(_peArray_14_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_14_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_14_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_14_TDATA),
		.s_axi_control_ARREADY(sum_14_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_14_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_14_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_14_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_14_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_14_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_14_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_14_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_14_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_14_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_14_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_14_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_14_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_14_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_14_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_14_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_14_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_14_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_14_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_14_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_14_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_14_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_14_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_14_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_14_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_14_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_14_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_14_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_14_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_14_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_14_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_14_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_14_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_14_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_14_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_14_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_14_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_14_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_14_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_14_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_14_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_14_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_14_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_14_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_14_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_14_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_14_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_14_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_14_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_14_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_14_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_14_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_14_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_14_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_14_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_14_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_14_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_14_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_14_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_14_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_14_m_axi_gmem_BUSER)
	);
	sum peArray_15_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_79_TREADY),
		.argOut_TVALID(_peArray_15_1_argOut_TVALID),
		.argOut_TDATA(_peArray_15_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_15_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_15_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_15_TDATA),
		.s_axi_control_ARREADY(sum_15_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_15_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_15_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_15_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_15_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_15_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_15_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_15_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_15_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_15_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_15_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_15_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_15_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_15_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_15_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_15_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_15_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_15_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_15_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_15_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_15_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_15_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_15_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_15_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_15_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_15_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_15_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_15_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_15_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_15_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_15_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_15_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_15_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_15_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_15_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_15_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_15_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_15_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_15_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_15_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_15_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_15_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_15_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_15_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_15_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_15_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_15_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_15_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_15_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_15_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_15_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_15_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_15_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_15_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_15_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_15_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_15_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_15_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_15_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_15_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_15_m_axi_gmem_BUSER)
	);
	sum peArray_16_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_80_TREADY),
		.argOut_TVALID(_peArray_16_1_argOut_TVALID),
		.argOut_TDATA(_peArray_16_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_16_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_16_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_16_TDATA),
		.s_axi_control_ARREADY(sum_16_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_16_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_16_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_16_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_16_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_16_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_16_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_16_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_16_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_16_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_16_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_16_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_16_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_16_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_16_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_16_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_16_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_16_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_16_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_16_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_16_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_16_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_16_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_16_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_16_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_16_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_16_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_16_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_16_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_16_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_16_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_16_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_16_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_16_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_16_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_16_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_16_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_16_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_16_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_16_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_16_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_16_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_16_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_16_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_16_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_16_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_16_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_16_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_16_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_16_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_16_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_16_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_16_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_16_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_16_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_16_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_16_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_16_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_16_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_16_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_16_m_axi_gmem_BUSER)
	);
	sum peArray_17_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_81_TREADY),
		.argOut_TVALID(_peArray_17_1_argOut_TVALID),
		.argOut_TDATA(_peArray_17_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_17_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_17_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_17_TDATA),
		.s_axi_control_ARREADY(sum_17_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_17_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_17_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_17_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_17_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_17_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_17_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_17_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_17_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_17_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_17_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_17_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_17_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_17_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_17_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_17_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_17_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_17_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_17_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_17_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_17_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_17_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_17_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_17_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_17_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_17_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_17_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_17_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_17_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_17_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_17_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_17_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_17_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_17_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_17_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_17_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_17_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_17_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_17_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_17_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_17_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_17_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_17_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_17_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_17_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_17_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_17_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_17_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_17_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_17_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_17_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_17_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_17_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_17_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_17_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_17_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_17_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_17_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_17_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_17_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_17_m_axi_gmem_BUSER)
	);
	sum peArray_18_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_82_TREADY),
		.argOut_TVALID(_peArray_18_1_argOut_TVALID),
		.argOut_TDATA(_peArray_18_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_18_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_18_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_18_TDATA),
		.s_axi_control_ARREADY(sum_18_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_18_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_18_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_18_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_18_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_18_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_18_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_18_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_18_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_18_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_18_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_18_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_18_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_18_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_18_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_18_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_18_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_18_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_18_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_18_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_18_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_18_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_18_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_18_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_18_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_18_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_18_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_18_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_18_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_18_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_18_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_18_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_18_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_18_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_18_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_18_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_18_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_18_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_18_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_18_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_18_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_18_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_18_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_18_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_18_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_18_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_18_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_18_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_18_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_18_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_18_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_18_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_18_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_18_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_18_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_18_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_18_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_18_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_18_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_18_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_18_m_axi_gmem_BUSER)
	);
	sum peArray_19_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_83_TREADY),
		.argOut_TVALID(_peArray_19_1_argOut_TVALID),
		.argOut_TDATA(_peArray_19_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_19_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_19_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_19_TDATA),
		.s_axi_control_ARREADY(sum_19_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_19_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_19_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_19_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_19_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_19_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_19_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_19_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_19_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_19_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_19_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_19_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_19_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_19_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_19_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_19_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_19_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_19_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_19_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_19_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_19_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_19_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_19_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_19_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_19_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_19_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_19_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_19_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_19_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_19_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_19_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_19_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_19_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_19_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_19_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_19_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_19_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_19_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_19_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_19_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_19_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_19_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_19_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_19_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_19_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_19_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_19_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_19_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_19_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_19_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_19_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_19_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_19_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_19_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_19_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_19_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_19_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_19_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_19_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_19_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_19_m_axi_gmem_BUSER)
	);
	sum peArray_20_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_84_TREADY),
		.argOut_TVALID(_peArray_20_1_argOut_TVALID),
		.argOut_TDATA(_peArray_20_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_20_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_20_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_20_TDATA),
		.s_axi_control_ARREADY(sum_20_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_20_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_20_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_20_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_20_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_20_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_20_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_20_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_20_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_20_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_20_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_20_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_20_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_20_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_20_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_20_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_20_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_20_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_20_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_20_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_20_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_20_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_20_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_20_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_20_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_20_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_20_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_20_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_20_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_20_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_20_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_20_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_20_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_20_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_20_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_20_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_20_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_20_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_20_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_20_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_20_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_20_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_20_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_20_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_20_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_20_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_20_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_20_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_20_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_20_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_20_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_20_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_20_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_20_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_20_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_20_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_20_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_20_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_20_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_20_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_20_m_axi_gmem_BUSER)
	);
	sum peArray_21_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_85_TREADY),
		.argOut_TVALID(_peArray_21_1_argOut_TVALID),
		.argOut_TDATA(_peArray_21_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_21_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_21_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_21_TDATA),
		.s_axi_control_ARREADY(sum_21_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_21_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_21_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_21_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_21_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_21_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_21_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_21_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_21_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_21_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_21_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_21_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_21_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_21_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_21_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_21_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_21_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_21_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_21_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_21_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_21_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_21_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_21_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_21_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_21_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_21_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_21_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_21_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_21_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_21_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_21_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_21_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_21_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_21_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_21_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_21_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_21_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_21_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_21_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_21_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_21_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_21_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_21_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_21_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_21_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_21_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_21_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_21_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_21_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_21_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_21_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_21_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_21_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_21_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_21_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_21_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_21_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_21_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_21_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_21_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_21_m_axi_gmem_BUSER)
	);
	sum peArray_22_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_86_TREADY),
		.argOut_TVALID(_peArray_22_1_argOut_TVALID),
		.argOut_TDATA(_peArray_22_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_22_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_22_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_22_TDATA),
		.s_axi_control_ARREADY(sum_22_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_22_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_22_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_22_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_22_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_22_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_22_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_22_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_22_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_22_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_22_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_22_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_22_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_22_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_22_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_22_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_22_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_22_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_22_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_22_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_22_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_22_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_22_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_22_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_22_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_22_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_22_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_22_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_22_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_22_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_22_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_22_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_22_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_22_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_22_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_22_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_22_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_22_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_22_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_22_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_22_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_22_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_22_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_22_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_22_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_22_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_22_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_22_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_22_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_22_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_22_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_22_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_22_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_22_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_22_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_22_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_22_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_22_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_22_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_22_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_22_m_axi_gmem_BUSER)
	);
	sum peArray_23_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_87_TREADY),
		.argOut_TVALID(_peArray_23_1_argOut_TVALID),
		.argOut_TDATA(_peArray_23_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_23_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_23_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_23_TDATA),
		.s_axi_control_ARREADY(sum_23_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_23_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_23_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_23_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_23_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_23_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_23_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_23_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_23_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_23_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_23_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_23_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_23_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_23_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_23_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_23_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_23_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_23_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_23_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_23_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_23_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_23_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_23_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_23_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_23_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_23_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_23_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_23_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_23_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_23_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_23_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_23_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_23_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_23_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_23_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_23_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_23_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_23_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_23_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_23_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_23_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_23_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_23_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_23_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_23_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_23_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_23_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_23_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_23_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_23_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_23_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_23_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_23_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_23_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_23_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_23_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_23_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_23_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_23_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_23_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_23_m_axi_gmem_BUSER)
	);
	sum peArray_24_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_88_TREADY),
		.argOut_TVALID(_peArray_24_1_argOut_TVALID),
		.argOut_TDATA(_peArray_24_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_24_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_24_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_24_TDATA),
		.s_axi_control_ARREADY(sum_24_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_24_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_24_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_24_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_24_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_24_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_24_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_24_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_24_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_24_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_24_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_24_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_24_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_24_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_24_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_24_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_24_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_24_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_24_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_24_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_24_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_24_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_24_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_24_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_24_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_24_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_24_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_24_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_24_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_24_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_24_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_24_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_24_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_24_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_24_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_24_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_24_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_24_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_24_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_24_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_24_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_24_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_24_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_24_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_24_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_24_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_24_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_24_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_24_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_24_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_24_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_24_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_24_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_24_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_24_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_24_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_24_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_24_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_24_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_24_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_24_m_axi_gmem_BUSER)
	);
	sum peArray_25_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_89_TREADY),
		.argOut_TVALID(_peArray_25_1_argOut_TVALID),
		.argOut_TDATA(_peArray_25_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_25_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_25_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_25_TDATA),
		.s_axi_control_ARREADY(sum_25_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_25_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_25_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_25_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_25_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_25_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_25_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_25_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_25_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_25_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_25_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_25_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_25_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_25_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_25_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_25_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_25_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_25_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_25_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_25_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_25_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_25_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_25_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_25_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_25_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_25_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_25_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_25_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_25_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_25_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_25_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_25_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_25_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_25_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_25_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_25_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_25_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_25_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_25_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_25_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_25_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_25_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_25_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_25_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_25_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_25_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_25_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_25_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_25_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_25_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_25_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_25_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_25_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_25_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_25_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_25_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_25_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_25_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_25_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_25_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_25_m_axi_gmem_BUSER)
	);
	sum peArray_26_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_90_TREADY),
		.argOut_TVALID(_peArray_26_1_argOut_TVALID),
		.argOut_TDATA(_peArray_26_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_26_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_26_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_26_TDATA),
		.s_axi_control_ARREADY(sum_26_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_26_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_26_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_26_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_26_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_26_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_26_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_26_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_26_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_26_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_26_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_26_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_26_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_26_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_26_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_26_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_26_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_26_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_26_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_26_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_26_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_26_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_26_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_26_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_26_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_26_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_26_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_26_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_26_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_26_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_26_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_26_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_26_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_26_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_26_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_26_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_26_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_26_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_26_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_26_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_26_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_26_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_26_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_26_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_26_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_26_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_26_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_26_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_26_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_26_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_26_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_26_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_26_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_26_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_26_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_26_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_26_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_26_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_26_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_26_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_26_m_axi_gmem_BUSER)
	);
	sum peArray_27_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_91_TREADY),
		.argOut_TVALID(_peArray_27_1_argOut_TVALID),
		.argOut_TDATA(_peArray_27_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_27_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_27_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_27_TDATA),
		.s_axi_control_ARREADY(sum_27_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_27_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_27_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_27_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_27_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_27_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_27_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_27_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_27_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_27_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_27_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_27_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_27_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_27_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_27_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_27_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_27_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_27_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_27_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_27_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_27_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_27_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_27_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_27_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_27_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_27_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_27_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_27_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_27_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_27_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_27_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_27_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_27_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_27_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_27_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_27_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_27_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_27_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_27_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_27_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_27_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_27_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_27_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_27_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_27_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_27_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_27_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_27_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_27_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_27_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_27_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_27_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_27_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_27_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_27_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_27_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_27_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_27_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_27_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_27_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_27_m_axi_gmem_BUSER)
	);
	sum peArray_28_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_92_TREADY),
		.argOut_TVALID(_peArray_28_1_argOut_TVALID),
		.argOut_TDATA(_peArray_28_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_28_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_28_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_28_TDATA),
		.s_axi_control_ARREADY(sum_28_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_28_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_28_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_28_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_28_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_28_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_28_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_28_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_28_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_28_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_28_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_28_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_28_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_28_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_28_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_28_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_28_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_28_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_28_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_28_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_28_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_28_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_28_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_28_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_28_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_28_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_28_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_28_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_28_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_28_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_28_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_28_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_28_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_28_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_28_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_28_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_28_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_28_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_28_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_28_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_28_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_28_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_28_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_28_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_28_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_28_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_28_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_28_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_28_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_28_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_28_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_28_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_28_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_28_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_28_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_28_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_28_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_28_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_28_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_28_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_28_m_axi_gmem_BUSER)
	);
	sum peArray_29_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_93_TREADY),
		.argOut_TVALID(_peArray_29_1_argOut_TVALID),
		.argOut_TDATA(_peArray_29_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_29_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_29_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_29_TDATA),
		.s_axi_control_ARREADY(sum_29_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_29_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_29_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_29_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_29_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_29_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_29_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_29_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_29_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_29_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_29_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_29_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_29_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_29_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_29_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_29_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_29_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_29_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_29_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_29_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_29_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_29_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_29_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_29_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_29_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_29_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_29_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_29_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_29_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_29_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_29_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_29_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_29_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_29_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_29_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_29_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_29_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_29_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_29_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_29_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_29_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_29_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_29_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_29_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_29_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_29_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_29_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_29_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_29_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_29_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_29_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_29_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_29_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_29_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_29_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_29_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_29_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_29_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_29_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_29_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_29_m_axi_gmem_BUSER)
	);
	sum peArray_30_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_94_TREADY),
		.argOut_TVALID(_peArray_30_1_argOut_TVALID),
		.argOut_TDATA(_peArray_30_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_30_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_30_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_30_TDATA),
		.s_axi_control_ARREADY(sum_30_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_30_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_30_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_30_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_30_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_30_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_30_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_30_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_30_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_30_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_30_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_30_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_30_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_30_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_30_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_30_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_30_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_30_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_30_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_30_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_30_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_30_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_30_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_30_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_30_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_30_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_30_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_30_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_30_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_30_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_30_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_30_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_30_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_30_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_30_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_30_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_30_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_30_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_30_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_30_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_30_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_30_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_30_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_30_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_30_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_30_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_30_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_30_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_30_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_30_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_30_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_30_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_30_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_30_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_30_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_30_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_30_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_30_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_30_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_30_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_30_m_axi_gmem_BUSER)
	);
	sum peArray_31_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_95_TREADY),
		.argOut_TVALID(_peArray_31_1_argOut_TVALID),
		.argOut_TDATA(_peArray_31_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_31_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_31_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_31_TDATA),
		.s_axi_control_ARREADY(sum_31_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_31_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_31_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_31_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_31_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_31_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_31_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_31_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_31_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_31_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_31_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_31_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_31_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_31_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_31_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_31_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_31_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_31_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_31_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_31_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_31_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_31_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_31_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_31_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_31_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_31_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_31_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_31_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_31_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_31_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_31_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_31_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_31_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_31_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_31_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_31_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_31_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_31_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_31_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_31_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_31_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_31_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_31_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_31_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_31_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_31_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_31_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_31_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_31_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_31_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_31_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_31_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_31_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_31_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_31_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_31_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_31_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_31_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_31_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_31_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_31_m_axi_gmem_BUSER)
	);
	sum peArray_32_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_96_TREADY),
		.argOut_TVALID(_peArray_32_1_argOut_TVALID),
		.argOut_TDATA(_peArray_32_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_32_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_32_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_32_TDATA),
		.s_axi_control_ARREADY(sum_32_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_32_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_32_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_32_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_32_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_32_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_32_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_32_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_32_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_32_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_32_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_32_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_32_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_32_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_32_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_32_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_32_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_32_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_32_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_32_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_32_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_32_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_32_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_32_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_32_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_32_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_32_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_32_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_32_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_32_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_32_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_32_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_32_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_32_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_32_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_32_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_32_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_32_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_32_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_32_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_32_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_32_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_32_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_32_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_32_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_32_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_32_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_32_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_32_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_32_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_32_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_32_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_32_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_32_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_32_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_32_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_32_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_32_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_32_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_32_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_32_m_axi_gmem_BUSER)
	);
	sum peArray_33_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_97_TREADY),
		.argOut_TVALID(_peArray_33_1_argOut_TVALID),
		.argOut_TDATA(_peArray_33_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_33_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_33_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_33_TDATA),
		.s_axi_control_ARREADY(sum_33_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_33_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_33_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_33_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_33_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_33_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_33_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_33_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_33_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_33_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_33_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_33_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_33_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_33_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_33_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_33_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_33_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_33_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_33_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_33_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_33_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_33_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_33_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_33_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_33_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_33_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_33_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_33_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_33_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_33_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_33_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_33_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_33_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_33_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_33_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_33_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_33_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_33_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_33_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_33_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_33_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_33_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_33_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_33_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_33_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_33_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_33_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_33_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_33_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_33_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_33_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_33_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_33_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_33_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_33_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_33_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_33_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_33_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_33_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_33_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_33_m_axi_gmem_BUSER)
	);
	sum peArray_34_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_98_TREADY),
		.argOut_TVALID(_peArray_34_1_argOut_TVALID),
		.argOut_TDATA(_peArray_34_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_34_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_34_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_34_TDATA),
		.s_axi_control_ARREADY(sum_34_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_34_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_34_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_34_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_34_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_34_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_34_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_34_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_34_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_34_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_34_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_34_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_34_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_34_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_34_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_34_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_34_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_34_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_34_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_34_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_34_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_34_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_34_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_34_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_34_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_34_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_34_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_34_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_34_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_34_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_34_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_34_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_34_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_34_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_34_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_34_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_34_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_34_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_34_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_34_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_34_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_34_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_34_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_34_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_34_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_34_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_34_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_34_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_34_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_34_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_34_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_34_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_34_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_34_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_34_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_34_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_34_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_34_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_34_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_34_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_34_m_axi_gmem_BUSER)
	);
	sum peArray_35_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_99_TREADY),
		.argOut_TVALID(_peArray_35_1_argOut_TVALID),
		.argOut_TDATA(_peArray_35_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_35_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_35_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_35_TDATA),
		.s_axi_control_ARREADY(sum_35_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_35_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_35_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_35_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_35_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_35_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_35_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_35_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_35_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_35_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_35_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_35_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_35_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_35_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_35_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_35_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_35_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_35_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_35_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_35_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_35_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_35_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_35_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_35_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_35_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_35_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_35_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_35_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_35_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_35_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_35_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_35_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_35_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_35_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_35_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_35_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_35_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_35_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_35_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_35_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_35_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_35_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_35_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_35_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_35_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_35_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_35_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_35_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_35_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_35_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_35_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_35_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_35_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_35_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_35_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_35_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_35_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_35_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_35_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_35_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_35_m_axi_gmem_BUSER)
	);
	sum peArray_36_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_100_TREADY),
		.argOut_TVALID(_peArray_36_1_argOut_TVALID),
		.argOut_TDATA(_peArray_36_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_36_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_36_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_36_TDATA),
		.s_axi_control_ARREADY(sum_36_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_36_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_36_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_36_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_36_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_36_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_36_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_36_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_36_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_36_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_36_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_36_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_36_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_36_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_36_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_36_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_36_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_36_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_36_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_36_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_36_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_36_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_36_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_36_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_36_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_36_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_36_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_36_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_36_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_36_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_36_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_36_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_36_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_36_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_36_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_36_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_36_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_36_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_36_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_36_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_36_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_36_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_36_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_36_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_36_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_36_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_36_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_36_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_36_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_36_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_36_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_36_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_36_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_36_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_36_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_36_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_36_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_36_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_36_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_36_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_36_m_axi_gmem_BUSER)
	);
	sum peArray_37_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_101_TREADY),
		.argOut_TVALID(_peArray_37_1_argOut_TVALID),
		.argOut_TDATA(_peArray_37_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_37_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_37_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_37_TDATA),
		.s_axi_control_ARREADY(sum_37_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_37_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_37_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_37_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_37_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_37_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_37_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_37_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_37_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_37_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_37_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_37_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_37_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_37_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_37_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_37_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_37_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_37_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_37_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_37_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_37_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_37_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_37_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_37_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_37_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_37_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_37_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_37_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_37_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_37_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_37_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_37_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_37_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_37_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_37_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_37_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_37_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_37_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_37_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_37_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_37_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_37_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_37_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_37_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_37_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_37_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_37_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_37_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_37_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_37_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_37_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_37_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_37_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_37_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_37_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_37_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_37_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_37_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_37_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_37_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_37_m_axi_gmem_BUSER)
	);
	sum peArray_38_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_102_TREADY),
		.argOut_TVALID(_peArray_38_1_argOut_TVALID),
		.argOut_TDATA(_peArray_38_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_38_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_38_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_38_TDATA),
		.s_axi_control_ARREADY(sum_38_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_38_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_38_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_38_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_38_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_38_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_38_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_38_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_38_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_38_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_38_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_38_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_38_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_38_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_38_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_38_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_38_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_38_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_38_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_38_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_38_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_38_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_38_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_38_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_38_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_38_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_38_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_38_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_38_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_38_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_38_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_38_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_38_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_38_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_38_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_38_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_38_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_38_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_38_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_38_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_38_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_38_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_38_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_38_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_38_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_38_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_38_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_38_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_38_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_38_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_38_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_38_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_38_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_38_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_38_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_38_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_38_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_38_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_38_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_38_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_38_m_axi_gmem_BUSER)
	);
	sum peArray_39_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_103_TREADY),
		.argOut_TVALID(_peArray_39_1_argOut_TVALID),
		.argOut_TDATA(_peArray_39_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_39_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_39_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_39_TDATA),
		.s_axi_control_ARREADY(sum_39_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_39_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_39_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_39_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_39_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_39_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_39_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_39_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_39_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_39_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_39_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_39_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_39_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_39_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_39_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_39_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_39_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_39_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_39_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_39_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_39_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_39_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_39_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_39_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_39_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_39_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_39_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_39_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_39_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_39_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_39_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_39_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_39_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_39_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_39_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_39_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_39_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_39_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_39_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_39_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_39_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_39_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_39_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_39_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_39_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_39_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_39_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_39_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_39_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_39_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_39_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_39_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_39_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_39_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_39_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_39_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_39_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_39_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_39_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_39_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_39_m_axi_gmem_BUSER)
	);
	sum peArray_40_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_104_TREADY),
		.argOut_TVALID(_peArray_40_1_argOut_TVALID),
		.argOut_TDATA(_peArray_40_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_40_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_40_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_40_TDATA),
		.s_axi_control_ARREADY(sum_40_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_40_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_40_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_40_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_40_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_40_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_40_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_40_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_40_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_40_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_40_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_40_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_40_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_40_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_40_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_40_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_40_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_40_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_40_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_40_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_40_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_40_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_40_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_40_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_40_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_40_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_40_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_40_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_40_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_40_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_40_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_40_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_40_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_40_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_40_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_40_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_40_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_40_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_40_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_40_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_40_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_40_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_40_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_40_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_40_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_40_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_40_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_40_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_40_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_40_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_40_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_40_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_40_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_40_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_40_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_40_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_40_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_40_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_40_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_40_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_40_m_axi_gmem_BUSER)
	);
	sum peArray_41_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_105_TREADY),
		.argOut_TVALID(_peArray_41_1_argOut_TVALID),
		.argOut_TDATA(_peArray_41_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_41_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_41_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_41_TDATA),
		.s_axi_control_ARREADY(sum_41_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_41_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_41_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_41_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_41_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_41_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_41_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_41_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_41_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_41_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_41_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_41_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_41_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_41_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_41_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_41_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_41_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_41_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_41_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_41_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_41_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_41_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_41_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_41_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_41_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_41_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_41_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_41_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_41_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_41_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_41_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_41_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_41_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_41_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_41_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_41_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_41_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_41_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_41_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_41_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_41_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_41_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_41_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_41_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_41_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_41_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_41_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_41_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_41_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_41_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_41_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_41_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_41_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_41_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_41_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_41_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_41_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_41_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_41_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_41_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_41_m_axi_gmem_BUSER)
	);
	sum peArray_42_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_106_TREADY),
		.argOut_TVALID(_peArray_42_1_argOut_TVALID),
		.argOut_TDATA(_peArray_42_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_42_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_42_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_42_TDATA),
		.s_axi_control_ARREADY(sum_42_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_42_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_42_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_42_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_42_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_42_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_42_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_42_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_42_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_42_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_42_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_42_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_42_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_42_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_42_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_42_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_42_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_42_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_42_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_42_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_42_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_42_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_42_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_42_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_42_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_42_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_42_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_42_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_42_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_42_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_42_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_42_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_42_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_42_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_42_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_42_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_42_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_42_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_42_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_42_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_42_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_42_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_42_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_42_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_42_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_42_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_42_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_42_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_42_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_42_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_42_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_42_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_42_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_42_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_42_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_42_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_42_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_42_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_42_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_42_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_42_m_axi_gmem_BUSER)
	);
	sum peArray_43_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_107_TREADY),
		.argOut_TVALID(_peArray_43_1_argOut_TVALID),
		.argOut_TDATA(_peArray_43_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_43_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_43_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_43_TDATA),
		.s_axi_control_ARREADY(sum_43_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_43_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_43_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_43_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_43_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_43_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_43_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_43_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_43_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_43_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_43_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_43_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_43_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_43_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_43_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_43_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_43_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_43_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_43_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_43_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_43_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_43_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_43_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_43_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_43_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_43_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_43_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_43_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_43_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_43_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_43_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_43_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_43_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_43_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_43_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_43_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_43_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_43_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_43_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_43_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_43_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_43_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_43_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_43_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_43_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_43_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_43_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_43_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_43_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_43_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_43_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_43_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_43_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_43_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_43_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_43_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_43_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_43_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_43_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_43_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_43_m_axi_gmem_BUSER)
	);
	sum peArray_44_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_108_TREADY),
		.argOut_TVALID(_peArray_44_1_argOut_TVALID),
		.argOut_TDATA(_peArray_44_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_44_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_44_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_44_TDATA),
		.s_axi_control_ARREADY(sum_44_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_44_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_44_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_44_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_44_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_44_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_44_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_44_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_44_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_44_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_44_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_44_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_44_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_44_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_44_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_44_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_44_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_44_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_44_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_44_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_44_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_44_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_44_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_44_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_44_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_44_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_44_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_44_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_44_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_44_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_44_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_44_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_44_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_44_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_44_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_44_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_44_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_44_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_44_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_44_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_44_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_44_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_44_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_44_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_44_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_44_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_44_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_44_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_44_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_44_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_44_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_44_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_44_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_44_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_44_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_44_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_44_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_44_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_44_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_44_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_44_m_axi_gmem_BUSER)
	);
	sum peArray_45_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_109_TREADY),
		.argOut_TVALID(_peArray_45_1_argOut_TVALID),
		.argOut_TDATA(_peArray_45_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_45_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_45_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_45_TDATA),
		.s_axi_control_ARREADY(sum_45_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_45_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_45_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_45_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_45_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_45_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_45_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_45_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_45_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_45_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_45_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_45_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_45_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_45_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_45_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_45_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_45_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_45_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_45_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_45_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_45_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_45_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_45_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_45_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_45_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_45_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_45_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_45_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_45_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_45_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_45_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_45_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_45_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_45_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_45_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_45_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_45_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_45_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_45_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_45_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_45_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_45_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_45_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_45_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_45_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_45_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_45_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_45_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_45_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_45_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_45_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_45_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_45_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_45_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_45_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_45_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_45_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_45_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_45_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_45_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_45_m_axi_gmem_BUSER)
	);
	sum peArray_46_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_110_TREADY),
		.argOut_TVALID(_peArray_46_1_argOut_TVALID),
		.argOut_TDATA(_peArray_46_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_46_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_46_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_46_TDATA),
		.s_axi_control_ARREADY(sum_46_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_46_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_46_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_46_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_46_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_46_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_46_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_46_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_46_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_46_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_46_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_46_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_46_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_46_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_46_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_46_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_46_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_46_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_46_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_46_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_46_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_46_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_46_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_46_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_46_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_46_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_46_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_46_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_46_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_46_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_46_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_46_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_46_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_46_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_46_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_46_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_46_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_46_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_46_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_46_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_46_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_46_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_46_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_46_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_46_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_46_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_46_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_46_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_46_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_46_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_46_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_46_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_46_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_46_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_46_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_46_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_46_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_46_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_46_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_46_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_46_m_axi_gmem_BUSER)
	);
	sum peArray_47_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_111_TREADY),
		.argOut_TVALID(_peArray_47_1_argOut_TVALID),
		.argOut_TDATA(_peArray_47_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_47_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_47_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_47_TDATA),
		.s_axi_control_ARREADY(sum_47_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_47_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_47_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_47_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_47_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_47_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_47_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_47_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_47_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_47_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_47_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_47_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_47_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_47_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_47_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_47_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_47_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_47_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_47_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_47_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_47_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_47_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_47_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_47_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_47_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_47_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_47_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_47_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_47_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_47_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_47_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_47_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_47_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_47_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_47_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_47_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_47_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_47_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_47_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_47_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_47_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_47_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_47_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_47_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_47_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_47_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_47_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_47_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_47_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_47_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_47_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_47_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_47_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_47_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_47_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_47_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_47_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_47_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_47_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_47_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_47_m_axi_gmem_BUSER)
	);
	sum peArray_48_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_112_TREADY),
		.argOut_TVALID(_peArray_48_1_argOut_TVALID),
		.argOut_TDATA(_peArray_48_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_48_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_48_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_48_TDATA),
		.s_axi_control_ARREADY(sum_48_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_48_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_48_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_48_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_48_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_48_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_48_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_48_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_48_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_48_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_48_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_48_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_48_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_48_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_48_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_48_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_48_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_48_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_48_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_48_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_48_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_48_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_48_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_48_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_48_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_48_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_48_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_48_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_48_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_48_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_48_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_48_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_48_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_48_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_48_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_48_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_48_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_48_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_48_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_48_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_48_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_48_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_48_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_48_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_48_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_48_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_48_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_48_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_48_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_48_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_48_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_48_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_48_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_48_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_48_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_48_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_48_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_48_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_48_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_48_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_48_m_axi_gmem_BUSER)
	);
	sum peArray_49_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_113_TREADY),
		.argOut_TVALID(_peArray_49_1_argOut_TVALID),
		.argOut_TDATA(_peArray_49_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_49_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_49_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_49_TDATA),
		.s_axi_control_ARREADY(sum_49_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_49_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_49_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_49_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_49_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_49_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_49_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_49_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_49_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_49_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_49_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_49_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_49_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_49_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_49_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_49_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_49_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_49_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_49_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_49_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_49_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_49_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_49_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_49_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_49_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_49_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_49_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_49_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_49_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_49_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_49_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_49_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_49_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_49_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_49_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_49_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_49_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_49_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_49_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_49_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_49_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_49_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_49_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_49_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_49_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_49_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_49_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_49_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_49_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_49_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_49_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_49_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_49_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_49_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_49_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_49_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_49_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_49_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_49_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_49_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_49_m_axi_gmem_BUSER)
	);
	sum peArray_50_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_114_TREADY),
		.argOut_TVALID(_peArray_50_1_argOut_TVALID),
		.argOut_TDATA(_peArray_50_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_50_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_50_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_50_TDATA),
		.s_axi_control_ARREADY(sum_50_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_50_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_50_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_50_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_50_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_50_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_50_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_50_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_50_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_50_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_50_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_50_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_50_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_50_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_50_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_50_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_50_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_50_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_50_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_50_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_50_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_50_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_50_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_50_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_50_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_50_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_50_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_50_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_50_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_50_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_50_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_50_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_50_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_50_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_50_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_50_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_50_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_50_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_50_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_50_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_50_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_50_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_50_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_50_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_50_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_50_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_50_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_50_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_50_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_50_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_50_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_50_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_50_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_50_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_50_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_50_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_50_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_50_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_50_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_50_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_50_m_axi_gmem_BUSER)
	);
	sum peArray_51_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_115_TREADY),
		.argOut_TVALID(_peArray_51_1_argOut_TVALID),
		.argOut_TDATA(_peArray_51_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_51_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_51_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_51_TDATA),
		.s_axi_control_ARREADY(sum_51_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_51_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_51_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_51_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_51_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_51_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_51_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_51_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_51_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_51_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_51_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_51_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_51_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_51_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_51_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_51_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_51_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_51_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_51_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_51_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_51_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_51_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_51_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_51_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_51_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_51_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_51_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_51_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_51_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_51_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_51_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_51_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_51_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_51_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_51_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_51_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_51_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_51_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_51_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_51_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_51_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_51_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_51_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_51_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_51_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_51_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_51_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_51_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_51_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_51_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_51_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_51_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_51_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_51_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_51_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_51_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_51_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_51_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_51_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_51_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_51_m_axi_gmem_BUSER)
	);
	sum peArray_52_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_116_TREADY),
		.argOut_TVALID(_peArray_52_1_argOut_TVALID),
		.argOut_TDATA(_peArray_52_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_52_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_52_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_52_TDATA),
		.s_axi_control_ARREADY(sum_52_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_52_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_52_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_52_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_52_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_52_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_52_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_52_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_52_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_52_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_52_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_52_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_52_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_52_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_52_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_52_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_52_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_52_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_52_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_52_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_52_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_52_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_52_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_52_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_52_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_52_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_52_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_52_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_52_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_52_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_52_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_52_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_52_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_52_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_52_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_52_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_52_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_52_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_52_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_52_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_52_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_52_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_52_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_52_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_52_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_52_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_52_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_52_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_52_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_52_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_52_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_52_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_52_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_52_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_52_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_52_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_52_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_52_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_52_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_52_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_52_m_axi_gmem_BUSER)
	);
	sum peArray_53_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_117_TREADY),
		.argOut_TVALID(_peArray_53_1_argOut_TVALID),
		.argOut_TDATA(_peArray_53_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_53_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_53_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_53_TDATA),
		.s_axi_control_ARREADY(sum_53_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_53_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_53_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_53_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_53_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_53_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_53_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_53_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_53_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_53_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_53_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_53_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_53_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_53_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_53_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_53_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_53_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_53_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_53_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_53_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_53_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_53_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_53_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_53_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_53_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_53_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_53_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_53_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_53_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_53_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_53_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_53_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_53_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_53_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_53_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_53_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_53_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_53_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_53_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_53_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_53_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_53_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_53_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_53_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_53_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_53_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_53_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_53_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_53_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_53_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_53_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_53_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_53_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_53_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_53_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_53_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_53_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_53_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_53_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_53_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_53_m_axi_gmem_BUSER)
	);
	sum peArray_54_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_118_TREADY),
		.argOut_TVALID(_peArray_54_1_argOut_TVALID),
		.argOut_TDATA(_peArray_54_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_54_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_54_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_54_TDATA),
		.s_axi_control_ARREADY(sum_54_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_54_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_54_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_54_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_54_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_54_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_54_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_54_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_54_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_54_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_54_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_54_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_54_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_54_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_54_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_54_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_54_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_54_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_54_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_54_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_54_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_54_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_54_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_54_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_54_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_54_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_54_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_54_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_54_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_54_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_54_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_54_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_54_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_54_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_54_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_54_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_54_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_54_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_54_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_54_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_54_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_54_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_54_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_54_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_54_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_54_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_54_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_54_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_54_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_54_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_54_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_54_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_54_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_54_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_54_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_54_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_54_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_54_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_54_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_54_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_54_m_axi_gmem_BUSER)
	);
	sum peArray_55_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_119_TREADY),
		.argOut_TVALID(_peArray_55_1_argOut_TVALID),
		.argOut_TDATA(_peArray_55_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_55_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_55_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_55_TDATA),
		.s_axi_control_ARREADY(sum_55_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_55_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_55_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_55_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_55_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_55_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_55_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_55_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_55_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_55_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_55_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_55_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_55_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_55_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_55_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_55_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_55_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_55_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_55_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_55_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_55_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_55_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_55_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_55_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_55_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_55_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_55_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_55_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_55_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_55_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_55_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_55_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_55_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_55_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_55_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_55_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_55_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_55_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_55_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_55_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_55_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_55_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_55_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_55_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_55_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_55_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_55_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_55_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_55_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_55_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_55_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_55_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_55_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_55_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_55_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_55_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_55_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_55_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_55_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_55_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_55_m_axi_gmem_BUSER)
	);
	sum peArray_56_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_120_TREADY),
		.argOut_TVALID(_peArray_56_1_argOut_TVALID),
		.argOut_TDATA(_peArray_56_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_56_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_56_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_56_TDATA),
		.s_axi_control_ARREADY(sum_56_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_56_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_56_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_56_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_56_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_56_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_56_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_56_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_56_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_56_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_56_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_56_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_56_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_56_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_56_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_56_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_56_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_56_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_56_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_56_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_56_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_56_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_56_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_56_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_56_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_56_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_56_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_56_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_56_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_56_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_56_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_56_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_56_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_56_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_56_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_56_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_56_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_56_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_56_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_56_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_56_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_56_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_56_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_56_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_56_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_56_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_56_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_56_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_56_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_56_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_56_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_56_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_56_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_56_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_56_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_56_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_56_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_56_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_56_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_56_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_56_m_axi_gmem_BUSER)
	);
	sum peArray_57_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_121_TREADY),
		.argOut_TVALID(_peArray_57_1_argOut_TVALID),
		.argOut_TDATA(_peArray_57_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_57_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_57_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_57_TDATA),
		.s_axi_control_ARREADY(sum_57_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_57_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_57_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_57_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_57_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_57_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_57_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_57_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_57_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_57_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_57_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_57_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_57_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_57_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_57_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_57_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_57_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_57_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_57_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_57_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_57_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_57_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_57_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_57_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_57_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_57_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_57_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_57_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_57_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_57_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_57_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_57_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_57_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_57_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_57_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_57_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_57_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_57_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_57_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_57_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_57_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_57_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_57_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_57_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_57_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_57_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_57_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_57_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_57_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_57_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_57_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_57_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_57_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_57_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_57_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_57_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_57_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_57_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_57_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_57_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_57_m_axi_gmem_BUSER)
	);
	sum peArray_58_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_122_TREADY),
		.argOut_TVALID(_peArray_58_1_argOut_TVALID),
		.argOut_TDATA(_peArray_58_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_58_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_58_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_58_TDATA),
		.s_axi_control_ARREADY(sum_58_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_58_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_58_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_58_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_58_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_58_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_58_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_58_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_58_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_58_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_58_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_58_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_58_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_58_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_58_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_58_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_58_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_58_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_58_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_58_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_58_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_58_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_58_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_58_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_58_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_58_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_58_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_58_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_58_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_58_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_58_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_58_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_58_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_58_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_58_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_58_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_58_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_58_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_58_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_58_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_58_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_58_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_58_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_58_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_58_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_58_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_58_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_58_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_58_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_58_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_58_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_58_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_58_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_58_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_58_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_58_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_58_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_58_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_58_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_58_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_58_m_axi_gmem_BUSER)
	);
	sum peArray_59_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_123_TREADY),
		.argOut_TVALID(_peArray_59_1_argOut_TVALID),
		.argOut_TDATA(_peArray_59_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_59_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_59_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_59_TDATA),
		.s_axi_control_ARREADY(sum_59_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_59_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_59_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_59_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_59_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_59_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_59_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_59_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_59_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_59_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_59_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_59_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_59_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_59_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_59_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_59_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_59_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_59_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_59_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_59_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_59_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_59_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_59_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_59_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_59_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_59_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_59_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_59_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_59_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_59_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_59_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_59_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_59_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_59_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_59_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_59_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_59_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_59_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_59_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_59_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_59_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_59_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_59_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_59_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_59_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_59_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_59_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_59_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_59_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_59_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_59_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_59_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_59_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_59_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_59_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_59_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_59_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_59_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_59_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_59_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_59_m_axi_gmem_BUSER)
	);
	sum peArray_60_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_124_TREADY),
		.argOut_TVALID(_peArray_60_1_argOut_TVALID),
		.argOut_TDATA(_peArray_60_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_60_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_60_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_60_TDATA),
		.s_axi_control_ARREADY(sum_60_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_60_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_60_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_60_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_60_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_60_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_60_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_60_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_60_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_60_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_60_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_60_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_60_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_60_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_60_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_60_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_60_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_60_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_60_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_60_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_60_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_60_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_60_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_60_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_60_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_60_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_60_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_60_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_60_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_60_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_60_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_60_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_60_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_60_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_60_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_60_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_60_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_60_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_60_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_60_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_60_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_60_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_60_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_60_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_60_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_60_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_60_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_60_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_60_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_60_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_60_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_60_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_60_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_60_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_60_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_60_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_60_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_60_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_60_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_60_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_60_m_axi_gmem_BUSER)
	);
	sum peArray_61_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_125_TREADY),
		.argOut_TVALID(_peArray_61_1_argOut_TVALID),
		.argOut_TDATA(_peArray_61_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_61_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_61_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_61_TDATA),
		.s_axi_control_ARREADY(sum_61_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_61_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_61_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_61_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_61_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_61_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_61_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_61_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_61_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_61_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_61_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_61_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_61_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_61_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_61_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_61_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_61_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_61_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_61_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_61_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_61_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_61_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_61_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_61_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_61_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_61_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_61_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_61_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_61_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_61_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_61_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_61_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_61_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_61_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_61_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_61_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_61_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_61_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_61_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_61_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_61_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_61_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_61_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_61_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_61_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_61_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_61_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_61_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_61_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_61_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_61_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_61_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_61_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_61_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_61_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_61_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_61_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_61_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_61_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_61_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_61_m_axi_gmem_BUSER)
	);
	sum peArray_62_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_126_TREADY),
		.argOut_TVALID(_peArray_62_1_argOut_TVALID),
		.argOut_TDATA(_peArray_62_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_62_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_62_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_62_TDATA),
		.s_axi_control_ARREADY(sum_62_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_62_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_62_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_62_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_62_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_62_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_62_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_62_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_62_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_62_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_62_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_62_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_62_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_62_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_62_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_62_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_62_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_62_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_62_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_62_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_62_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_62_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_62_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_62_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_62_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_62_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_62_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_62_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_62_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_62_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_62_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_62_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_62_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_62_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_62_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_62_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_62_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_62_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_62_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_62_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_62_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_62_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_62_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_62_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_62_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_62_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_62_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_62_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_62_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_62_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_62_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_62_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_62_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_62_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_62_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_62_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_62_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_62_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_62_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_62_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_62_m_axi_gmem_BUSER)
	);
	sum peArray_63_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_127_TREADY),
		.argOut_TVALID(_peArray_63_1_argOut_TVALID),
		.argOut_TDATA(_peArray_63_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_63_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_63_TVALID),
		.taskIn_TDATA(_Scheduler_1_io_export_taskOut_63_TDATA),
		.s_axi_control_ARREADY(sum_63_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(sum_63_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(sum_63_s_axi_control_ARADDR),
		.s_axi_control_RREADY(sum_63_s_axi_control_RREADY),
		.s_axi_control_RVALID(sum_63_s_axi_control_RVALID),
		.s_axi_control_RDATA(sum_63_s_axi_control_RDATA),
		.s_axi_control_RRESP(sum_63_s_axi_control_RRESP),
		.s_axi_control_AWREADY(sum_63_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(sum_63_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(sum_63_s_axi_control_AWADDR),
		.s_axi_control_WREADY(sum_63_s_axi_control_WREADY),
		.s_axi_control_WVALID(sum_63_s_axi_control_WVALID),
		.s_axi_control_WDATA(sum_63_s_axi_control_WDATA),
		.s_axi_control_WSTRB(sum_63_s_axi_control_WSTRB),
		.s_axi_control_BREADY(sum_63_s_axi_control_BREADY),
		.s_axi_control_BVALID(sum_63_s_axi_control_BVALID),
		.s_axi_control_BRESP(sum_63_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(sum_63_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(sum_63_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(sum_63_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(sum_63_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(sum_63_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(sum_63_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(sum_63_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(sum_63_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(sum_63_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(sum_63_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(sum_63_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(sum_63_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(sum_63_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(sum_63_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(sum_63_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(sum_63_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(sum_63_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(sum_63_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(sum_63_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(sum_63_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(sum_63_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(sum_63_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(sum_63_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(sum_63_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(sum_63_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(sum_63_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(sum_63_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(sum_63_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(sum_63_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(sum_63_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(sum_63_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(sum_63_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(sum_63_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(sum_63_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(sum_63_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(sum_63_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(sum_63_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(sum_63_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(sum_63_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(sum_63_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(sum_63_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(sum_63_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(sum_63_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(sum_63_m_axi_gmem_BUSER)
	);
	Scheduler_1 Scheduler_1(
		.clock(clock),
		.reset(reset),
		.io_export_taskOut_0_TREADY(_peArray_0_1_taskIn_TREADY),
		.io_export_taskOut_0_TVALID(_Scheduler_1_io_export_taskOut_0_TVALID),
		.io_export_taskOut_0_TDATA(_Scheduler_1_io_export_taskOut_0_TDATA),
		.io_export_taskOut_1_TREADY(_peArray_1_1_taskIn_TREADY),
		.io_export_taskOut_1_TVALID(_Scheduler_1_io_export_taskOut_1_TVALID),
		.io_export_taskOut_1_TDATA(_Scheduler_1_io_export_taskOut_1_TDATA),
		.io_export_taskOut_2_TREADY(_peArray_2_1_taskIn_TREADY),
		.io_export_taskOut_2_TVALID(_Scheduler_1_io_export_taskOut_2_TVALID),
		.io_export_taskOut_2_TDATA(_Scheduler_1_io_export_taskOut_2_TDATA),
		.io_export_taskOut_3_TREADY(_peArray_3_1_taskIn_TREADY),
		.io_export_taskOut_3_TVALID(_Scheduler_1_io_export_taskOut_3_TVALID),
		.io_export_taskOut_3_TDATA(_Scheduler_1_io_export_taskOut_3_TDATA),
		.io_export_taskOut_4_TREADY(_peArray_4_1_taskIn_TREADY),
		.io_export_taskOut_4_TVALID(_Scheduler_1_io_export_taskOut_4_TVALID),
		.io_export_taskOut_4_TDATA(_Scheduler_1_io_export_taskOut_4_TDATA),
		.io_export_taskOut_5_TREADY(_peArray_5_1_taskIn_TREADY),
		.io_export_taskOut_5_TVALID(_Scheduler_1_io_export_taskOut_5_TVALID),
		.io_export_taskOut_5_TDATA(_Scheduler_1_io_export_taskOut_5_TDATA),
		.io_export_taskOut_6_TREADY(_peArray_6_1_taskIn_TREADY),
		.io_export_taskOut_6_TVALID(_Scheduler_1_io_export_taskOut_6_TVALID),
		.io_export_taskOut_6_TDATA(_Scheduler_1_io_export_taskOut_6_TDATA),
		.io_export_taskOut_7_TREADY(_peArray_7_1_taskIn_TREADY),
		.io_export_taskOut_7_TVALID(_Scheduler_1_io_export_taskOut_7_TVALID),
		.io_export_taskOut_7_TDATA(_Scheduler_1_io_export_taskOut_7_TDATA),
		.io_export_taskOut_8_TREADY(_peArray_8_1_taskIn_TREADY),
		.io_export_taskOut_8_TVALID(_Scheduler_1_io_export_taskOut_8_TVALID),
		.io_export_taskOut_8_TDATA(_Scheduler_1_io_export_taskOut_8_TDATA),
		.io_export_taskOut_9_TREADY(_peArray_9_1_taskIn_TREADY),
		.io_export_taskOut_9_TVALID(_Scheduler_1_io_export_taskOut_9_TVALID),
		.io_export_taskOut_9_TDATA(_Scheduler_1_io_export_taskOut_9_TDATA),
		.io_export_taskOut_10_TREADY(_peArray_10_1_taskIn_TREADY),
		.io_export_taskOut_10_TVALID(_Scheduler_1_io_export_taskOut_10_TVALID),
		.io_export_taskOut_10_TDATA(_Scheduler_1_io_export_taskOut_10_TDATA),
		.io_export_taskOut_11_TREADY(_peArray_11_1_taskIn_TREADY),
		.io_export_taskOut_11_TVALID(_Scheduler_1_io_export_taskOut_11_TVALID),
		.io_export_taskOut_11_TDATA(_Scheduler_1_io_export_taskOut_11_TDATA),
		.io_export_taskOut_12_TREADY(_peArray_12_1_taskIn_TREADY),
		.io_export_taskOut_12_TVALID(_Scheduler_1_io_export_taskOut_12_TVALID),
		.io_export_taskOut_12_TDATA(_Scheduler_1_io_export_taskOut_12_TDATA),
		.io_export_taskOut_13_TREADY(_peArray_13_1_taskIn_TREADY),
		.io_export_taskOut_13_TVALID(_Scheduler_1_io_export_taskOut_13_TVALID),
		.io_export_taskOut_13_TDATA(_Scheduler_1_io_export_taskOut_13_TDATA),
		.io_export_taskOut_14_TREADY(_peArray_14_1_taskIn_TREADY),
		.io_export_taskOut_14_TVALID(_Scheduler_1_io_export_taskOut_14_TVALID),
		.io_export_taskOut_14_TDATA(_Scheduler_1_io_export_taskOut_14_TDATA),
		.io_export_taskOut_15_TREADY(_peArray_15_1_taskIn_TREADY),
		.io_export_taskOut_15_TVALID(_Scheduler_1_io_export_taskOut_15_TVALID),
		.io_export_taskOut_15_TDATA(_Scheduler_1_io_export_taskOut_15_TDATA),
		.io_export_taskOut_16_TREADY(_peArray_16_1_taskIn_TREADY),
		.io_export_taskOut_16_TVALID(_Scheduler_1_io_export_taskOut_16_TVALID),
		.io_export_taskOut_16_TDATA(_Scheduler_1_io_export_taskOut_16_TDATA),
		.io_export_taskOut_17_TREADY(_peArray_17_1_taskIn_TREADY),
		.io_export_taskOut_17_TVALID(_Scheduler_1_io_export_taskOut_17_TVALID),
		.io_export_taskOut_17_TDATA(_Scheduler_1_io_export_taskOut_17_TDATA),
		.io_export_taskOut_18_TREADY(_peArray_18_1_taskIn_TREADY),
		.io_export_taskOut_18_TVALID(_Scheduler_1_io_export_taskOut_18_TVALID),
		.io_export_taskOut_18_TDATA(_Scheduler_1_io_export_taskOut_18_TDATA),
		.io_export_taskOut_19_TREADY(_peArray_19_1_taskIn_TREADY),
		.io_export_taskOut_19_TVALID(_Scheduler_1_io_export_taskOut_19_TVALID),
		.io_export_taskOut_19_TDATA(_Scheduler_1_io_export_taskOut_19_TDATA),
		.io_export_taskOut_20_TREADY(_peArray_20_1_taskIn_TREADY),
		.io_export_taskOut_20_TVALID(_Scheduler_1_io_export_taskOut_20_TVALID),
		.io_export_taskOut_20_TDATA(_Scheduler_1_io_export_taskOut_20_TDATA),
		.io_export_taskOut_21_TREADY(_peArray_21_1_taskIn_TREADY),
		.io_export_taskOut_21_TVALID(_Scheduler_1_io_export_taskOut_21_TVALID),
		.io_export_taskOut_21_TDATA(_Scheduler_1_io_export_taskOut_21_TDATA),
		.io_export_taskOut_22_TREADY(_peArray_22_1_taskIn_TREADY),
		.io_export_taskOut_22_TVALID(_Scheduler_1_io_export_taskOut_22_TVALID),
		.io_export_taskOut_22_TDATA(_Scheduler_1_io_export_taskOut_22_TDATA),
		.io_export_taskOut_23_TREADY(_peArray_23_1_taskIn_TREADY),
		.io_export_taskOut_23_TVALID(_Scheduler_1_io_export_taskOut_23_TVALID),
		.io_export_taskOut_23_TDATA(_Scheduler_1_io_export_taskOut_23_TDATA),
		.io_export_taskOut_24_TREADY(_peArray_24_1_taskIn_TREADY),
		.io_export_taskOut_24_TVALID(_Scheduler_1_io_export_taskOut_24_TVALID),
		.io_export_taskOut_24_TDATA(_Scheduler_1_io_export_taskOut_24_TDATA),
		.io_export_taskOut_25_TREADY(_peArray_25_1_taskIn_TREADY),
		.io_export_taskOut_25_TVALID(_Scheduler_1_io_export_taskOut_25_TVALID),
		.io_export_taskOut_25_TDATA(_Scheduler_1_io_export_taskOut_25_TDATA),
		.io_export_taskOut_26_TREADY(_peArray_26_1_taskIn_TREADY),
		.io_export_taskOut_26_TVALID(_Scheduler_1_io_export_taskOut_26_TVALID),
		.io_export_taskOut_26_TDATA(_Scheduler_1_io_export_taskOut_26_TDATA),
		.io_export_taskOut_27_TREADY(_peArray_27_1_taskIn_TREADY),
		.io_export_taskOut_27_TVALID(_Scheduler_1_io_export_taskOut_27_TVALID),
		.io_export_taskOut_27_TDATA(_Scheduler_1_io_export_taskOut_27_TDATA),
		.io_export_taskOut_28_TREADY(_peArray_28_1_taskIn_TREADY),
		.io_export_taskOut_28_TVALID(_Scheduler_1_io_export_taskOut_28_TVALID),
		.io_export_taskOut_28_TDATA(_Scheduler_1_io_export_taskOut_28_TDATA),
		.io_export_taskOut_29_TREADY(_peArray_29_1_taskIn_TREADY),
		.io_export_taskOut_29_TVALID(_Scheduler_1_io_export_taskOut_29_TVALID),
		.io_export_taskOut_29_TDATA(_Scheduler_1_io_export_taskOut_29_TDATA),
		.io_export_taskOut_30_TREADY(_peArray_30_1_taskIn_TREADY),
		.io_export_taskOut_30_TVALID(_Scheduler_1_io_export_taskOut_30_TVALID),
		.io_export_taskOut_30_TDATA(_Scheduler_1_io_export_taskOut_30_TDATA),
		.io_export_taskOut_31_TREADY(_peArray_31_1_taskIn_TREADY),
		.io_export_taskOut_31_TVALID(_Scheduler_1_io_export_taskOut_31_TVALID),
		.io_export_taskOut_31_TDATA(_Scheduler_1_io_export_taskOut_31_TDATA),
		.io_export_taskOut_32_TREADY(_peArray_32_1_taskIn_TREADY),
		.io_export_taskOut_32_TVALID(_Scheduler_1_io_export_taskOut_32_TVALID),
		.io_export_taskOut_32_TDATA(_Scheduler_1_io_export_taskOut_32_TDATA),
		.io_export_taskOut_33_TREADY(_peArray_33_1_taskIn_TREADY),
		.io_export_taskOut_33_TVALID(_Scheduler_1_io_export_taskOut_33_TVALID),
		.io_export_taskOut_33_TDATA(_Scheduler_1_io_export_taskOut_33_TDATA),
		.io_export_taskOut_34_TREADY(_peArray_34_1_taskIn_TREADY),
		.io_export_taskOut_34_TVALID(_Scheduler_1_io_export_taskOut_34_TVALID),
		.io_export_taskOut_34_TDATA(_Scheduler_1_io_export_taskOut_34_TDATA),
		.io_export_taskOut_35_TREADY(_peArray_35_1_taskIn_TREADY),
		.io_export_taskOut_35_TVALID(_Scheduler_1_io_export_taskOut_35_TVALID),
		.io_export_taskOut_35_TDATA(_Scheduler_1_io_export_taskOut_35_TDATA),
		.io_export_taskOut_36_TREADY(_peArray_36_1_taskIn_TREADY),
		.io_export_taskOut_36_TVALID(_Scheduler_1_io_export_taskOut_36_TVALID),
		.io_export_taskOut_36_TDATA(_Scheduler_1_io_export_taskOut_36_TDATA),
		.io_export_taskOut_37_TREADY(_peArray_37_1_taskIn_TREADY),
		.io_export_taskOut_37_TVALID(_Scheduler_1_io_export_taskOut_37_TVALID),
		.io_export_taskOut_37_TDATA(_Scheduler_1_io_export_taskOut_37_TDATA),
		.io_export_taskOut_38_TREADY(_peArray_38_1_taskIn_TREADY),
		.io_export_taskOut_38_TVALID(_Scheduler_1_io_export_taskOut_38_TVALID),
		.io_export_taskOut_38_TDATA(_Scheduler_1_io_export_taskOut_38_TDATA),
		.io_export_taskOut_39_TREADY(_peArray_39_1_taskIn_TREADY),
		.io_export_taskOut_39_TVALID(_Scheduler_1_io_export_taskOut_39_TVALID),
		.io_export_taskOut_39_TDATA(_Scheduler_1_io_export_taskOut_39_TDATA),
		.io_export_taskOut_40_TREADY(_peArray_40_1_taskIn_TREADY),
		.io_export_taskOut_40_TVALID(_Scheduler_1_io_export_taskOut_40_TVALID),
		.io_export_taskOut_40_TDATA(_Scheduler_1_io_export_taskOut_40_TDATA),
		.io_export_taskOut_41_TREADY(_peArray_41_1_taskIn_TREADY),
		.io_export_taskOut_41_TVALID(_Scheduler_1_io_export_taskOut_41_TVALID),
		.io_export_taskOut_41_TDATA(_Scheduler_1_io_export_taskOut_41_TDATA),
		.io_export_taskOut_42_TREADY(_peArray_42_1_taskIn_TREADY),
		.io_export_taskOut_42_TVALID(_Scheduler_1_io_export_taskOut_42_TVALID),
		.io_export_taskOut_42_TDATA(_Scheduler_1_io_export_taskOut_42_TDATA),
		.io_export_taskOut_43_TREADY(_peArray_43_1_taskIn_TREADY),
		.io_export_taskOut_43_TVALID(_Scheduler_1_io_export_taskOut_43_TVALID),
		.io_export_taskOut_43_TDATA(_Scheduler_1_io_export_taskOut_43_TDATA),
		.io_export_taskOut_44_TREADY(_peArray_44_1_taskIn_TREADY),
		.io_export_taskOut_44_TVALID(_Scheduler_1_io_export_taskOut_44_TVALID),
		.io_export_taskOut_44_TDATA(_Scheduler_1_io_export_taskOut_44_TDATA),
		.io_export_taskOut_45_TREADY(_peArray_45_1_taskIn_TREADY),
		.io_export_taskOut_45_TVALID(_Scheduler_1_io_export_taskOut_45_TVALID),
		.io_export_taskOut_45_TDATA(_Scheduler_1_io_export_taskOut_45_TDATA),
		.io_export_taskOut_46_TREADY(_peArray_46_1_taskIn_TREADY),
		.io_export_taskOut_46_TVALID(_Scheduler_1_io_export_taskOut_46_TVALID),
		.io_export_taskOut_46_TDATA(_Scheduler_1_io_export_taskOut_46_TDATA),
		.io_export_taskOut_47_TREADY(_peArray_47_1_taskIn_TREADY),
		.io_export_taskOut_47_TVALID(_Scheduler_1_io_export_taskOut_47_TVALID),
		.io_export_taskOut_47_TDATA(_Scheduler_1_io_export_taskOut_47_TDATA),
		.io_export_taskOut_48_TREADY(_peArray_48_1_taskIn_TREADY),
		.io_export_taskOut_48_TVALID(_Scheduler_1_io_export_taskOut_48_TVALID),
		.io_export_taskOut_48_TDATA(_Scheduler_1_io_export_taskOut_48_TDATA),
		.io_export_taskOut_49_TREADY(_peArray_49_1_taskIn_TREADY),
		.io_export_taskOut_49_TVALID(_Scheduler_1_io_export_taskOut_49_TVALID),
		.io_export_taskOut_49_TDATA(_Scheduler_1_io_export_taskOut_49_TDATA),
		.io_export_taskOut_50_TREADY(_peArray_50_1_taskIn_TREADY),
		.io_export_taskOut_50_TVALID(_Scheduler_1_io_export_taskOut_50_TVALID),
		.io_export_taskOut_50_TDATA(_Scheduler_1_io_export_taskOut_50_TDATA),
		.io_export_taskOut_51_TREADY(_peArray_51_1_taskIn_TREADY),
		.io_export_taskOut_51_TVALID(_Scheduler_1_io_export_taskOut_51_TVALID),
		.io_export_taskOut_51_TDATA(_Scheduler_1_io_export_taskOut_51_TDATA),
		.io_export_taskOut_52_TREADY(_peArray_52_1_taskIn_TREADY),
		.io_export_taskOut_52_TVALID(_Scheduler_1_io_export_taskOut_52_TVALID),
		.io_export_taskOut_52_TDATA(_Scheduler_1_io_export_taskOut_52_TDATA),
		.io_export_taskOut_53_TREADY(_peArray_53_1_taskIn_TREADY),
		.io_export_taskOut_53_TVALID(_Scheduler_1_io_export_taskOut_53_TVALID),
		.io_export_taskOut_53_TDATA(_Scheduler_1_io_export_taskOut_53_TDATA),
		.io_export_taskOut_54_TREADY(_peArray_54_1_taskIn_TREADY),
		.io_export_taskOut_54_TVALID(_Scheduler_1_io_export_taskOut_54_TVALID),
		.io_export_taskOut_54_TDATA(_Scheduler_1_io_export_taskOut_54_TDATA),
		.io_export_taskOut_55_TREADY(_peArray_55_1_taskIn_TREADY),
		.io_export_taskOut_55_TVALID(_Scheduler_1_io_export_taskOut_55_TVALID),
		.io_export_taskOut_55_TDATA(_Scheduler_1_io_export_taskOut_55_TDATA),
		.io_export_taskOut_56_TREADY(_peArray_56_1_taskIn_TREADY),
		.io_export_taskOut_56_TVALID(_Scheduler_1_io_export_taskOut_56_TVALID),
		.io_export_taskOut_56_TDATA(_Scheduler_1_io_export_taskOut_56_TDATA),
		.io_export_taskOut_57_TREADY(_peArray_57_1_taskIn_TREADY),
		.io_export_taskOut_57_TVALID(_Scheduler_1_io_export_taskOut_57_TVALID),
		.io_export_taskOut_57_TDATA(_Scheduler_1_io_export_taskOut_57_TDATA),
		.io_export_taskOut_58_TREADY(_peArray_58_1_taskIn_TREADY),
		.io_export_taskOut_58_TVALID(_Scheduler_1_io_export_taskOut_58_TVALID),
		.io_export_taskOut_58_TDATA(_Scheduler_1_io_export_taskOut_58_TDATA),
		.io_export_taskOut_59_TREADY(_peArray_59_1_taskIn_TREADY),
		.io_export_taskOut_59_TVALID(_Scheduler_1_io_export_taskOut_59_TVALID),
		.io_export_taskOut_59_TDATA(_Scheduler_1_io_export_taskOut_59_TDATA),
		.io_export_taskOut_60_TREADY(_peArray_60_1_taskIn_TREADY),
		.io_export_taskOut_60_TVALID(_Scheduler_1_io_export_taskOut_60_TVALID),
		.io_export_taskOut_60_TDATA(_Scheduler_1_io_export_taskOut_60_TDATA),
		.io_export_taskOut_61_TREADY(_peArray_61_1_taskIn_TREADY),
		.io_export_taskOut_61_TVALID(_Scheduler_1_io_export_taskOut_61_TVALID),
		.io_export_taskOut_61_TDATA(_Scheduler_1_io_export_taskOut_61_TDATA),
		.io_export_taskOut_62_TREADY(_peArray_62_1_taskIn_TREADY),
		.io_export_taskOut_62_TVALID(_Scheduler_1_io_export_taskOut_62_TVALID),
		.io_export_taskOut_62_TDATA(_Scheduler_1_io_export_taskOut_62_TDATA),
		.io_export_taskOut_63_TREADY(_peArray_63_1_taskIn_TREADY),
		.io_export_taskOut_63_TVALID(_Scheduler_1_io_export_taskOut_63_TVALID),
		.io_export_taskOut_63_TDATA(_Scheduler_1_io_export_taskOut_63_TDATA),
		.io_internal_vss_axi_full_0_ar_ready(sum_schedulerAXI_0_ARREADY),
		.io_internal_vss_axi_full_0_ar_valid(sum_schedulerAXI_0_ARVALID),
		.io_internal_vss_axi_full_0_ar_bits_id(sum_schedulerAXI_0_ARID),
		.io_internal_vss_axi_full_0_ar_bits_addr(sum_schedulerAXI_0_ARADDR),
		.io_internal_vss_axi_full_0_ar_bits_len(sum_schedulerAXI_0_ARLEN),
		.io_internal_vss_axi_full_0_ar_bits_size(sum_schedulerAXI_0_ARSIZE),
		.io_internal_vss_axi_full_0_ar_bits_burst(sum_schedulerAXI_0_ARBURST),
		.io_internal_vss_axi_full_0_ar_bits_lock(sum_schedulerAXI_0_ARLOCK),
		.io_internal_vss_axi_full_0_ar_bits_cache(sum_schedulerAXI_0_ARCACHE),
		.io_internal_vss_axi_full_0_ar_bits_prot(sum_schedulerAXI_0_ARPROT),
		.io_internal_vss_axi_full_0_ar_bits_qos(sum_schedulerAXI_0_ARQOS),
		.io_internal_vss_axi_full_0_ar_bits_region(sum_schedulerAXI_0_ARREGION),
		.io_internal_vss_axi_full_0_r_ready(sum_schedulerAXI_0_RREADY),
		.io_internal_vss_axi_full_0_r_valid(sum_schedulerAXI_0_RVALID),
		.io_internal_vss_axi_full_0_r_bits_id(sum_schedulerAXI_0_RID),
		.io_internal_vss_axi_full_0_r_bits_data(sum_schedulerAXI_0_RDATA),
		.io_internal_vss_axi_full_0_r_bits_resp(sum_schedulerAXI_0_RRESP),
		.io_internal_vss_axi_full_0_r_bits_last(sum_schedulerAXI_0_RLAST),
		.io_internal_vss_axi_full_0_aw_ready(sum_schedulerAXI_0_AWREADY),
		.io_internal_vss_axi_full_0_aw_valid(sum_schedulerAXI_0_AWVALID),
		.io_internal_vss_axi_full_0_aw_bits_id(sum_schedulerAXI_0_AWID),
		.io_internal_vss_axi_full_0_aw_bits_addr(sum_schedulerAXI_0_AWADDR),
		.io_internal_vss_axi_full_0_aw_bits_len(sum_schedulerAXI_0_AWLEN),
		.io_internal_vss_axi_full_0_aw_bits_size(sum_schedulerAXI_0_AWSIZE),
		.io_internal_vss_axi_full_0_aw_bits_burst(sum_schedulerAXI_0_AWBURST),
		.io_internal_vss_axi_full_0_aw_bits_lock(sum_schedulerAXI_0_AWLOCK),
		.io_internal_vss_axi_full_0_aw_bits_cache(sum_schedulerAXI_0_AWCACHE),
		.io_internal_vss_axi_full_0_aw_bits_prot(sum_schedulerAXI_0_AWPROT),
		.io_internal_vss_axi_full_0_aw_bits_qos(sum_schedulerAXI_0_AWQOS),
		.io_internal_vss_axi_full_0_aw_bits_region(sum_schedulerAXI_0_AWREGION),
		.io_internal_vss_axi_full_0_w_ready(sum_schedulerAXI_0_WREADY),
		.io_internal_vss_axi_full_0_w_valid(sum_schedulerAXI_0_WVALID),
		.io_internal_vss_axi_full_0_w_bits_data(sum_schedulerAXI_0_WDATA),
		.io_internal_vss_axi_full_0_w_bits_strb(sum_schedulerAXI_0_WSTRB),
		.io_internal_vss_axi_full_0_w_bits_last(sum_schedulerAXI_0_WLAST),
		.io_internal_vss_axi_full_0_b_ready(sum_schedulerAXI_0_BREADY),
		.io_internal_vss_axi_full_0_b_valid(sum_schedulerAXI_0_BVALID),
		.io_internal_vss_axi_full_0_b_bits_id(sum_schedulerAXI_0_BID),
		.io_internal_vss_axi_full_0_b_bits_resp(sum_schedulerAXI_0_BRESP),
		.io_internal_axi_mgmt_vss_0_ar_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_ar_ready),
		.io_internal_axi_mgmt_vss_0_ar_valid(_demux_m_axil_2_ar_valid),
		.io_internal_axi_mgmt_vss_0_ar_bits_addr(_demux_m_axil_2_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_ar_bits_prot(_demux_m_axil_2_ar_bits_prot),
		.io_internal_axi_mgmt_vss_0_r_ready(_demux_m_axil_2_r_ready),
		.io_internal_axi_mgmt_vss_0_r_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_valid),
		.io_internal_axi_mgmt_vss_0_r_bits_data(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_internal_axi_mgmt_vss_0_r_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_internal_axi_mgmt_vss_0_aw_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_aw_ready),
		.io_internal_axi_mgmt_vss_0_aw_valid(_demux_m_axil_2_aw_valid),
		.io_internal_axi_mgmt_vss_0_aw_bits_addr(_demux_m_axil_2_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_aw_bits_prot(_demux_m_axil_2_aw_bits_prot),
		.io_internal_axi_mgmt_vss_0_w_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_w_ready),
		.io_internal_axi_mgmt_vss_0_w_valid(_demux_m_axil_2_w_valid),
		.io_internal_axi_mgmt_vss_0_w_bits_data(_demux_m_axil_2_w_bits_data),
		.io_internal_axi_mgmt_vss_0_w_bits_strb(_demux_m_axil_2_w_bits_strb),
		.io_internal_axi_mgmt_vss_0_b_ready(_demux_m_axil_2_b_ready),
		.io_internal_axi_mgmt_vss_0_b_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_valid),
		.io_internal_axi_mgmt_vss_0_b_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.io_internal_axi_mgmt_vss_1_ar_ready(_Scheduler_1_io_internal_axi_mgmt_vss_1_ar_ready),
		.io_internal_axi_mgmt_vss_1_ar_valid(_demux_m_axil_3_ar_valid),
		.io_internal_axi_mgmt_vss_1_ar_bits_addr(_demux_m_axil_3_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_1_ar_bits_prot(_demux_m_axil_3_ar_bits_prot),
		.io_internal_axi_mgmt_vss_1_r_ready(_demux_m_axil_3_r_ready),
		.io_internal_axi_mgmt_vss_1_r_valid(_Scheduler_1_io_internal_axi_mgmt_vss_1_r_valid),
		.io_internal_axi_mgmt_vss_1_r_bits_data(_Scheduler_1_io_internal_axi_mgmt_vss_1_r_bits_data),
		.io_internal_axi_mgmt_vss_1_r_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_1_r_bits_resp),
		.io_internal_axi_mgmt_vss_1_aw_ready(_Scheduler_1_io_internal_axi_mgmt_vss_1_aw_ready),
		.io_internal_axi_mgmt_vss_1_aw_valid(_demux_m_axil_3_aw_valid),
		.io_internal_axi_mgmt_vss_1_aw_bits_addr(_demux_m_axil_3_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_1_aw_bits_prot(_demux_m_axil_3_aw_bits_prot),
		.io_internal_axi_mgmt_vss_1_w_ready(_Scheduler_1_io_internal_axi_mgmt_vss_1_w_ready),
		.io_internal_axi_mgmt_vss_1_w_valid(_demux_m_axil_3_w_valid),
		.io_internal_axi_mgmt_vss_1_w_bits_data(_demux_m_axil_3_w_bits_data),
		.io_internal_axi_mgmt_vss_1_w_bits_strb(_demux_m_axil_3_w_bits_strb),
		.io_internal_axi_mgmt_vss_1_b_ready(_demux_m_axil_3_b_ready),
		.io_internal_axi_mgmt_vss_1_b_valid(_Scheduler_1_io_internal_axi_mgmt_vss_1_b_valid),
		.io_internal_axi_mgmt_vss_1_b_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_1_b_bits_resp),
		.connArgumentNotifier_0_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_0_ctrl_serveStealReq_valid),
		.connArgumentNotifier_0_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_0_ctrl_serveStealReq_ready),
		.connArgumentNotifier_0_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_0_data_qOutTask_ready),
		.connArgumentNotifier_0_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_0_data_qOutTask_valid),
		.connArgumentNotifier_0_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_0_data_qOutTask_bits),
		.connArgumentNotifier_1_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_1_ctrl_serveStealReq_valid),
		.connArgumentNotifier_1_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_1_ctrl_serveStealReq_ready),
		.connArgumentNotifier_1_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_1_data_qOutTask_ready),
		.connArgumentNotifier_1_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_1_data_qOutTask_valid),
		.connArgumentNotifier_1_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_1_data_qOutTask_bits),
		.connArgumentNotifier_2_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_2_ctrl_serveStealReq_valid),
		.connArgumentNotifier_2_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_2_ctrl_serveStealReq_ready),
		.connArgumentNotifier_2_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_2_data_qOutTask_ready),
		.connArgumentNotifier_2_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_2_data_qOutTask_valid),
		.connArgumentNotifier_2_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_2_data_qOutTask_bits),
		.connArgumentNotifier_3_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_3_ctrl_serveStealReq_valid),
		.connArgumentNotifier_3_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_3_ctrl_serveStealReq_ready),
		.connArgumentNotifier_3_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_3_data_qOutTask_ready),
		.connArgumentNotifier_3_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_3_data_qOutTask_valid),
		.connArgumentNotifier_3_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_3_data_qOutTask_bits),
		.connArgumentNotifier_4_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_4_ctrl_serveStealReq_valid),
		.connArgumentNotifier_4_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_4_ctrl_serveStealReq_ready),
		.connArgumentNotifier_4_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_4_data_qOutTask_ready),
		.connArgumentNotifier_4_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_4_data_qOutTask_valid),
		.connArgumentNotifier_4_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_4_data_qOutTask_bits),
		.connArgumentNotifier_5_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_5_ctrl_serveStealReq_valid),
		.connArgumentNotifier_5_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_5_ctrl_serveStealReq_ready),
		.connArgumentNotifier_5_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_5_data_qOutTask_ready),
		.connArgumentNotifier_5_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_5_data_qOutTask_valid),
		.connArgumentNotifier_5_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_5_data_qOutTask_bits),
		.connArgumentNotifier_6_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_6_ctrl_serveStealReq_valid),
		.connArgumentNotifier_6_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_6_ctrl_serveStealReq_ready),
		.connArgumentNotifier_6_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_6_data_qOutTask_ready),
		.connArgumentNotifier_6_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_6_data_qOutTask_valid),
		.connArgumentNotifier_6_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_6_data_qOutTask_bits),
		.connArgumentNotifier_7_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_7_ctrl_serveStealReq_valid),
		.connArgumentNotifier_7_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_7_ctrl_serveStealReq_ready),
		.connArgumentNotifier_7_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_7_data_qOutTask_ready),
		.connArgumentNotifier_7_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_7_data_qOutTask_valid),
		.connArgumentNotifier_7_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_7_data_qOutTask_bits),
		.connArgumentNotifier_8_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_8_ctrl_serveStealReq_valid),
		.connArgumentNotifier_8_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_8_ctrl_serveStealReq_ready),
		.connArgumentNotifier_8_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_8_data_qOutTask_ready),
		.connArgumentNotifier_8_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_8_data_qOutTask_valid),
		.connArgumentNotifier_8_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_8_data_qOutTask_bits),
		.connArgumentNotifier_9_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_9_ctrl_serveStealReq_valid),
		.connArgumentNotifier_9_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_9_ctrl_serveStealReq_ready),
		.connArgumentNotifier_9_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_9_data_qOutTask_ready),
		.connArgumentNotifier_9_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_9_data_qOutTask_valid),
		.connArgumentNotifier_9_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_9_data_qOutTask_bits),
		.connArgumentNotifier_10_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_10_ctrl_serveStealReq_valid),
		.connArgumentNotifier_10_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_10_ctrl_serveStealReq_ready),
		.connArgumentNotifier_10_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_10_data_qOutTask_ready),
		.connArgumentNotifier_10_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_10_data_qOutTask_valid),
		.connArgumentNotifier_10_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_10_data_qOutTask_bits),
		.connArgumentNotifier_11_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_11_ctrl_serveStealReq_valid),
		.connArgumentNotifier_11_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_11_ctrl_serveStealReq_ready),
		.connArgumentNotifier_11_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_11_data_qOutTask_ready),
		.connArgumentNotifier_11_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_11_data_qOutTask_valid),
		.connArgumentNotifier_11_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_11_data_qOutTask_bits),
		.connArgumentNotifier_12_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_12_ctrl_serveStealReq_valid),
		.connArgumentNotifier_12_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_12_ctrl_serveStealReq_ready),
		.connArgumentNotifier_12_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_12_data_qOutTask_ready),
		.connArgumentNotifier_12_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_12_data_qOutTask_valid),
		.connArgumentNotifier_12_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_12_data_qOutTask_bits),
		.connArgumentNotifier_13_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_13_ctrl_serveStealReq_valid),
		.connArgumentNotifier_13_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_13_ctrl_serveStealReq_ready),
		.connArgumentNotifier_13_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_13_data_qOutTask_ready),
		.connArgumentNotifier_13_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_13_data_qOutTask_valid),
		.connArgumentNotifier_13_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_13_data_qOutTask_bits),
		.connArgumentNotifier_14_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_14_ctrl_serveStealReq_valid),
		.connArgumentNotifier_14_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_14_ctrl_serveStealReq_ready),
		.connArgumentNotifier_14_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_14_data_qOutTask_ready),
		.connArgumentNotifier_14_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_14_data_qOutTask_valid),
		.connArgumentNotifier_14_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_14_data_qOutTask_bits),
		.connArgumentNotifier_15_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_15_ctrl_serveStealReq_valid),
		.connArgumentNotifier_15_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_15_ctrl_serveStealReq_ready),
		.connArgumentNotifier_15_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_15_data_qOutTask_ready),
		.connArgumentNotifier_15_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_15_data_qOutTask_valid),
		.connArgumentNotifier_15_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_15_data_qOutTask_bits)
	);
	Allocator Allocator(
		.clock(clock),
		.reset(reset),
		.io_export_closureOut_0_TREADY(_peArray_0_closureIn_TREADY),
		.io_export_closureOut_0_TVALID(_Allocator_io_export_closureOut_0_TVALID),
		.io_export_closureOut_0_TDATA(_Allocator_io_export_closureOut_0_TDATA),
		.io_export_closureOut_1_TREADY(_peArray_1_closureIn_TREADY),
		.io_export_closureOut_1_TVALID(_Allocator_io_export_closureOut_1_TVALID),
		.io_export_closureOut_1_TDATA(_Allocator_io_export_closureOut_1_TDATA),
		.io_export_closureOut_2_TREADY(_peArray_2_closureIn_TREADY),
		.io_export_closureOut_2_TVALID(_Allocator_io_export_closureOut_2_TVALID),
		.io_export_closureOut_2_TDATA(_Allocator_io_export_closureOut_2_TDATA),
		.io_export_closureOut_3_TREADY(_peArray_3_closureIn_TREADY),
		.io_export_closureOut_3_TVALID(_Allocator_io_export_closureOut_3_TVALID),
		.io_export_closureOut_3_TDATA(_Allocator_io_export_closureOut_3_TDATA),
		.io_export_closureOut_4_TREADY(_peArray_4_closureIn_TREADY),
		.io_export_closureOut_4_TVALID(_Allocator_io_export_closureOut_4_TVALID),
		.io_export_closureOut_4_TDATA(_Allocator_io_export_closureOut_4_TDATA),
		.io_export_closureOut_5_TREADY(_peArray_5_closureIn_TREADY),
		.io_export_closureOut_5_TVALID(_Allocator_io_export_closureOut_5_TVALID),
		.io_export_closureOut_5_TDATA(_Allocator_io_export_closureOut_5_TDATA),
		.io_export_closureOut_6_TREADY(_peArray_6_closureIn_TREADY),
		.io_export_closureOut_6_TVALID(_Allocator_io_export_closureOut_6_TVALID),
		.io_export_closureOut_6_TDATA(_Allocator_io_export_closureOut_6_TDATA),
		.io_export_closureOut_7_TREADY(_peArray_7_closureIn_TREADY),
		.io_export_closureOut_7_TVALID(_Allocator_io_export_closureOut_7_TVALID),
		.io_export_closureOut_7_TDATA(_Allocator_io_export_closureOut_7_TDATA),
		.io_export_closureOut_8_TREADY(_peArray_8_closureIn_TREADY),
		.io_export_closureOut_8_TVALID(_Allocator_io_export_closureOut_8_TVALID),
		.io_export_closureOut_8_TDATA(_Allocator_io_export_closureOut_8_TDATA),
		.io_export_closureOut_9_TREADY(_peArray_9_closureIn_TREADY),
		.io_export_closureOut_9_TVALID(_Allocator_io_export_closureOut_9_TVALID),
		.io_export_closureOut_9_TDATA(_Allocator_io_export_closureOut_9_TDATA),
		.io_export_closureOut_10_TREADY(_peArray_10_closureIn_TREADY),
		.io_export_closureOut_10_TVALID(_Allocator_io_export_closureOut_10_TVALID),
		.io_export_closureOut_10_TDATA(_Allocator_io_export_closureOut_10_TDATA),
		.io_export_closureOut_11_TREADY(_peArray_11_closureIn_TREADY),
		.io_export_closureOut_11_TVALID(_Allocator_io_export_closureOut_11_TVALID),
		.io_export_closureOut_11_TDATA(_Allocator_io_export_closureOut_11_TDATA),
		.io_export_closureOut_12_TREADY(_peArray_12_closureIn_TREADY),
		.io_export_closureOut_12_TVALID(_Allocator_io_export_closureOut_12_TVALID),
		.io_export_closureOut_12_TDATA(_Allocator_io_export_closureOut_12_TDATA),
		.io_export_closureOut_13_TREADY(_peArray_13_closureIn_TREADY),
		.io_export_closureOut_13_TVALID(_Allocator_io_export_closureOut_13_TVALID),
		.io_export_closureOut_13_TDATA(_Allocator_io_export_closureOut_13_TDATA),
		.io_export_closureOut_14_TREADY(_peArray_14_closureIn_TREADY),
		.io_export_closureOut_14_TVALID(_Allocator_io_export_closureOut_14_TVALID),
		.io_export_closureOut_14_TDATA(_Allocator_io_export_closureOut_14_TDATA),
		.io_export_closureOut_15_TREADY(_peArray_15_closureIn_TREADY),
		.io_export_closureOut_15_TVALID(_Allocator_io_export_closureOut_15_TVALID),
		.io_export_closureOut_15_TDATA(_Allocator_io_export_closureOut_15_TDATA),
		.io_export_closureOut_16_TREADY(_peArray_16_closureIn_TREADY),
		.io_export_closureOut_16_TVALID(_Allocator_io_export_closureOut_16_TVALID),
		.io_export_closureOut_16_TDATA(_Allocator_io_export_closureOut_16_TDATA),
		.io_export_closureOut_17_TREADY(_peArray_17_closureIn_TREADY),
		.io_export_closureOut_17_TVALID(_Allocator_io_export_closureOut_17_TVALID),
		.io_export_closureOut_17_TDATA(_Allocator_io_export_closureOut_17_TDATA),
		.io_export_closureOut_18_TREADY(_peArray_18_closureIn_TREADY),
		.io_export_closureOut_18_TVALID(_Allocator_io_export_closureOut_18_TVALID),
		.io_export_closureOut_18_TDATA(_Allocator_io_export_closureOut_18_TDATA),
		.io_export_closureOut_19_TREADY(_peArray_19_closureIn_TREADY),
		.io_export_closureOut_19_TVALID(_Allocator_io_export_closureOut_19_TVALID),
		.io_export_closureOut_19_TDATA(_Allocator_io_export_closureOut_19_TDATA),
		.io_export_closureOut_20_TREADY(_peArray_20_closureIn_TREADY),
		.io_export_closureOut_20_TVALID(_Allocator_io_export_closureOut_20_TVALID),
		.io_export_closureOut_20_TDATA(_Allocator_io_export_closureOut_20_TDATA),
		.io_export_closureOut_21_TREADY(_peArray_21_closureIn_TREADY),
		.io_export_closureOut_21_TVALID(_Allocator_io_export_closureOut_21_TVALID),
		.io_export_closureOut_21_TDATA(_Allocator_io_export_closureOut_21_TDATA),
		.io_export_closureOut_22_TREADY(_peArray_22_closureIn_TREADY),
		.io_export_closureOut_22_TVALID(_Allocator_io_export_closureOut_22_TVALID),
		.io_export_closureOut_22_TDATA(_Allocator_io_export_closureOut_22_TDATA),
		.io_export_closureOut_23_TREADY(_peArray_23_closureIn_TREADY),
		.io_export_closureOut_23_TVALID(_Allocator_io_export_closureOut_23_TVALID),
		.io_export_closureOut_23_TDATA(_Allocator_io_export_closureOut_23_TDATA),
		.io_export_closureOut_24_TREADY(_peArray_24_closureIn_TREADY),
		.io_export_closureOut_24_TVALID(_Allocator_io_export_closureOut_24_TVALID),
		.io_export_closureOut_24_TDATA(_Allocator_io_export_closureOut_24_TDATA),
		.io_export_closureOut_25_TREADY(_peArray_25_closureIn_TREADY),
		.io_export_closureOut_25_TVALID(_Allocator_io_export_closureOut_25_TVALID),
		.io_export_closureOut_25_TDATA(_Allocator_io_export_closureOut_25_TDATA),
		.io_export_closureOut_26_TREADY(_peArray_26_closureIn_TREADY),
		.io_export_closureOut_26_TVALID(_Allocator_io_export_closureOut_26_TVALID),
		.io_export_closureOut_26_TDATA(_Allocator_io_export_closureOut_26_TDATA),
		.io_export_closureOut_27_TREADY(_peArray_27_closureIn_TREADY),
		.io_export_closureOut_27_TVALID(_Allocator_io_export_closureOut_27_TVALID),
		.io_export_closureOut_27_TDATA(_Allocator_io_export_closureOut_27_TDATA),
		.io_export_closureOut_28_TREADY(_peArray_28_closureIn_TREADY),
		.io_export_closureOut_28_TVALID(_Allocator_io_export_closureOut_28_TVALID),
		.io_export_closureOut_28_TDATA(_Allocator_io_export_closureOut_28_TDATA),
		.io_export_closureOut_29_TREADY(_peArray_29_closureIn_TREADY),
		.io_export_closureOut_29_TVALID(_Allocator_io_export_closureOut_29_TVALID),
		.io_export_closureOut_29_TDATA(_Allocator_io_export_closureOut_29_TDATA),
		.io_export_closureOut_30_TREADY(_peArray_30_closureIn_TREADY),
		.io_export_closureOut_30_TVALID(_Allocator_io_export_closureOut_30_TVALID),
		.io_export_closureOut_30_TDATA(_Allocator_io_export_closureOut_30_TDATA),
		.io_export_closureOut_31_TREADY(_peArray_31_closureIn_TREADY),
		.io_export_closureOut_31_TVALID(_Allocator_io_export_closureOut_31_TVALID),
		.io_export_closureOut_31_TDATA(_Allocator_io_export_closureOut_31_TDATA),
		.io_export_closureOut_32_TREADY(_peArray_32_closureIn_TREADY),
		.io_export_closureOut_32_TVALID(_Allocator_io_export_closureOut_32_TVALID),
		.io_export_closureOut_32_TDATA(_Allocator_io_export_closureOut_32_TDATA),
		.io_export_closureOut_33_TREADY(_peArray_33_closureIn_TREADY),
		.io_export_closureOut_33_TVALID(_Allocator_io_export_closureOut_33_TVALID),
		.io_export_closureOut_33_TDATA(_Allocator_io_export_closureOut_33_TDATA),
		.io_export_closureOut_34_TREADY(_peArray_34_closureIn_TREADY),
		.io_export_closureOut_34_TVALID(_Allocator_io_export_closureOut_34_TVALID),
		.io_export_closureOut_34_TDATA(_Allocator_io_export_closureOut_34_TDATA),
		.io_export_closureOut_35_TREADY(_peArray_35_closureIn_TREADY),
		.io_export_closureOut_35_TVALID(_Allocator_io_export_closureOut_35_TVALID),
		.io_export_closureOut_35_TDATA(_Allocator_io_export_closureOut_35_TDATA),
		.io_export_closureOut_36_TREADY(_peArray_36_closureIn_TREADY),
		.io_export_closureOut_36_TVALID(_Allocator_io_export_closureOut_36_TVALID),
		.io_export_closureOut_36_TDATA(_Allocator_io_export_closureOut_36_TDATA),
		.io_export_closureOut_37_TREADY(_peArray_37_closureIn_TREADY),
		.io_export_closureOut_37_TVALID(_Allocator_io_export_closureOut_37_TVALID),
		.io_export_closureOut_37_TDATA(_Allocator_io_export_closureOut_37_TDATA),
		.io_export_closureOut_38_TREADY(_peArray_38_closureIn_TREADY),
		.io_export_closureOut_38_TVALID(_Allocator_io_export_closureOut_38_TVALID),
		.io_export_closureOut_38_TDATA(_Allocator_io_export_closureOut_38_TDATA),
		.io_export_closureOut_39_TREADY(_peArray_39_closureIn_TREADY),
		.io_export_closureOut_39_TVALID(_Allocator_io_export_closureOut_39_TVALID),
		.io_export_closureOut_39_TDATA(_Allocator_io_export_closureOut_39_TDATA),
		.io_export_closureOut_40_TREADY(_peArray_40_closureIn_TREADY),
		.io_export_closureOut_40_TVALID(_Allocator_io_export_closureOut_40_TVALID),
		.io_export_closureOut_40_TDATA(_Allocator_io_export_closureOut_40_TDATA),
		.io_export_closureOut_41_TREADY(_peArray_41_closureIn_TREADY),
		.io_export_closureOut_41_TVALID(_Allocator_io_export_closureOut_41_TVALID),
		.io_export_closureOut_41_TDATA(_Allocator_io_export_closureOut_41_TDATA),
		.io_export_closureOut_42_TREADY(_peArray_42_closureIn_TREADY),
		.io_export_closureOut_42_TVALID(_Allocator_io_export_closureOut_42_TVALID),
		.io_export_closureOut_42_TDATA(_Allocator_io_export_closureOut_42_TDATA),
		.io_export_closureOut_43_TREADY(_peArray_43_closureIn_TREADY),
		.io_export_closureOut_43_TVALID(_Allocator_io_export_closureOut_43_TVALID),
		.io_export_closureOut_43_TDATA(_Allocator_io_export_closureOut_43_TDATA),
		.io_export_closureOut_44_TREADY(_peArray_44_closureIn_TREADY),
		.io_export_closureOut_44_TVALID(_Allocator_io_export_closureOut_44_TVALID),
		.io_export_closureOut_44_TDATA(_Allocator_io_export_closureOut_44_TDATA),
		.io_export_closureOut_45_TREADY(_peArray_45_closureIn_TREADY),
		.io_export_closureOut_45_TVALID(_Allocator_io_export_closureOut_45_TVALID),
		.io_export_closureOut_45_TDATA(_Allocator_io_export_closureOut_45_TDATA),
		.io_export_closureOut_46_TREADY(_peArray_46_closureIn_TREADY),
		.io_export_closureOut_46_TVALID(_Allocator_io_export_closureOut_46_TVALID),
		.io_export_closureOut_46_TDATA(_Allocator_io_export_closureOut_46_TDATA),
		.io_export_closureOut_47_TREADY(_peArray_47_closureIn_TREADY),
		.io_export_closureOut_47_TVALID(_Allocator_io_export_closureOut_47_TVALID),
		.io_export_closureOut_47_TDATA(_Allocator_io_export_closureOut_47_TDATA),
		.io_export_closureOut_48_TREADY(_peArray_48_closureIn_TREADY),
		.io_export_closureOut_48_TVALID(_Allocator_io_export_closureOut_48_TVALID),
		.io_export_closureOut_48_TDATA(_Allocator_io_export_closureOut_48_TDATA),
		.io_export_closureOut_49_TREADY(_peArray_49_closureIn_TREADY),
		.io_export_closureOut_49_TVALID(_Allocator_io_export_closureOut_49_TVALID),
		.io_export_closureOut_49_TDATA(_Allocator_io_export_closureOut_49_TDATA),
		.io_export_closureOut_50_TREADY(_peArray_50_closureIn_TREADY),
		.io_export_closureOut_50_TVALID(_Allocator_io_export_closureOut_50_TVALID),
		.io_export_closureOut_50_TDATA(_Allocator_io_export_closureOut_50_TDATA),
		.io_export_closureOut_51_TREADY(_peArray_51_closureIn_TREADY),
		.io_export_closureOut_51_TVALID(_Allocator_io_export_closureOut_51_TVALID),
		.io_export_closureOut_51_TDATA(_Allocator_io_export_closureOut_51_TDATA),
		.io_export_closureOut_52_TREADY(_peArray_52_closureIn_TREADY),
		.io_export_closureOut_52_TVALID(_Allocator_io_export_closureOut_52_TVALID),
		.io_export_closureOut_52_TDATA(_Allocator_io_export_closureOut_52_TDATA),
		.io_export_closureOut_53_TREADY(_peArray_53_closureIn_TREADY),
		.io_export_closureOut_53_TVALID(_Allocator_io_export_closureOut_53_TVALID),
		.io_export_closureOut_53_TDATA(_Allocator_io_export_closureOut_53_TDATA),
		.io_export_closureOut_54_TREADY(_peArray_54_closureIn_TREADY),
		.io_export_closureOut_54_TVALID(_Allocator_io_export_closureOut_54_TVALID),
		.io_export_closureOut_54_TDATA(_Allocator_io_export_closureOut_54_TDATA),
		.io_export_closureOut_55_TREADY(_peArray_55_closureIn_TREADY),
		.io_export_closureOut_55_TVALID(_Allocator_io_export_closureOut_55_TVALID),
		.io_export_closureOut_55_TDATA(_Allocator_io_export_closureOut_55_TDATA),
		.io_export_closureOut_56_TREADY(_peArray_56_closureIn_TREADY),
		.io_export_closureOut_56_TVALID(_Allocator_io_export_closureOut_56_TVALID),
		.io_export_closureOut_56_TDATA(_Allocator_io_export_closureOut_56_TDATA),
		.io_export_closureOut_57_TREADY(_peArray_57_closureIn_TREADY),
		.io_export_closureOut_57_TVALID(_Allocator_io_export_closureOut_57_TVALID),
		.io_export_closureOut_57_TDATA(_Allocator_io_export_closureOut_57_TDATA),
		.io_export_closureOut_58_TREADY(_peArray_58_closureIn_TREADY),
		.io_export_closureOut_58_TVALID(_Allocator_io_export_closureOut_58_TVALID),
		.io_export_closureOut_58_TDATA(_Allocator_io_export_closureOut_58_TDATA),
		.io_export_closureOut_59_TREADY(_peArray_59_closureIn_TREADY),
		.io_export_closureOut_59_TVALID(_Allocator_io_export_closureOut_59_TVALID),
		.io_export_closureOut_59_TDATA(_Allocator_io_export_closureOut_59_TDATA),
		.io_export_closureOut_60_TREADY(_peArray_60_closureIn_TREADY),
		.io_export_closureOut_60_TVALID(_Allocator_io_export_closureOut_60_TVALID),
		.io_export_closureOut_60_TDATA(_Allocator_io_export_closureOut_60_TDATA),
		.io_export_closureOut_61_TREADY(_peArray_61_closureIn_TREADY),
		.io_export_closureOut_61_TVALID(_Allocator_io_export_closureOut_61_TVALID),
		.io_export_closureOut_61_TDATA(_Allocator_io_export_closureOut_61_TDATA),
		.io_export_closureOut_62_TREADY(_peArray_62_closureIn_TREADY),
		.io_export_closureOut_62_TVALID(_Allocator_io_export_closureOut_62_TVALID),
		.io_export_closureOut_62_TDATA(_Allocator_io_export_closureOut_62_TDATA),
		.io_export_closureOut_63_TREADY(_peArray_63_closureIn_TREADY),
		.io_export_closureOut_63_TVALID(_Allocator_io_export_closureOut_63_TVALID),
		.io_export_closureOut_63_TDATA(_Allocator_io_export_closureOut_63_TDATA),
		.io_internal_vcas_axi_full_0_ar_ready(sum_closureAllocatorAXI_0_ARREADY),
		.io_internal_vcas_axi_full_0_ar_valid(sum_closureAllocatorAXI_0_ARVALID),
		.io_internal_vcas_axi_full_0_ar_bits_id(sum_closureAllocatorAXI_0_ARID),
		.io_internal_vcas_axi_full_0_ar_bits_addr(sum_closureAllocatorAXI_0_ARADDR),
		.io_internal_vcas_axi_full_0_ar_bits_len(sum_closureAllocatorAXI_0_ARLEN),
		.io_internal_vcas_axi_full_0_ar_bits_size(sum_closureAllocatorAXI_0_ARSIZE),
		.io_internal_vcas_axi_full_0_ar_bits_burst(sum_closureAllocatorAXI_0_ARBURST),
		.io_internal_vcas_axi_full_0_ar_bits_lock(sum_closureAllocatorAXI_0_ARLOCK),
		.io_internal_vcas_axi_full_0_ar_bits_cache(sum_closureAllocatorAXI_0_ARCACHE),
		.io_internal_vcas_axi_full_0_ar_bits_prot(sum_closureAllocatorAXI_0_ARPROT),
		.io_internal_vcas_axi_full_0_ar_bits_qos(sum_closureAllocatorAXI_0_ARQOS),
		.io_internal_vcas_axi_full_0_ar_bits_region(sum_closureAllocatorAXI_0_ARREGION),
		.io_internal_vcas_axi_full_0_r_ready(sum_closureAllocatorAXI_0_RREADY),
		.io_internal_vcas_axi_full_0_r_valid(sum_closureAllocatorAXI_0_RVALID),
		.io_internal_vcas_axi_full_0_r_bits_id(sum_closureAllocatorAXI_0_RID),
		.io_internal_vcas_axi_full_0_r_bits_data(sum_closureAllocatorAXI_0_RDATA),
		.io_internal_vcas_axi_full_0_r_bits_resp(sum_closureAllocatorAXI_0_RRESP),
		.io_internal_vcas_axi_full_0_r_bits_last(sum_closureAllocatorAXI_0_RLAST),
		.io_internal_vcas_axi_full_0_aw_ready(sum_closureAllocatorAXI_0_AWREADY),
		.io_internal_vcas_axi_full_0_aw_valid(sum_closureAllocatorAXI_0_AWVALID),
		.io_internal_vcas_axi_full_0_aw_bits_id(sum_closureAllocatorAXI_0_AWID),
		.io_internal_vcas_axi_full_0_aw_bits_addr(sum_closureAllocatorAXI_0_AWADDR),
		.io_internal_vcas_axi_full_0_aw_bits_len(sum_closureAllocatorAXI_0_AWLEN),
		.io_internal_vcas_axi_full_0_aw_bits_size(sum_closureAllocatorAXI_0_AWSIZE),
		.io_internal_vcas_axi_full_0_aw_bits_burst(sum_closureAllocatorAXI_0_AWBURST),
		.io_internal_vcas_axi_full_0_aw_bits_lock(sum_closureAllocatorAXI_0_AWLOCK),
		.io_internal_vcas_axi_full_0_aw_bits_cache(sum_closureAllocatorAXI_0_AWCACHE),
		.io_internal_vcas_axi_full_0_aw_bits_prot(sum_closureAllocatorAXI_0_AWPROT),
		.io_internal_vcas_axi_full_0_aw_bits_qos(sum_closureAllocatorAXI_0_AWQOS),
		.io_internal_vcas_axi_full_0_aw_bits_region(sum_closureAllocatorAXI_0_AWREGION),
		.io_internal_vcas_axi_full_0_w_ready(sum_closureAllocatorAXI_0_WREADY),
		.io_internal_vcas_axi_full_0_w_valid(sum_closureAllocatorAXI_0_WVALID),
		.io_internal_vcas_axi_full_0_w_bits_data(sum_closureAllocatorAXI_0_WDATA),
		.io_internal_vcas_axi_full_0_w_bits_strb(sum_closureAllocatorAXI_0_WSTRB),
		.io_internal_vcas_axi_full_0_w_bits_last(sum_closureAllocatorAXI_0_WLAST),
		.io_internal_vcas_axi_full_0_b_ready(sum_closureAllocatorAXI_0_BREADY),
		.io_internal_vcas_axi_full_0_b_valid(sum_closureAllocatorAXI_0_BVALID),
		.io_internal_vcas_axi_full_0_b_bits_id(sum_closureAllocatorAXI_0_BID),
		.io_internal_vcas_axi_full_0_b_bits_resp(sum_closureAllocatorAXI_0_BRESP),
		.io_internal_axi_mgmt_vcas_0_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_0_ar_ready),
		.io_internal_axi_mgmt_vcas_0_ar_valid(_demux_m_axil_4_ar_valid),
		.io_internal_axi_mgmt_vcas_0_ar_bits_addr(_demux_m_axil_4_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_0_ar_bits_prot(_demux_m_axil_4_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_0_r_ready(_demux_m_axil_4_r_ready),
		.io_internal_axi_mgmt_vcas_0_r_valid(_Allocator_io_internal_axi_mgmt_vcas_0_r_valid),
		.io_internal_axi_mgmt_vcas_0_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_data),
		.io_internal_axi_mgmt_vcas_0_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_resp),
		.io_internal_axi_mgmt_vcas_0_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_0_aw_ready),
		.io_internal_axi_mgmt_vcas_0_aw_valid(_demux_m_axil_4_aw_valid),
		.io_internal_axi_mgmt_vcas_0_aw_bits_addr(_demux_m_axil_4_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_0_aw_bits_prot(_demux_m_axil_4_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_0_w_ready(_Allocator_io_internal_axi_mgmt_vcas_0_w_ready),
		.io_internal_axi_mgmt_vcas_0_w_valid(_demux_m_axil_4_w_valid),
		.io_internal_axi_mgmt_vcas_0_w_bits_data(_demux_m_axil_4_w_bits_data),
		.io_internal_axi_mgmt_vcas_0_w_bits_strb(_demux_m_axil_4_w_bits_strb),
		.io_internal_axi_mgmt_vcas_0_b_ready(_demux_m_axil_4_b_ready),
		.io_internal_axi_mgmt_vcas_0_b_valid(_Allocator_io_internal_axi_mgmt_vcas_0_b_valid),
		.io_internal_axi_mgmt_vcas_0_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_b_bits_resp),
		.io_internal_axi_mgmt_vcas_1_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_1_ar_ready),
		.io_internal_axi_mgmt_vcas_1_ar_valid(_demux_m_axil_5_ar_valid),
		.io_internal_axi_mgmt_vcas_1_ar_bits_addr(_demux_m_axil_5_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_1_ar_bits_prot(_demux_m_axil_5_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_1_r_ready(_demux_m_axil_5_r_ready),
		.io_internal_axi_mgmt_vcas_1_r_valid(_Allocator_io_internal_axi_mgmt_vcas_1_r_valid),
		.io_internal_axi_mgmt_vcas_1_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_data),
		.io_internal_axi_mgmt_vcas_1_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_resp),
		.io_internal_axi_mgmt_vcas_1_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_1_aw_ready),
		.io_internal_axi_mgmt_vcas_1_aw_valid(_demux_m_axil_5_aw_valid),
		.io_internal_axi_mgmt_vcas_1_aw_bits_addr(_demux_m_axil_5_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_1_aw_bits_prot(_demux_m_axil_5_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_1_w_ready(_Allocator_io_internal_axi_mgmt_vcas_1_w_ready),
		.io_internal_axi_mgmt_vcas_1_w_valid(_demux_m_axil_5_w_valid),
		.io_internal_axi_mgmt_vcas_1_w_bits_data(_demux_m_axil_5_w_bits_data),
		.io_internal_axi_mgmt_vcas_1_w_bits_strb(_demux_m_axil_5_w_bits_strb),
		.io_internal_axi_mgmt_vcas_1_b_ready(_demux_m_axil_5_b_ready),
		.io_internal_axi_mgmt_vcas_1_b_valid(_Allocator_io_internal_axi_mgmt_vcas_1_b_valid),
		.io_internal_axi_mgmt_vcas_1_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_b_bits_resp),
		.io_internal_axi_mgmt_vcas_2_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_2_ar_ready),
		.io_internal_axi_mgmt_vcas_2_ar_valid(_demux_m_axil_6_ar_valid),
		.io_internal_axi_mgmt_vcas_2_ar_bits_addr(_demux_m_axil_6_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_2_ar_bits_prot(_demux_m_axil_6_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_2_r_ready(_demux_m_axil_6_r_ready),
		.io_internal_axi_mgmt_vcas_2_r_valid(_Allocator_io_internal_axi_mgmt_vcas_2_r_valid),
		.io_internal_axi_mgmt_vcas_2_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_data),
		.io_internal_axi_mgmt_vcas_2_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_resp),
		.io_internal_axi_mgmt_vcas_2_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_2_aw_ready),
		.io_internal_axi_mgmt_vcas_2_aw_valid(_demux_m_axil_6_aw_valid),
		.io_internal_axi_mgmt_vcas_2_aw_bits_addr(_demux_m_axil_6_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_2_aw_bits_prot(_demux_m_axil_6_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_2_w_ready(_Allocator_io_internal_axi_mgmt_vcas_2_w_ready),
		.io_internal_axi_mgmt_vcas_2_w_valid(_demux_m_axil_6_w_valid),
		.io_internal_axi_mgmt_vcas_2_w_bits_data(_demux_m_axil_6_w_bits_data),
		.io_internal_axi_mgmt_vcas_2_w_bits_strb(_demux_m_axil_6_w_bits_strb),
		.io_internal_axi_mgmt_vcas_2_b_ready(_demux_m_axil_6_b_ready),
		.io_internal_axi_mgmt_vcas_2_b_valid(_Allocator_io_internal_axi_mgmt_vcas_2_b_valid),
		.io_internal_axi_mgmt_vcas_2_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_b_bits_resp),
		.io_internal_axi_mgmt_vcas_3_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_3_ar_ready),
		.io_internal_axi_mgmt_vcas_3_ar_valid(_demux_m_axil_7_ar_valid),
		.io_internal_axi_mgmt_vcas_3_ar_bits_addr(_demux_m_axil_7_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_3_ar_bits_prot(_demux_m_axil_7_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_3_r_ready(_demux_m_axil_7_r_ready),
		.io_internal_axi_mgmt_vcas_3_r_valid(_Allocator_io_internal_axi_mgmt_vcas_3_r_valid),
		.io_internal_axi_mgmt_vcas_3_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_data),
		.io_internal_axi_mgmt_vcas_3_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_resp),
		.io_internal_axi_mgmt_vcas_3_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_3_aw_ready),
		.io_internal_axi_mgmt_vcas_3_aw_valid(_demux_m_axil_7_aw_valid),
		.io_internal_axi_mgmt_vcas_3_aw_bits_addr(_demux_m_axil_7_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_3_aw_bits_prot(_demux_m_axil_7_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_3_w_ready(_Allocator_io_internal_axi_mgmt_vcas_3_w_ready),
		.io_internal_axi_mgmt_vcas_3_w_valid(_demux_m_axil_7_w_valid),
		.io_internal_axi_mgmt_vcas_3_w_bits_data(_demux_m_axil_7_w_bits_data),
		.io_internal_axi_mgmt_vcas_3_w_bits_strb(_demux_m_axil_7_w_bits_strb),
		.io_internal_axi_mgmt_vcas_3_b_ready(_demux_m_axil_7_b_ready),
		.io_internal_axi_mgmt_vcas_3_b_valid(_Allocator_io_internal_axi_mgmt_vcas_3_b_valid),
		.io_internal_axi_mgmt_vcas_3_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_b_bits_resp)
	);
	ArgumentNotifier ArgumentNotifier(
		.clock(clock),
		.reset(reset),
		.io_export_argIn_0_TREADY(_ArgumentNotifier_io_export_argIn_0_TREADY),
		.io_export_argIn_0_TVALID(_peArray_0_argOut_TVALID),
		.io_export_argIn_0_TDATA(_peArray_0_argOut_TDATA),
		.io_export_argIn_1_TREADY(_ArgumentNotifier_io_export_argIn_1_TREADY),
		.io_export_argIn_1_TVALID(_peArray_1_argOut_TVALID),
		.io_export_argIn_1_TDATA(_peArray_1_argOut_TDATA),
		.io_export_argIn_2_TREADY(_ArgumentNotifier_io_export_argIn_2_TREADY),
		.io_export_argIn_2_TVALID(_peArray_2_argOut_TVALID),
		.io_export_argIn_2_TDATA(_peArray_2_argOut_TDATA),
		.io_export_argIn_3_TREADY(_ArgumentNotifier_io_export_argIn_3_TREADY),
		.io_export_argIn_3_TVALID(_peArray_3_argOut_TVALID),
		.io_export_argIn_3_TDATA(_peArray_3_argOut_TDATA),
		.io_export_argIn_4_TREADY(_ArgumentNotifier_io_export_argIn_4_TREADY),
		.io_export_argIn_4_TVALID(_peArray_4_argOut_TVALID),
		.io_export_argIn_4_TDATA(_peArray_4_argOut_TDATA),
		.io_export_argIn_5_TREADY(_ArgumentNotifier_io_export_argIn_5_TREADY),
		.io_export_argIn_5_TVALID(_peArray_5_argOut_TVALID),
		.io_export_argIn_5_TDATA(_peArray_5_argOut_TDATA),
		.io_export_argIn_6_TREADY(_ArgumentNotifier_io_export_argIn_6_TREADY),
		.io_export_argIn_6_TVALID(_peArray_6_argOut_TVALID),
		.io_export_argIn_6_TDATA(_peArray_6_argOut_TDATA),
		.io_export_argIn_7_TREADY(_ArgumentNotifier_io_export_argIn_7_TREADY),
		.io_export_argIn_7_TVALID(_peArray_7_argOut_TVALID),
		.io_export_argIn_7_TDATA(_peArray_7_argOut_TDATA),
		.io_export_argIn_8_TREADY(_ArgumentNotifier_io_export_argIn_8_TREADY),
		.io_export_argIn_8_TVALID(_peArray_8_argOut_TVALID),
		.io_export_argIn_8_TDATA(_peArray_8_argOut_TDATA),
		.io_export_argIn_9_TREADY(_ArgumentNotifier_io_export_argIn_9_TREADY),
		.io_export_argIn_9_TVALID(_peArray_9_argOut_TVALID),
		.io_export_argIn_9_TDATA(_peArray_9_argOut_TDATA),
		.io_export_argIn_10_TREADY(_ArgumentNotifier_io_export_argIn_10_TREADY),
		.io_export_argIn_10_TVALID(_peArray_10_argOut_TVALID),
		.io_export_argIn_10_TDATA(_peArray_10_argOut_TDATA),
		.io_export_argIn_11_TREADY(_ArgumentNotifier_io_export_argIn_11_TREADY),
		.io_export_argIn_11_TVALID(_peArray_11_argOut_TVALID),
		.io_export_argIn_11_TDATA(_peArray_11_argOut_TDATA),
		.io_export_argIn_12_TREADY(_ArgumentNotifier_io_export_argIn_12_TREADY),
		.io_export_argIn_12_TVALID(_peArray_12_argOut_TVALID),
		.io_export_argIn_12_TDATA(_peArray_12_argOut_TDATA),
		.io_export_argIn_13_TREADY(_ArgumentNotifier_io_export_argIn_13_TREADY),
		.io_export_argIn_13_TVALID(_peArray_13_argOut_TVALID),
		.io_export_argIn_13_TDATA(_peArray_13_argOut_TDATA),
		.io_export_argIn_14_TREADY(_ArgumentNotifier_io_export_argIn_14_TREADY),
		.io_export_argIn_14_TVALID(_peArray_14_argOut_TVALID),
		.io_export_argIn_14_TDATA(_peArray_14_argOut_TDATA),
		.io_export_argIn_15_TREADY(_ArgumentNotifier_io_export_argIn_15_TREADY),
		.io_export_argIn_15_TVALID(_peArray_15_argOut_TVALID),
		.io_export_argIn_15_TDATA(_peArray_15_argOut_TDATA),
		.io_export_argIn_16_TREADY(_ArgumentNotifier_io_export_argIn_16_TREADY),
		.io_export_argIn_16_TVALID(_peArray_16_argOut_TVALID),
		.io_export_argIn_16_TDATA(_peArray_16_argOut_TDATA),
		.io_export_argIn_17_TREADY(_ArgumentNotifier_io_export_argIn_17_TREADY),
		.io_export_argIn_17_TVALID(_peArray_17_argOut_TVALID),
		.io_export_argIn_17_TDATA(_peArray_17_argOut_TDATA),
		.io_export_argIn_18_TREADY(_ArgumentNotifier_io_export_argIn_18_TREADY),
		.io_export_argIn_18_TVALID(_peArray_18_argOut_TVALID),
		.io_export_argIn_18_TDATA(_peArray_18_argOut_TDATA),
		.io_export_argIn_19_TREADY(_ArgumentNotifier_io_export_argIn_19_TREADY),
		.io_export_argIn_19_TVALID(_peArray_19_argOut_TVALID),
		.io_export_argIn_19_TDATA(_peArray_19_argOut_TDATA),
		.io_export_argIn_20_TREADY(_ArgumentNotifier_io_export_argIn_20_TREADY),
		.io_export_argIn_20_TVALID(_peArray_20_argOut_TVALID),
		.io_export_argIn_20_TDATA(_peArray_20_argOut_TDATA),
		.io_export_argIn_21_TREADY(_ArgumentNotifier_io_export_argIn_21_TREADY),
		.io_export_argIn_21_TVALID(_peArray_21_argOut_TVALID),
		.io_export_argIn_21_TDATA(_peArray_21_argOut_TDATA),
		.io_export_argIn_22_TREADY(_ArgumentNotifier_io_export_argIn_22_TREADY),
		.io_export_argIn_22_TVALID(_peArray_22_argOut_TVALID),
		.io_export_argIn_22_TDATA(_peArray_22_argOut_TDATA),
		.io_export_argIn_23_TREADY(_ArgumentNotifier_io_export_argIn_23_TREADY),
		.io_export_argIn_23_TVALID(_peArray_23_argOut_TVALID),
		.io_export_argIn_23_TDATA(_peArray_23_argOut_TDATA),
		.io_export_argIn_24_TREADY(_ArgumentNotifier_io_export_argIn_24_TREADY),
		.io_export_argIn_24_TVALID(_peArray_24_argOut_TVALID),
		.io_export_argIn_24_TDATA(_peArray_24_argOut_TDATA),
		.io_export_argIn_25_TREADY(_ArgumentNotifier_io_export_argIn_25_TREADY),
		.io_export_argIn_25_TVALID(_peArray_25_argOut_TVALID),
		.io_export_argIn_25_TDATA(_peArray_25_argOut_TDATA),
		.io_export_argIn_26_TREADY(_ArgumentNotifier_io_export_argIn_26_TREADY),
		.io_export_argIn_26_TVALID(_peArray_26_argOut_TVALID),
		.io_export_argIn_26_TDATA(_peArray_26_argOut_TDATA),
		.io_export_argIn_27_TREADY(_ArgumentNotifier_io_export_argIn_27_TREADY),
		.io_export_argIn_27_TVALID(_peArray_27_argOut_TVALID),
		.io_export_argIn_27_TDATA(_peArray_27_argOut_TDATA),
		.io_export_argIn_28_TREADY(_ArgumentNotifier_io_export_argIn_28_TREADY),
		.io_export_argIn_28_TVALID(_peArray_28_argOut_TVALID),
		.io_export_argIn_28_TDATA(_peArray_28_argOut_TDATA),
		.io_export_argIn_29_TREADY(_ArgumentNotifier_io_export_argIn_29_TREADY),
		.io_export_argIn_29_TVALID(_peArray_29_argOut_TVALID),
		.io_export_argIn_29_TDATA(_peArray_29_argOut_TDATA),
		.io_export_argIn_30_TREADY(_ArgumentNotifier_io_export_argIn_30_TREADY),
		.io_export_argIn_30_TVALID(_peArray_30_argOut_TVALID),
		.io_export_argIn_30_TDATA(_peArray_30_argOut_TDATA),
		.io_export_argIn_31_TREADY(_ArgumentNotifier_io_export_argIn_31_TREADY),
		.io_export_argIn_31_TVALID(_peArray_31_argOut_TVALID),
		.io_export_argIn_31_TDATA(_peArray_31_argOut_TDATA),
		.io_export_argIn_32_TREADY(_ArgumentNotifier_io_export_argIn_32_TREADY),
		.io_export_argIn_32_TVALID(_peArray_32_argOut_TVALID),
		.io_export_argIn_32_TDATA(_peArray_32_argOut_TDATA),
		.io_export_argIn_33_TREADY(_ArgumentNotifier_io_export_argIn_33_TREADY),
		.io_export_argIn_33_TVALID(_peArray_33_argOut_TVALID),
		.io_export_argIn_33_TDATA(_peArray_33_argOut_TDATA),
		.io_export_argIn_34_TREADY(_ArgumentNotifier_io_export_argIn_34_TREADY),
		.io_export_argIn_34_TVALID(_peArray_34_argOut_TVALID),
		.io_export_argIn_34_TDATA(_peArray_34_argOut_TDATA),
		.io_export_argIn_35_TREADY(_ArgumentNotifier_io_export_argIn_35_TREADY),
		.io_export_argIn_35_TVALID(_peArray_35_argOut_TVALID),
		.io_export_argIn_35_TDATA(_peArray_35_argOut_TDATA),
		.io_export_argIn_36_TREADY(_ArgumentNotifier_io_export_argIn_36_TREADY),
		.io_export_argIn_36_TVALID(_peArray_36_argOut_TVALID),
		.io_export_argIn_36_TDATA(_peArray_36_argOut_TDATA),
		.io_export_argIn_37_TREADY(_ArgumentNotifier_io_export_argIn_37_TREADY),
		.io_export_argIn_37_TVALID(_peArray_37_argOut_TVALID),
		.io_export_argIn_37_TDATA(_peArray_37_argOut_TDATA),
		.io_export_argIn_38_TREADY(_ArgumentNotifier_io_export_argIn_38_TREADY),
		.io_export_argIn_38_TVALID(_peArray_38_argOut_TVALID),
		.io_export_argIn_38_TDATA(_peArray_38_argOut_TDATA),
		.io_export_argIn_39_TREADY(_ArgumentNotifier_io_export_argIn_39_TREADY),
		.io_export_argIn_39_TVALID(_peArray_39_argOut_TVALID),
		.io_export_argIn_39_TDATA(_peArray_39_argOut_TDATA),
		.io_export_argIn_40_TREADY(_ArgumentNotifier_io_export_argIn_40_TREADY),
		.io_export_argIn_40_TVALID(_peArray_40_argOut_TVALID),
		.io_export_argIn_40_TDATA(_peArray_40_argOut_TDATA),
		.io_export_argIn_41_TREADY(_ArgumentNotifier_io_export_argIn_41_TREADY),
		.io_export_argIn_41_TVALID(_peArray_41_argOut_TVALID),
		.io_export_argIn_41_TDATA(_peArray_41_argOut_TDATA),
		.io_export_argIn_42_TREADY(_ArgumentNotifier_io_export_argIn_42_TREADY),
		.io_export_argIn_42_TVALID(_peArray_42_argOut_TVALID),
		.io_export_argIn_42_TDATA(_peArray_42_argOut_TDATA),
		.io_export_argIn_43_TREADY(_ArgumentNotifier_io_export_argIn_43_TREADY),
		.io_export_argIn_43_TVALID(_peArray_43_argOut_TVALID),
		.io_export_argIn_43_TDATA(_peArray_43_argOut_TDATA),
		.io_export_argIn_44_TREADY(_ArgumentNotifier_io_export_argIn_44_TREADY),
		.io_export_argIn_44_TVALID(_peArray_44_argOut_TVALID),
		.io_export_argIn_44_TDATA(_peArray_44_argOut_TDATA),
		.io_export_argIn_45_TREADY(_ArgumentNotifier_io_export_argIn_45_TREADY),
		.io_export_argIn_45_TVALID(_peArray_45_argOut_TVALID),
		.io_export_argIn_45_TDATA(_peArray_45_argOut_TDATA),
		.io_export_argIn_46_TREADY(_ArgumentNotifier_io_export_argIn_46_TREADY),
		.io_export_argIn_46_TVALID(_peArray_46_argOut_TVALID),
		.io_export_argIn_46_TDATA(_peArray_46_argOut_TDATA),
		.io_export_argIn_47_TREADY(_ArgumentNotifier_io_export_argIn_47_TREADY),
		.io_export_argIn_47_TVALID(_peArray_47_argOut_TVALID),
		.io_export_argIn_47_TDATA(_peArray_47_argOut_TDATA),
		.io_export_argIn_48_TREADY(_ArgumentNotifier_io_export_argIn_48_TREADY),
		.io_export_argIn_48_TVALID(_peArray_48_argOut_TVALID),
		.io_export_argIn_48_TDATA(_peArray_48_argOut_TDATA),
		.io_export_argIn_49_TREADY(_ArgumentNotifier_io_export_argIn_49_TREADY),
		.io_export_argIn_49_TVALID(_peArray_49_argOut_TVALID),
		.io_export_argIn_49_TDATA(_peArray_49_argOut_TDATA),
		.io_export_argIn_50_TREADY(_ArgumentNotifier_io_export_argIn_50_TREADY),
		.io_export_argIn_50_TVALID(_peArray_50_argOut_TVALID),
		.io_export_argIn_50_TDATA(_peArray_50_argOut_TDATA),
		.io_export_argIn_51_TREADY(_ArgumentNotifier_io_export_argIn_51_TREADY),
		.io_export_argIn_51_TVALID(_peArray_51_argOut_TVALID),
		.io_export_argIn_51_TDATA(_peArray_51_argOut_TDATA),
		.io_export_argIn_52_TREADY(_ArgumentNotifier_io_export_argIn_52_TREADY),
		.io_export_argIn_52_TVALID(_peArray_52_argOut_TVALID),
		.io_export_argIn_52_TDATA(_peArray_52_argOut_TDATA),
		.io_export_argIn_53_TREADY(_ArgumentNotifier_io_export_argIn_53_TREADY),
		.io_export_argIn_53_TVALID(_peArray_53_argOut_TVALID),
		.io_export_argIn_53_TDATA(_peArray_53_argOut_TDATA),
		.io_export_argIn_54_TREADY(_ArgumentNotifier_io_export_argIn_54_TREADY),
		.io_export_argIn_54_TVALID(_peArray_54_argOut_TVALID),
		.io_export_argIn_54_TDATA(_peArray_54_argOut_TDATA),
		.io_export_argIn_55_TREADY(_ArgumentNotifier_io_export_argIn_55_TREADY),
		.io_export_argIn_55_TVALID(_peArray_55_argOut_TVALID),
		.io_export_argIn_55_TDATA(_peArray_55_argOut_TDATA),
		.io_export_argIn_56_TREADY(_ArgumentNotifier_io_export_argIn_56_TREADY),
		.io_export_argIn_56_TVALID(_peArray_56_argOut_TVALID),
		.io_export_argIn_56_TDATA(_peArray_56_argOut_TDATA),
		.io_export_argIn_57_TREADY(_ArgumentNotifier_io_export_argIn_57_TREADY),
		.io_export_argIn_57_TVALID(_peArray_57_argOut_TVALID),
		.io_export_argIn_57_TDATA(_peArray_57_argOut_TDATA),
		.io_export_argIn_58_TREADY(_ArgumentNotifier_io_export_argIn_58_TREADY),
		.io_export_argIn_58_TVALID(_peArray_58_argOut_TVALID),
		.io_export_argIn_58_TDATA(_peArray_58_argOut_TDATA),
		.io_export_argIn_59_TREADY(_ArgumentNotifier_io_export_argIn_59_TREADY),
		.io_export_argIn_59_TVALID(_peArray_59_argOut_TVALID),
		.io_export_argIn_59_TDATA(_peArray_59_argOut_TDATA),
		.io_export_argIn_60_TREADY(_ArgumentNotifier_io_export_argIn_60_TREADY),
		.io_export_argIn_60_TVALID(_peArray_60_argOut_TVALID),
		.io_export_argIn_60_TDATA(_peArray_60_argOut_TDATA),
		.io_export_argIn_61_TREADY(_ArgumentNotifier_io_export_argIn_61_TREADY),
		.io_export_argIn_61_TVALID(_peArray_61_argOut_TVALID),
		.io_export_argIn_61_TDATA(_peArray_61_argOut_TDATA),
		.io_export_argIn_62_TREADY(_ArgumentNotifier_io_export_argIn_62_TREADY),
		.io_export_argIn_62_TVALID(_peArray_62_argOut_TVALID),
		.io_export_argIn_62_TDATA(_peArray_62_argOut_TDATA),
		.io_export_argIn_63_TREADY(_ArgumentNotifier_io_export_argIn_63_TREADY),
		.io_export_argIn_63_TVALID(_peArray_63_argOut_TVALID),
		.io_export_argIn_63_TDATA(_peArray_63_argOut_TDATA),
		.io_export_argIn_64_TREADY(_ArgumentNotifier_io_export_argIn_64_TREADY),
		.io_export_argIn_64_TVALID(_peArray_0_1_argOut_TVALID),
		.io_export_argIn_64_TDATA(_peArray_0_1_argOut_TDATA),
		.io_export_argIn_65_TREADY(_ArgumentNotifier_io_export_argIn_65_TREADY),
		.io_export_argIn_65_TVALID(_peArray_1_1_argOut_TVALID),
		.io_export_argIn_65_TDATA(_peArray_1_1_argOut_TDATA),
		.io_export_argIn_66_TREADY(_ArgumentNotifier_io_export_argIn_66_TREADY),
		.io_export_argIn_66_TVALID(_peArray_2_1_argOut_TVALID),
		.io_export_argIn_66_TDATA(_peArray_2_1_argOut_TDATA),
		.io_export_argIn_67_TREADY(_ArgumentNotifier_io_export_argIn_67_TREADY),
		.io_export_argIn_67_TVALID(_peArray_3_1_argOut_TVALID),
		.io_export_argIn_67_TDATA(_peArray_3_1_argOut_TDATA),
		.io_export_argIn_68_TREADY(_ArgumentNotifier_io_export_argIn_68_TREADY),
		.io_export_argIn_68_TVALID(_peArray_4_1_argOut_TVALID),
		.io_export_argIn_68_TDATA(_peArray_4_1_argOut_TDATA),
		.io_export_argIn_69_TREADY(_ArgumentNotifier_io_export_argIn_69_TREADY),
		.io_export_argIn_69_TVALID(_peArray_5_1_argOut_TVALID),
		.io_export_argIn_69_TDATA(_peArray_5_1_argOut_TDATA),
		.io_export_argIn_70_TREADY(_ArgumentNotifier_io_export_argIn_70_TREADY),
		.io_export_argIn_70_TVALID(_peArray_6_1_argOut_TVALID),
		.io_export_argIn_70_TDATA(_peArray_6_1_argOut_TDATA),
		.io_export_argIn_71_TREADY(_ArgumentNotifier_io_export_argIn_71_TREADY),
		.io_export_argIn_71_TVALID(_peArray_7_1_argOut_TVALID),
		.io_export_argIn_71_TDATA(_peArray_7_1_argOut_TDATA),
		.io_export_argIn_72_TREADY(_ArgumentNotifier_io_export_argIn_72_TREADY),
		.io_export_argIn_72_TVALID(_peArray_8_1_argOut_TVALID),
		.io_export_argIn_72_TDATA(_peArray_8_1_argOut_TDATA),
		.io_export_argIn_73_TREADY(_ArgumentNotifier_io_export_argIn_73_TREADY),
		.io_export_argIn_73_TVALID(_peArray_9_1_argOut_TVALID),
		.io_export_argIn_73_TDATA(_peArray_9_1_argOut_TDATA),
		.io_export_argIn_74_TREADY(_ArgumentNotifier_io_export_argIn_74_TREADY),
		.io_export_argIn_74_TVALID(_peArray_10_1_argOut_TVALID),
		.io_export_argIn_74_TDATA(_peArray_10_1_argOut_TDATA),
		.io_export_argIn_75_TREADY(_ArgumentNotifier_io_export_argIn_75_TREADY),
		.io_export_argIn_75_TVALID(_peArray_11_1_argOut_TVALID),
		.io_export_argIn_75_TDATA(_peArray_11_1_argOut_TDATA),
		.io_export_argIn_76_TREADY(_ArgumentNotifier_io_export_argIn_76_TREADY),
		.io_export_argIn_76_TVALID(_peArray_12_1_argOut_TVALID),
		.io_export_argIn_76_TDATA(_peArray_12_1_argOut_TDATA),
		.io_export_argIn_77_TREADY(_ArgumentNotifier_io_export_argIn_77_TREADY),
		.io_export_argIn_77_TVALID(_peArray_13_1_argOut_TVALID),
		.io_export_argIn_77_TDATA(_peArray_13_1_argOut_TDATA),
		.io_export_argIn_78_TREADY(_ArgumentNotifier_io_export_argIn_78_TREADY),
		.io_export_argIn_78_TVALID(_peArray_14_1_argOut_TVALID),
		.io_export_argIn_78_TDATA(_peArray_14_1_argOut_TDATA),
		.io_export_argIn_79_TREADY(_ArgumentNotifier_io_export_argIn_79_TREADY),
		.io_export_argIn_79_TVALID(_peArray_15_1_argOut_TVALID),
		.io_export_argIn_79_TDATA(_peArray_15_1_argOut_TDATA),
		.io_export_argIn_80_TREADY(_ArgumentNotifier_io_export_argIn_80_TREADY),
		.io_export_argIn_80_TVALID(_peArray_16_1_argOut_TVALID),
		.io_export_argIn_80_TDATA(_peArray_16_1_argOut_TDATA),
		.io_export_argIn_81_TREADY(_ArgumentNotifier_io_export_argIn_81_TREADY),
		.io_export_argIn_81_TVALID(_peArray_17_1_argOut_TVALID),
		.io_export_argIn_81_TDATA(_peArray_17_1_argOut_TDATA),
		.io_export_argIn_82_TREADY(_ArgumentNotifier_io_export_argIn_82_TREADY),
		.io_export_argIn_82_TVALID(_peArray_18_1_argOut_TVALID),
		.io_export_argIn_82_TDATA(_peArray_18_1_argOut_TDATA),
		.io_export_argIn_83_TREADY(_ArgumentNotifier_io_export_argIn_83_TREADY),
		.io_export_argIn_83_TVALID(_peArray_19_1_argOut_TVALID),
		.io_export_argIn_83_TDATA(_peArray_19_1_argOut_TDATA),
		.io_export_argIn_84_TREADY(_ArgumentNotifier_io_export_argIn_84_TREADY),
		.io_export_argIn_84_TVALID(_peArray_20_1_argOut_TVALID),
		.io_export_argIn_84_TDATA(_peArray_20_1_argOut_TDATA),
		.io_export_argIn_85_TREADY(_ArgumentNotifier_io_export_argIn_85_TREADY),
		.io_export_argIn_85_TVALID(_peArray_21_1_argOut_TVALID),
		.io_export_argIn_85_TDATA(_peArray_21_1_argOut_TDATA),
		.io_export_argIn_86_TREADY(_ArgumentNotifier_io_export_argIn_86_TREADY),
		.io_export_argIn_86_TVALID(_peArray_22_1_argOut_TVALID),
		.io_export_argIn_86_TDATA(_peArray_22_1_argOut_TDATA),
		.io_export_argIn_87_TREADY(_ArgumentNotifier_io_export_argIn_87_TREADY),
		.io_export_argIn_87_TVALID(_peArray_23_1_argOut_TVALID),
		.io_export_argIn_87_TDATA(_peArray_23_1_argOut_TDATA),
		.io_export_argIn_88_TREADY(_ArgumentNotifier_io_export_argIn_88_TREADY),
		.io_export_argIn_88_TVALID(_peArray_24_1_argOut_TVALID),
		.io_export_argIn_88_TDATA(_peArray_24_1_argOut_TDATA),
		.io_export_argIn_89_TREADY(_ArgumentNotifier_io_export_argIn_89_TREADY),
		.io_export_argIn_89_TVALID(_peArray_25_1_argOut_TVALID),
		.io_export_argIn_89_TDATA(_peArray_25_1_argOut_TDATA),
		.io_export_argIn_90_TREADY(_ArgumentNotifier_io_export_argIn_90_TREADY),
		.io_export_argIn_90_TVALID(_peArray_26_1_argOut_TVALID),
		.io_export_argIn_90_TDATA(_peArray_26_1_argOut_TDATA),
		.io_export_argIn_91_TREADY(_ArgumentNotifier_io_export_argIn_91_TREADY),
		.io_export_argIn_91_TVALID(_peArray_27_1_argOut_TVALID),
		.io_export_argIn_91_TDATA(_peArray_27_1_argOut_TDATA),
		.io_export_argIn_92_TREADY(_ArgumentNotifier_io_export_argIn_92_TREADY),
		.io_export_argIn_92_TVALID(_peArray_28_1_argOut_TVALID),
		.io_export_argIn_92_TDATA(_peArray_28_1_argOut_TDATA),
		.io_export_argIn_93_TREADY(_ArgumentNotifier_io_export_argIn_93_TREADY),
		.io_export_argIn_93_TVALID(_peArray_29_1_argOut_TVALID),
		.io_export_argIn_93_TDATA(_peArray_29_1_argOut_TDATA),
		.io_export_argIn_94_TREADY(_ArgumentNotifier_io_export_argIn_94_TREADY),
		.io_export_argIn_94_TVALID(_peArray_30_1_argOut_TVALID),
		.io_export_argIn_94_TDATA(_peArray_30_1_argOut_TDATA),
		.io_export_argIn_95_TREADY(_ArgumentNotifier_io_export_argIn_95_TREADY),
		.io_export_argIn_95_TVALID(_peArray_31_1_argOut_TVALID),
		.io_export_argIn_95_TDATA(_peArray_31_1_argOut_TDATA),
		.io_export_argIn_96_TREADY(_ArgumentNotifier_io_export_argIn_96_TREADY),
		.io_export_argIn_96_TVALID(_peArray_32_1_argOut_TVALID),
		.io_export_argIn_96_TDATA(_peArray_32_1_argOut_TDATA),
		.io_export_argIn_97_TREADY(_ArgumentNotifier_io_export_argIn_97_TREADY),
		.io_export_argIn_97_TVALID(_peArray_33_1_argOut_TVALID),
		.io_export_argIn_97_TDATA(_peArray_33_1_argOut_TDATA),
		.io_export_argIn_98_TREADY(_ArgumentNotifier_io_export_argIn_98_TREADY),
		.io_export_argIn_98_TVALID(_peArray_34_1_argOut_TVALID),
		.io_export_argIn_98_TDATA(_peArray_34_1_argOut_TDATA),
		.io_export_argIn_99_TREADY(_ArgumentNotifier_io_export_argIn_99_TREADY),
		.io_export_argIn_99_TVALID(_peArray_35_1_argOut_TVALID),
		.io_export_argIn_99_TDATA(_peArray_35_1_argOut_TDATA),
		.io_export_argIn_100_TREADY(_ArgumentNotifier_io_export_argIn_100_TREADY),
		.io_export_argIn_100_TVALID(_peArray_36_1_argOut_TVALID),
		.io_export_argIn_100_TDATA(_peArray_36_1_argOut_TDATA),
		.io_export_argIn_101_TREADY(_ArgumentNotifier_io_export_argIn_101_TREADY),
		.io_export_argIn_101_TVALID(_peArray_37_1_argOut_TVALID),
		.io_export_argIn_101_TDATA(_peArray_37_1_argOut_TDATA),
		.io_export_argIn_102_TREADY(_ArgumentNotifier_io_export_argIn_102_TREADY),
		.io_export_argIn_102_TVALID(_peArray_38_1_argOut_TVALID),
		.io_export_argIn_102_TDATA(_peArray_38_1_argOut_TDATA),
		.io_export_argIn_103_TREADY(_ArgumentNotifier_io_export_argIn_103_TREADY),
		.io_export_argIn_103_TVALID(_peArray_39_1_argOut_TVALID),
		.io_export_argIn_103_TDATA(_peArray_39_1_argOut_TDATA),
		.io_export_argIn_104_TREADY(_ArgumentNotifier_io_export_argIn_104_TREADY),
		.io_export_argIn_104_TVALID(_peArray_40_1_argOut_TVALID),
		.io_export_argIn_104_TDATA(_peArray_40_1_argOut_TDATA),
		.io_export_argIn_105_TREADY(_ArgumentNotifier_io_export_argIn_105_TREADY),
		.io_export_argIn_105_TVALID(_peArray_41_1_argOut_TVALID),
		.io_export_argIn_105_TDATA(_peArray_41_1_argOut_TDATA),
		.io_export_argIn_106_TREADY(_ArgumentNotifier_io_export_argIn_106_TREADY),
		.io_export_argIn_106_TVALID(_peArray_42_1_argOut_TVALID),
		.io_export_argIn_106_TDATA(_peArray_42_1_argOut_TDATA),
		.io_export_argIn_107_TREADY(_ArgumentNotifier_io_export_argIn_107_TREADY),
		.io_export_argIn_107_TVALID(_peArray_43_1_argOut_TVALID),
		.io_export_argIn_107_TDATA(_peArray_43_1_argOut_TDATA),
		.io_export_argIn_108_TREADY(_ArgumentNotifier_io_export_argIn_108_TREADY),
		.io_export_argIn_108_TVALID(_peArray_44_1_argOut_TVALID),
		.io_export_argIn_108_TDATA(_peArray_44_1_argOut_TDATA),
		.io_export_argIn_109_TREADY(_ArgumentNotifier_io_export_argIn_109_TREADY),
		.io_export_argIn_109_TVALID(_peArray_45_1_argOut_TVALID),
		.io_export_argIn_109_TDATA(_peArray_45_1_argOut_TDATA),
		.io_export_argIn_110_TREADY(_ArgumentNotifier_io_export_argIn_110_TREADY),
		.io_export_argIn_110_TVALID(_peArray_46_1_argOut_TVALID),
		.io_export_argIn_110_TDATA(_peArray_46_1_argOut_TDATA),
		.io_export_argIn_111_TREADY(_ArgumentNotifier_io_export_argIn_111_TREADY),
		.io_export_argIn_111_TVALID(_peArray_47_1_argOut_TVALID),
		.io_export_argIn_111_TDATA(_peArray_47_1_argOut_TDATA),
		.io_export_argIn_112_TREADY(_ArgumentNotifier_io_export_argIn_112_TREADY),
		.io_export_argIn_112_TVALID(_peArray_48_1_argOut_TVALID),
		.io_export_argIn_112_TDATA(_peArray_48_1_argOut_TDATA),
		.io_export_argIn_113_TREADY(_ArgumentNotifier_io_export_argIn_113_TREADY),
		.io_export_argIn_113_TVALID(_peArray_49_1_argOut_TVALID),
		.io_export_argIn_113_TDATA(_peArray_49_1_argOut_TDATA),
		.io_export_argIn_114_TREADY(_ArgumentNotifier_io_export_argIn_114_TREADY),
		.io_export_argIn_114_TVALID(_peArray_50_1_argOut_TVALID),
		.io_export_argIn_114_TDATA(_peArray_50_1_argOut_TDATA),
		.io_export_argIn_115_TREADY(_ArgumentNotifier_io_export_argIn_115_TREADY),
		.io_export_argIn_115_TVALID(_peArray_51_1_argOut_TVALID),
		.io_export_argIn_115_TDATA(_peArray_51_1_argOut_TDATA),
		.io_export_argIn_116_TREADY(_ArgumentNotifier_io_export_argIn_116_TREADY),
		.io_export_argIn_116_TVALID(_peArray_52_1_argOut_TVALID),
		.io_export_argIn_116_TDATA(_peArray_52_1_argOut_TDATA),
		.io_export_argIn_117_TREADY(_ArgumentNotifier_io_export_argIn_117_TREADY),
		.io_export_argIn_117_TVALID(_peArray_53_1_argOut_TVALID),
		.io_export_argIn_117_TDATA(_peArray_53_1_argOut_TDATA),
		.io_export_argIn_118_TREADY(_ArgumentNotifier_io_export_argIn_118_TREADY),
		.io_export_argIn_118_TVALID(_peArray_54_1_argOut_TVALID),
		.io_export_argIn_118_TDATA(_peArray_54_1_argOut_TDATA),
		.io_export_argIn_119_TREADY(_ArgumentNotifier_io_export_argIn_119_TREADY),
		.io_export_argIn_119_TVALID(_peArray_55_1_argOut_TVALID),
		.io_export_argIn_119_TDATA(_peArray_55_1_argOut_TDATA),
		.io_export_argIn_120_TREADY(_ArgumentNotifier_io_export_argIn_120_TREADY),
		.io_export_argIn_120_TVALID(_peArray_56_1_argOut_TVALID),
		.io_export_argIn_120_TDATA(_peArray_56_1_argOut_TDATA),
		.io_export_argIn_121_TREADY(_ArgumentNotifier_io_export_argIn_121_TREADY),
		.io_export_argIn_121_TVALID(_peArray_57_1_argOut_TVALID),
		.io_export_argIn_121_TDATA(_peArray_57_1_argOut_TDATA),
		.io_export_argIn_122_TREADY(_ArgumentNotifier_io_export_argIn_122_TREADY),
		.io_export_argIn_122_TVALID(_peArray_58_1_argOut_TVALID),
		.io_export_argIn_122_TDATA(_peArray_58_1_argOut_TDATA),
		.io_export_argIn_123_TREADY(_ArgumentNotifier_io_export_argIn_123_TREADY),
		.io_export_argIn_123_TVALID(_peArray_59_1_argOut_TVALID),
		.io_export_argIn_123_TDATA(_peArray_59_1_argOut_TDATA),
		.io_export_argIn_124_TREADY(_ArgumentNotifier_io_export_argIn_124_TREADY),
		.io_export_argIn_124_TVALID(_peArray_60_1_argOut_TVALID),
		.io_export_argIn_124_TDATA(_peArray_60_1_argOut_TDATA),
		.io_export_argIn_125_TREADY(_ArgumentNotifier_io_export_argIn_125_TREADY),
		.io_export_argIn_125_TVALID(_peArray_61_1_argOut_TVALID),
		.io_export_argIn_125_TDATA(_peArray_61_1_argOut_TDATA),
		.io_export_argIn_126_TREADY(_ArgumentNotifier_io_export_argIn_126_TREADY),
		.io_export_argIn_126_TVALID(_peArray_62_1_argOut_TVALID),
		.io_export_argIn_126_TDATA(_peArray_62_1_argOut_TDATA),
		.io_export_argIn_127_TREADY(_ArgumentNotifier_io_export_argIn_127_TREADY),
		.io_export_argIn_127_TVALID(_peArray_63_1_argOut_TVALID),
		.io_export_argIn_127_TDATA(_peArray_63_1_argOut_TDATA),
		.connStealNtw_0_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_0_ctrl_serveStealReq_valid),
		.connStealNtw_0_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_0_ctrl_serveStealReq_ready),
		.connStealNtw_0_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_0_data_qOutTask_ready),
		.connStealNtw_0_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_0_data_qOutTask_valid),
		.connStealNtw_0_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_0_data_qOutTask_bits),
		.connStealNtw_1_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_1_ctrl_serveStealReq_valid),
		.connStealNtw_1_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_1_ctrl_serveStealReq_ready),
		.connStealNtw_1_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_1_data_qOutTask_ready),
		.connStealNtw_1_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_1_data_qOutTask_valid),
		.connStealNtw_1_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_1_data_qOutTask_bits),
		.connStealNtw_2_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_2_ctrl_serveStealReq_valid),
		.connStealNtw_2_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_2_ctrl_serveStealReq_ready),
		.connStealNtw_2_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_2_data_qOutTask_ready),
		.connStealNtw_2_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_2_data_qOutTask_valid),
		.connStealNtw_2_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_2_data_qOutTask_bits),
		.connStealNtw_3_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_3_ctrl_serveStealReq_valid),
		.connStealNtw_3_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_3_ctrl_serveStealReq_ready),
		.connStealNtw_3_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_3_data_qOutTask_ready),
		.connStealNtw_3_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_3_data_qOutTask_valid),
		.connStealNtw_3_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_3_data_qOutTask_bits),
		.connStealNtw_4_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_4_ctrl_serveStealReq_valid),
		.connStealNtw_4_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_4_ctrl_serveStealReq_ready),
		.connStealNtw_4_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_4_data_qOutTask_ready),
		.connStealNtw_4_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_4_data_qOutTask_valid),
		.connStealNtw_4_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_4_data_qOutTask_bits),
		.connStealNtw_5_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_5_ctrl_serveStealReq_valid),
		.connStealNtw_5_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_5_ctrl_serveStealReq_ready),
		.connStealNtw_5_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_5_data_qOutTask_ready),
		.connStealNtw_5_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_5_data_qOutTask_valid),
		.connStealNtw_5_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_5_data_qOutTask_bits),
		.connStealNtw_6_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_6_ctrl_serveStealReq_valid),
		.connStealNtw_6_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_6_ctrl_serveStealReq_ready),
		.connStealNtw_6_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_6_data_qOutTask_ready),
		.connStealNtw_6_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_6_data_qOutTask_valid),
		.connStealNtw_6_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_6_data_qOutTask_bits),
		.connStealNtw_7_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_7_ctrl_serveStealReq_valid),
		.connStealNtw_7_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_7_ctrl_serveStealReq_ready),
		.connStealNtw_7_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_7_data_qOutTask_ready),
		.connStealNtw_7_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_7_data_qOutTask_valid),
		.connStealNtw_7_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_7_data_qOutTask_bits),
		.connStealNtw_8_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_8_ctrl_serveStealReq_valid),
		.connStealNtw_8_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_8_ctrl_serveStealReq_ready),
		.connStealNtw_8_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_8_data_qOutTask_ready),
		.connStealNtw_8_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_8_data_qOutTask_valid),
		.connStealNtw_8_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_8_data_qOutTask_bits),
		.connStealNtw_9_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_9_ctrl_serveStealReq_valid),
		.connStealNtw_9_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_9_ctrl_serveStealReq_ready),
		.connStealNtw_9_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_9_data_qOutTask_ready),
		.connStealNtw_9_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_9_data_qOutTask_valid),
		.connStealNtw_9_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_9_data_qOutTask_bits),
		.connStealNtw_10_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_10_ctrl_serveStealReq_valid),
		.connStealNtw_10_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_10_ctrl_serveStealReq_ready),
		.connStealNtw_10_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_10_data_qOutTask_ready),
		.connStealNtw_10_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_10_data_qOutTask_valid),
		.connStealNtw_10_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_10_data_qOutTask_bits),
		.connStealNtw_11_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_11_ctrl_serveStealReq_valid),
		.connStealNtw_11_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_11_ctrl_serveStealReq_ready),
		.connStealNtw_11_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_11_data_qOutTask_ready),
		.connStealNtw_11_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_11_data_qOutTask_valid),
		.connStealNtw_11_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_11_data_qOutTask_bits),
		.connStealNtw_12_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_12_ctrl_serveStealReq_valid),
		.connStealNtw_12_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_12_ctrl_serveStealReq_ready),
		.connStealNtw_12_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_12_data_qOutTask_ready),
		.connStealNtw_12_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_12_data_qOutTask_valid),
		.connStealNtw_12_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_12_data_qOutTask_bits),
		.connStealNtw_13_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_13_ctrl_serveStealReq_valid),
		.connStealNtw_13_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_13_ctrl_serveStealReq_ready),
		.connStealNtw_13_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_13_data_qOutTask_ready),
		.connStealNtw_13_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_13_data_qOutTask_valid),
		.connStealNtw_13_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_13_data_qOutTask_bits),
		.connStealNtw_14_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_14_ctrl_serveStealReq_valid),
		.connStealNtw_14_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_14_ctrl_serveStealReq_ready),
		.connStealNtw_14_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_14_data_qOutTask_ready),
		.connStealNtw_14_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_14_data_qOutTask_valid),
		.connStealNtw_14_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_14_data_qOutTask_bits),
		.connStealNtw_15_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_15_ctrl_serveStealReq_valid),
		.connStealNtw_15_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_15_ctrl_serveStealReq_ready),
		.connStealNtw_15_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_15_data_qOutTask_ready),
		.connStealNtw_15_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_15_data_qOutTask_valid),
		.connStealNtw_15_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_15_data_qOutTask_bits),
		.axi_full_argRoute_0_ar_ready(sum_argumentNotifierAXI_0_ARREADY),
		.axi_full_argRoute_0_ar_valid(sum_argumentNotifierAXI_0_ARVALID),
		.axi_full_argRoute_0_ar_bits_id(sum_argumentNotifierAXI_0_ARID),
		.axi_full_argRoute_0_ar_bits_addr(sum_argumentNotifierAXI_0_ARADDR),
		.axi_full_argRoute_0_ar_bits_len(sum_argumentNotifierAXI_0_ARLEN),
		.axi_full_argRoute_0_ar_bits_size(sum_argumentNotifierAXI_0_ARSIZE),
		.axi_full_argRoute_0_ar_bits_burst(sum_argumentNotifierAXI_0_ARBURST),
		.axi_full_argRoute_0_ar_bits_lock(sum_argumentNotifierAXI_0_ARLOCK),
		.axi_full_argRoute_0_ar_bits_cache(sum_argumentNotifierAXI_0_ARCACHE),
		.axi_full_argRoute_0_ar_bits_prot(sum_argumentNotifierAXI_0_ARPROT),
		.axi_full_argRoute_0_ar_bits_qos(sum_argumentNotifierAXI_0_ARQOS),
		.axi_full_argRoute_0_ar_bits_region(sum_argumentNotifierAXI_0_ARREGION),
		.axi_full_argRoute_0_r_ready(sum_argumentNotifierAXI_0_RREADY),
		.axi_full_argRoute_0_r_valid(sum_argumentNotifierAXI_0_RVALID),
		.axi_full_argRoute_0_r_bits_id(sum_argumentNotifierAXI_0_RID),
		.axi_full_argRoute_0_r_bits_data(sum_argumentNotifierAXI_0_RDATA),
		.axi_full_argRoute_0_r_bits_resp(sum_argumentNotifierAXI_0_RRESP),
		.axi_full_argRoute_0_r_bits_last(sum_argumentNotifierAXI_0_RLAST),
		.axi_full_argRoute_0_aw_ready(sum_argumentNotifierAXI_0_AWREADY),
		.axi_full_argRoute_0_aw_valid(sum_argumentNotifierAXI_0_AWVALID),
		.axi_full_argRoute_0_aw_bits_id(sum_argumentNotifierAXI_0_AWID),
		.axi_full_argRoute_0_aw_bits_addr(sum_argumentNotifierAXI_0_AWADDR),
		.axi_full_argRoute_0_aw_bits_len(sum_argumentNotifierAXI_0_AWLEN),
		.axi_full_argRoute_0_aw_bits_size(sum_argumentNotifierAXI_0_AWSIZE),
		.axi_full_argRoute_0_aw_bits_burst(sum_argumentNotifierAXI_0_AWBURST),
		.axi_full_argRoute_0_aw_bits_lock(sum_argumentNotifierAXI_0_AWLOCK),
		.axi_full_argRoute_0_aw_bits_cache(sum_argumentNotifierAXI_0_AWCACHE),
		.axi_full_argRoute_0_aw_bits_prot(sum_argumentNotifierAXI_0_AWPROT),
		.axi_full_argRoute_0_aw_bits_qos(sum_argumentNotifierAXI_0_AWQOS),
		.axi_full_argRoute_0_aw_bits_region(sum_argumentNotifierAXI_0_AWREGION),
		.axi_full_argRoute_0_w_ready(sum_argumentNotifierAXI_0_WREADY),
		.axi_full_argRoute_0_w_valid(sum_argumentNotifierAXI_0_WVALID),
		.axi_full_argRoute_0_w_bits_data(sum_argumentNotifierAXI_0_WDATA),
		.axi_full_argRoute_0_w_bits_strb(sum_argumentNotifierAXI_0_WSTRB),
		.axi_full_argRoute_0_w_bits_last(sum_argumentNotifierAXI_0_WLAST),
		.axi_full_argRoute_0_b_ready(sum_argumentNotifierAXI_0_BREADY),
		.axi_full_argRoute_0_b_valid(sum_argumentNotifierAXI_0_BVALID),
		.axi_full_argRoute_0_b_bits_id(sum_argumentNotifierAXI_0_BID),
		.axi_full_argRoute_0_b_bits_resp(sum_argumentNotifierAXI_0_BRESP)
	);
endmodule
