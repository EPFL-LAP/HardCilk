module ram_2x15 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [14:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [14:0] W0_data;
	reg [14:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 15'bxxxxxxxxxxxxxxx);
endmodule
module Queue2_AddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_prot,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_prot
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [11:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_prot;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [11:0] io_deq_bits_addr;
	output wire [2:0] io_deq_bits_prot;
	wire [14:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x15 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_prot, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[11:0];
	assign io_deq_bits_prot = _ram_ext_R0_data[14:12];
endmodule
module ram_2x66 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [65:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [65:0] W0_data;
	reg [65:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 66'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_ReadDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	wire [65:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x66 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_resp, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[63:0];
	assign io_deq_bits_resp = _ram_ext_R0_data[65:64];
endmodule
module ram_2x72 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [71:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [71:0] W0_data;
	reg [71:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 72'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [7:0] io_enq_bits_strb;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [7:0] io_deq_bits_strb;
	wire [71:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x72 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_strb, io_enq_bits_data})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_data = _ram_ext_R0_data[63:0];
	assign io_deq_bits_strb = _ram_ext_R0_data[71:64];
endmodule
module ram_resp_2x2 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [1:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [1:0] W0_data;
	reg [1:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 2'bxx);
endmodule
module Queue2_WriteResponseChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [1:0] io_deq_bits_resp;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_resp_2x2 ram_resp_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_resp),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_resp)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module ram_8x3 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [2:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [2:0] R0_data;
	input [2:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [2:0] W0_data;
	reg [2:0] Memory [0:7];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 3'bxxx);
endmodule
module Queue8_UInt3 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits;
	wire io_enq_ready_0;
	wire [2:0] _ram_ext_R0_data;
	reg [2:0] enq_ptr_value;
	reg [2:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire io_deq_valid_0 = io_enq_valid | ~empty;
	wire do_deq = (~empty & io_deq_ready) & io_deq_valid_0;
	wire do_enq = (~(empty & io_deq_ready) & io_enq_ready_0) & io_enq_valid;
	assign io_enq_ready_0 = io_deq_ready | ~(ptr_match & maybe_full);
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 3'h0;
			deq_ptr_value <= 3'h0;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 3'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 3'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_8x3 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = io_enq_ready_0;
	assign io_deq_valid = io_deq_valid_0;
	assign io_deq_bits = (empty ? io_enq_bits : _ram_ext_R0_data);
endmodule
module elasticDemux (
	io_source_ready,
	io_source_valid,
	io_source_bits_addr,
	io_source_bits_prot,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_addr,
	io_sinks_0_bits_prot,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_addr,
	io_sinks_1_bits_prot,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_2_bits_addr,
	io_sinks_2_bits_prot,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_3_bits_addr,
	io_sinks_3_bits_prot,
	io_sinks_4_ready,
	io_sinks_4_valid,
	io_sinks_4_bits_addr,
	io_sinks_4_bits_prot,
	io_sinks_5_ready,
	io_sinks_5_valid,
	io_sinks_5_bits_addr,
	io_sinks_5_bits_prot,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [11:0] io_source_bits_addr;
	input [2:0] io_source_bits_prot;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [11:0] io_sinks_0_bits_addr;
	output wire [2:0] io_sinks_0_bits_prot;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [11:0] io_sinks_1_bits_addr;
	output wire [2:0] io_sinks_1_bits_prot;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	output wire [11:0] io_sinks_2_bits_addr;
	output wire [2:0] io_sinks_2_bits_prot;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire [11:0] io_sinks_3_bits_addr;
	output wire [2:0] io_sinks_3_bits_prot;
	input io_sinks_4_ready;
	output wire io_sinks_4_valid;
	output wire [11:0] io_sinks_4_bits_addr;
	output wire [2:0] io_sinks_4_bits_prot;
	input io_sinks_5_ready;
	output wire io_sinks_5_valid;
	output wire [11:0] io_sinks_5_bits_addr;
	output wire [2:0] io_sinks_5_bits_prot;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [7:0] _GEN = {io_sinks_0_ready, io_sinks_0_ready, io_sinks_5_ready, io_sinks_4_ready, io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 3'h0);
	assign io_sinks_0_bits_addr = io_source_bits_addr;
	assign io_sinks_0_bits_prot = io_source_bits_prot;
	assign io_sinks_1_valid = valid & (io_select_bits == 3'h1);
	assign io_sinks_1_bits_addr = io_source_bits_addr;
	assign io_sinks_1_bits_prot = io_source_bits_prot;
	assign io_sinks_2_valid = valid & (io_select_bits == 3'h2);
	assign io_sinks_2_bits_addr = io_source_bits_addr;
	assign io_sinks_2_bits_prot = io_source_bits_prot;
	assign io_sinks_3_valid = valid & (io_select_bits == 3'h3);
	assign io_sinks_3_bits_addr = io_source_bits_addr;
	assign io_sinks_3_bits_prot = io_source_bits_prot;
	assign io_sinks_4_valid = valid & (io_select_bits == 3'h4);
	assign io_sinks_4_bits_addr = io_source_bits_addr;
	assign io_sinks_4_bits_prot = io_source_bits_prot;
	assign io_sinks_5_valid = valid & (io_select_bits == 3'h5);
	assign io_sinks_5_bits_addr = io_source_bits_addr;
	assign io_sinks_5_bits_prot = io_source_bits_prot;
	assign io_select_ready = fire;
endmodule
module elasticMux (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_data,
	io_sources_0_bits_resp,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_data,
	io_sources_1_bits_resp,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_data,
	io_sources_2_bits_resp,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_data,
	io_sources_3_bits_resp,
	io_sources_4_ready,
	io_sources_4_valid,
	io_sources_4_bits_data,
	io_sources_4_bits_resp,
	io_sources_5_ready,
	io_sources_5_valid,
	io_sources_5_bits_data,
	io_sources_5_bits_resp,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_data,
	io_sink_bits_resp,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [63:0] io_sources_0_bits_data;
	input [1:0] io_sources_0_bits_resp;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [63:0] io_sources_1_bits_data;
	input [1:0] io_sources_1_bits_resp;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [63:0] io_sources_2_bits_data;
	input [1:0] io_sources_2_bits_resp;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [63:0] io_sources_3_bits_data;
	input [1:0] io_sources_3_bits_resp;
	output wire io_sources_4_ready;
	input io_sources_4_valid;
	input [63:0] io_sources_4_bits_data;
	input [1:0] io_sources_4_bits_resp;
	output wire io_sources_5_ready;
	input io_sources_5_valid;
	input [63:0] io_sources_5_bits_data;
	input [1:0] io_sources_5_bits_resp;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [63:0] io_sink_bits_data;
	output wire [1:0] io_sink_bits_resp;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire [7:0] _GEN = {io_sources_0_valid, io_sources_0_valid, io_sources_5_valid, io_sources_4_valid, io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [511:0] _GEN_0 = {io_sources_0_bits_data, io_sources_0_bits_data, io_sources_5_bits_data, io_sources_4_bits_data, io_sources_3_bits_data, io_sources_2_bits_data, io_sources_1_bits_data, io_sources_0_bits_data};
	wire [15:0] _GEN_1 = {io_sources_0_bits_resp, io_sources_0_bits_resp, io_sources_5_bits_resp, io_sources_4_bits_resp, io_sources_3_bits_resp, io_sources_2_bits_resp, io_sources_1_bits_resp, io_sources_0_bits_resp};
	wire valid = io_select_valid & _GEN[io_select_bits];
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & (io_select_bits == 3'h0);
	assign io_sources_1_ready = fire & (io_select_bits == 3'h1);
	assign io_sources_2_ready = fire & (io_select_bits == 3'h2);
	assign io_sources_3_ready = fire & (io_select_bits == 3'h3);
	assign io_sources_4_ready = fire & (io_select_bits == 3'h4);
	assign io_sources_5_ready = fire & (io_select_bits == 3'h5);
	assign io_sink_valid = valid;
	assign io_sink_bits_data = _GEN_0[io_select_bits * 64+:64];
	assign io_sink_bits_resp = _GEN_1[io_select_bits * 2+:2];
	assign io_select_ready = fire;
endmodule
module elasticDemux_2 (
	io_source_ready,
	io_source_valid,
	io_source_bits_data,
	io_source_bits_strb,
	io_sinks_0_ready,
	io_sinks_0_valid,
	io_sinks_0_bits_data,
	io_sinks_0_bits_strb,
	io_sinks_1_ready,
	io_sinks_1_valid,
	io_sinks_1_bits_data,
	io_sinks_1_bits_strb,
	io_sinks_2_ready,
	io_sinks_2_valid,
	io_sinks_2_bits_data,
	io_sinks_2_bits_strb,
	io_sinks_3_ready,
	io_sinks_3_valid,
	io_sinks_3_bits_data,
	io_sinks_3_bits_strb,
	io_sinks_4_ready,
	io_sinks_4_valid,
	io_sinks_4_bits_data,
	io_sinks_4_bits_strb,
	io_sinks_5_ready,
	io_sinks_5_valid,
	io_sinks_5_bits_data,
	io_sinks_5_bits_strb,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_source_ready;
	input io_source_valid;
	input [63:0] io_source_bits_data;
	input [7:0] io_source_bits_strb;
	input io_sinks_0_ready;
	output wire io_sinks_0_valid;
	output wire [63:0] io_sinks_0_bits_data;
	output wire [7:0] io_sinks_0_bits_strb;
	input io_sinks_1_ready;
	output wire io_sinks_1_valid;
	output wire [63:0] io_sinks_1_bits_data;
	output wire [7:0] io_sinks_1_bits_strb;
	input io_sinks_2_ready;
	output wire io_sinks_2_valid;
	output wire [63:0] io_sinks_2_bits_data;
	output wire [7:0] io_sinks_2_bits_strb;
	input io_sinks_3_ready;
	output wire io_sinks_3_valid;
	output wire [63:0] io_sinks_3_bits_data;
	output wire [7:0] io_sinks_3_bits_strb;
	input io_sinks_4_ready;
	output wire io_sinks_4_valid;
	output wire [63:0] io_sinks_4_bits_data;
	output wire [7:0] io_sinks_4_bits_strb;
	input io_sinks_5_ready;
	output wire io_sinks_5_valid;
	output wire [63:0] io_sinks_5_bits_data;
	output wire [7:0] io_sinks_5_bits_strb;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire valid = io_select_valid & io_source_valid;
	wire [7:0] _GEN = {io_sinks_0_ready, io_sinks_0_ready, io_sinks_5_ready, io_sinks_4_ready, io_sinks_3_ready, io_sinks_2_ready, io_sinks_1_ready, io_sinks_0_ready};
	wire fire = valid & _GEN[io_select_bits];
	assign io_source_ready = fire;
	assign io_sinks_0_valid = valid & (io_select_bits == 3'h0);
	assign io_sinks_0_bits_data = io_source_bits_data;
	assign io_sinks_0_bits_strb = io_source_bits_strb;
	assign io_sinks_1_valid = valid & (io_select_bits == 3'h1);
	assign io_sinks_1_bits_data = io_source_bits_data;
	assign io_sinks_1_bits_strb = io_source_bits_strb;
	assign io_sinks_2_valid = valid & (io_select_bits == 3'h2);
	assign io_sinks_2_bits_data = io_source_bits_data;
	assign io_sinks_2_bits_strb = io_source_bits_strb;
	assign io_sinks_3_valid = valid & (io_select_bits == 3'h3);
	assign io_sinks_3_bits_data = io_source_bits_data;
	assign io_sinks_3_bits_strb = io_source_bits_strb;
	assign io_sinks_4_valid = valid & (io_select_bits == 3'h4);
	assign io_sinks_4_bits_data = io_source_bits_data;
	assign io_sinks_4_bits_strb = io_source_bits_strb;
	assign io_sinks_5_valid = valid & (io_select_bits == 3'h5);
	assign io_sinks_5_bits_data = io_source_bits_data;
	assign io_sinks_5_bits_strb = io_source_bits_strb;
	assign io_select_ready = fire;
endmodule
module elasticMux_1 (
	io_sources_0_ready,
	io_sources_0_valid,
	io_sources_0_bits_resp,
	io_sources_1_ready,
	io_sources_1_valid,
	io_sources_1_bits_resp,
	io_sources_2_ready,
	io_sources_2_valid,
	io_sources_2_bits_resp,
	io_sources_3_ready,
	io_sources_3_valid,
	io_sources_3_bits_resp,
	io_sources_4_ready,
	io_sources_4_valid,
	io_sources_4_bits_resp,
	io_sources_5_ready,
	io_sources_5_valid,
	io_sources_5_bits_resp,
	io_sink_ready,
	io_sink_valid,
	io_sink_bits_resp,
	io_select_ready,
	io_select_valid,
	io_select_bits
);
	output wire io_sources_0_ready;
	input io_sources_0_valid;
	input [1:0] io_sources_0_bits_resp;
	output wire io_sources_1_ready;
	input io_sources_1_valid;
	input [1:0] io_sources_1_bits_resp;
	output wire io_sources_2_ready;
	input io_sources_2_valid;
	input [1:0] io_sources_2_bits_resp;
	output wire io_sources_3_ready;
	input io_sources_3_valid;
	input [1:0] io_sources_3_bits_resp;
	output wire io_sources_4_ready;
	input io_sources_4_valid;
	input [1:0] io_sources_4_bits_resp;
	output wire io_sources_5_ready;
	input io_sources_5_valid;
	input [1:0] io_sources_5_bits_resp;
	input io_sink_ready;
	output wire io_sink_valid;
	output wire [1:0] io_sink_bits_resp;
	output wire io_select_ready;
	input io_select_valid;
	input [2:0] io_select_bits;
	wire [7:0] _GEN = {io_sources_0_valid, io_sources_0_valid, io_sources_5_valid, io_sources_4_valid, io_sources_3_valid, io_sources_2_valid, io_sources_1_valid, io_sources_0_valid};
	wire [15:0] _GEN_0 = {io_sources_0_bits_resp, io_sources_0_bits_resp, io_sources_5_bits_resp, io_sources_4_bits_resp, io_sources_3_bits_resp, io_sources_2_bits_resp, io_sources_1_bits_resp, io_sources_0_bits_resp};
	wire valid = io_select_valid & _GEN[io_select_bits];
	wire fire = valid & io_sink_ready;
	assign io_sources_0_ready = fire & (io_select_bits == 3'h0);
	assign io_sources_1_ready = fire & (io_select_bits == 3'h1);
	assign io_sources_2_ready = fire & (io_select_bits == 3'h2);
	assign io_sources_3_ready = fire & (io_select_bits == 3'h3);
	assign io_sources_4_ready = fire & (io_select_bits == 3'h4);
	assign io_sources_5_ready = fire & (io_select_bits == 3'h5);
	assign io_sink_valid = valid;
	assign io_sink_bits_resp = _GEN_0[io_select_bits * 2+:2];
	assign io_select_ready = fire;
endmodule
module axi4LiteDemux (
	clock,
	reset,
	s_axil_ar_ready,
	s_axil_ar_valid,
	s_axil_ar_bits_addr,
	s_axil_ar_bits_prot,
	s_axil_r_ready,
	s_axil_r_valid,
	s_axil_r_bits_data,
	s_axil_r_bits_resp,
	s_axil_aw_ready,
	s_axil_aw_valid,
	s_axil_aw_bits_addr,
	s_axil_aw_bits_prot,
	s_axil_w_ready,
	s_axil_w_valid,
	s_axil_w_bits_data,
	s_axil_w_bits_strb,
	s_axil_b_ready,
	s_axil_b_valid,
	s_axil_b_bits_resp,
	m_axil_0_ar_ready,
	m_axil_0_ar_valid,
	m_axil_0_ar_bits_addr,
	m_axil_0_ar_bits_prot,
	m_axil_0_r_ready,
	m_axil_0_r_valid,
	m_axil_0_r_bits_data,
	m_axil_0_r_bits_resp,
	m_axil_0_aw_ready,
	m_axil_0_aw_valid,
	m_axil_0_aw_bits_addr,
	m_axil_0_aw_bits_prot,
	m_axil_0_w_ready,
	m_axil_0_w_valid,
	m_axil_0_w_bits_data,
	m_axil_0_w_bits_strb,
	m_axil_0_b_ready,
	m_axil_0_b_valid,
	m_axil_0_b_bits_resp,
	m_axil_1_ar_ready,
	m_axil_1_ar_valid,
	m_axil_1_ar_bits_addr,
	m_axil_1_ar_bits_prot,
	m_axil_1_r_ready,
	m_axil_1_r_valid,
	m_axil_1_r_bits_data,
	m_axil_1_r_bits_resp,
	m_axil_1_aw_ready,
	m_axil_1_aw_valid,
	m_axil_1_aw_bits_addr,
	m_axil_1_aw_bits_prot,
	m_axil_1_w_ready,
	m_axil_1_w_valid,
	m_axil_1_w_bits_data,
	m_axil_1_w_bits_strb,
	m_axil_1_b_ready,
	m_axil_1_b_valid,
	m_axil_1_b_bits_resp,
	m_axil_2_ar_ready,
	m_axil_2_ar_valid,
	m_axil_2_ar_bits_addr,
	m_axil_2_ar_bits_prot,
	m_axil_2_r_ready,
	m_axil_2_r_valid,
	m_axil_2_r_bits_data,
	m_axil_2_r_bits_resp,
	m_axil_2_aw_ready,
	m_axil_2_aw_valid,
	m_axil_2_aw_bits_addr,
	m_axil_2_aw_bits_prot,
	m_axil_2_w_ready,
	m_axil_2_w_valid,
	m_axil_2_w_bits_data,
	m_axil_2_w_bits_strb,
	m_axil_2_b_ready,
	m_axil_2_b_valid,
	m_axil_2_b_bits_resp,
	m_axil_3_ar_ready,
	m_axil_3_ar_valid,
	m_axil_3_ar_bits_addr,
	m_axil_3_ar_bits_prot,
	m_axil_3_r_ready,
	m_axil_3_r_valid,
	m_axil_3_r_bits_data,
	m_axil_3_r_bits_resp,
	m_axil_3_aw_ready,
	m_axil_3_aw_valid,
	m_axil_3_aw_bits_addr,
	m_axil_3_aw_bits_prot,
	m_axil_3_w_ready,
	m_axil_3_w_valid,
	m_axil_3_w_bits_data,
	m_axil_3_w_bits_strb,
	m_axil_3_b_ready,
	m_axil_3_b_valid,
	m_axil_3_b_bits_resp,
	m_axil_4_ar_ready,
	m_axil_4_ar_valid,
	m_axil_4_ar_bits_addr,
	m_axil_4_ar_bits_prot,
	m_axil_4_r_ready,
	m_axil_4_r_valid,
	m_axil_4_r_bits_data,
	m_axil_4_r_bits_resp,
	m_axil_4_aw_ready,
	m_axil_4_aw_valid,
	m_axil_4_aw_bits_addr,
	m_axil_4_aw_bits_prot,
	m_axil_4_w_ready,
	m_axil_4_w_valid,
	m_axil_4_w_bits_data,
	m_axil_4_w_bits_strb,
	m_axil_4_b_ready,
	m_axil_4_b_valid,
	m_axil_4_b_bits_resp,
	m_axil_5_ar_ready,
	m_axil_5_ar_valid,
	m_axil_5_ar_bits_addr,
	m_axil_5_ar_bits_prot,
	m_axil_5_r_ready,
	m_axil_5_r_valid,
	m_axil_5_r_bits_data,
	m_axil_5_r_bits_resp,
	m_axil_5_aw_ready,
	m_axil_5_aw_valid,
	m_axil_5_aw_bits_addr,
	m_axil_5_aw_bits_prot,
	m_axil_5_w_ready,
	m_axil_5_w_valid,
	m_axil_5_w_bits_data,
	m_axil_5_w_bits_strb,
	m_axil_5_b_ready,
	m_axil_5_b_valid,
	m_axil_5_b_bits_resp
);
	input clock;
	input reset;
	output wire s_axil_ar_ready;
	input s_axil_ar_valid;
	input [11:0] s_axil_ar_bits_addr;
	input [2:0] s_axil_ar_bits_prot;
	input s_axil_r_ready;
	output wire s_axil_r_valid;
	output wire [63:0] s_axil_r_bits_data;
	output wire [1:0] s_axil_r_bits_resp;
	output wire s_axil_aw_ready;
	input s_axil_aw_valid;
	input [11:0] s_axil_aw_bits_addr;
	input [2:0] s_axil_aw_bits_prot;
	output wire s_axil_w_ready;
	input s_axil_w_valid;
	input [63:0] s_axil_w_bits_data;
	input [7:0] s_axil_w_bits_strb;
	input s_axil_b_ready;
	output wire s_axil_b_valid;
	output wire [1:0] s_axil_b_bits_resp;
	input m_axil_0_ar_ready;
	output wire m_axil_0_ar_valid;
	output wire [11:0] m_axil_0_ar_bits_addr;
	output wire [2:0] m_axil_0_ar_bits_prot;
	output wire m_axil_0_r_ready;
	input m_axil_0_r_valid;
	input [63:0] m_axil_0_r_bits_data;
	input [1:0] m_axil_0_r_bits_resp;
	input m_axil_0_aw_ready;
	output wire m_axil_0_aw_valid;
	output wire [11:0] m_axil_0_aw_bits_addr;
	output wire [2:0] m_axil_0_aw_bits_prot;
	input m_axil_0_w_ready;
	output wire m_axil_0_w_valid;
	output wire [63:0] m_axil_0_w_bits_data;
	output wire [7:0] m_axil_0_w_bits_strb;
	output wire m_axil_0_b_ready;
	input m_axil_0_b_valid;
	input [1:0] m_axil_0_b_bits_resp;
	input m_axil_1_ar_ready;
	output wire m_axil_1_ar_valid;
	output wire [11:0] m_axil_1_ar_bits_addr;
	output wire [2:0] m_axil_1_ar_bits_prot;
	output wire m_axil_1_r_ready;
	input m_axil_1_r_valid;
	input [63:0] m_axil_1_r_bits_data;
	input [1:0] m_axil_1_r_bits_resp;
	input m_axil_1_aw_ready;
	output wire m_axil_1_aw_valid;
	output wire [11:0] m_axil_1_aw_bits_addr;
	output wire [2:0] m_axil_1_aw_bits_prot;
	input m_axil_1_w_ready;
	output wire m_axil_1_w_valid;
	output wire [63:0] m_axil_1_w_bits_data;
	output wire [7:0] m_axil_1_w_bits_strb;
	output wire m_axil_1_b_ready;
	input m_axil_1_b_valid;
	input [1:0] m_axil_1_b_bits_resp;
	input m_axil_2_ar_ready;
	output wire m_axil_2_ar_valid;
	output wire [11:0] m_axil_2_ar_bits_addr;
	output wire [2:0] m_axil_2_ar_bits_prot;
	output wire m_axil_2_r_ready;
	input m_axil_2_r_valid;
	input [63:0] m_axil_2_r_bits_data;
	input [1:0] m_axil_2_r_bits_resp;
	input m_axil_2_aw_ready;
	output wire m_axil_2_aw_valid;
	output wire [11:0] m_axil_2_aw_bits_addr;
	output wire [2:0] m_axil_2_aw_bits_prot;
	input m_axil_2_w_ready;
	output wire m_axil_2_w_valid;
	output wire [63:0] m_axil_2_w_bits_data;
	output wire [7:0] m_axil_2_w_bits_strb;
	output wire m_axil_2_b_ready;
	input m_axil_2_b_valid;
	input [1:0] m_axil_2_b_bits_resp;
	input m_axil_3_ar_ready;
	output wire m_axil_3_ar_valid;
	output wire [11:0] m_axil_3_ar_bits_addr;
	output wire [2:0] m_axil_3_ar_bits_prot;
	output wire m_axil_3_r_ready;
	input m_axil_3_r_valid;
	input [63:0] m_axil_3_r_bits_data;
	input [1:0] m_axil_3_r_bits_resp;
	input m_axil_3_aw_ready;
	output wire m_axil_3_aw_valid;
	output wire [11:0] m_axil_3_aw_bits_addr;
	output wire [2:0] m_axil_3_aw_bits_prot;
	input m_axil_3_w_ready;
	output wire m_axil_3_w_valid;
	output wire [63:0] m_axil_3_w_bits_data;
	output wire [7:0] m_axil_3_w_bits_strb;
	output wire m_axil_3_b_ready;
	input m_axil_3_b_valid;
	input [1:0] m_axil_3_b_bits_resp;
	input m_axil_4_ar_ready;
	output wire m_axil_4_ar_valid;
	output wire [11:0] m_axil_4_ar_bits_addr;
	output wire [2:0] m_axil_4_ar_bits_prot;
	output wire m_axil_4_r_ready;
	input m_axil_4_r_valid;
	input [63:0] m_axil_4_r_bits_data;
	input [1:0] m_axil_4_r_bits_resp;
	input m_axil_4_aw_ready;
	output wire m_axil_4_aw_valid;
	output wire [11:0] m_axil_4_aw_bits_addr;
	output wire [2:0] m_axil_4_aw_bits_prot;
	input m_axil_4_w_ready;
	output wire m_axil_4_w_valid;
	output wire [63:0] m_axil_4_w_bits_data;
	output wire [7:0] m_axil_4_w_bits_strb;
	output wire m_axil_4_b_ready;
	input m_axil_4_b_valid;
	input [1:0] m_axil_4_b_bits_resp;
	input m_axil_5_ar_ready;
	output wire m_axil_5_ar_valid;
	output wire [11:0] m_axil_5_ar_bits_addr;
	output wire [2:0] m_axil_5_ar_bits_prot;
	output wire m_axil_5_r_ready;
	input m_axil_5_r_valid;
	input [63:0] m_axil_5_r_bits_data;
	input [1:0] m_axil_5_r_bits_resp;
	input m_axil_5_aw_ready;
	output wire m_axil_5_aw_valid;
	output wire [11:0] m_axil_5_aw_bits_addr;
	output wire [2:0] m_axil_5_aw_bits_prot;
	input m_axil_5_w_ready;
	output wire m_axil_5_w_valid;
	output wire [63:0] m_axil_5_w_bits_data;
	output wire [7:0] m_axil_5_w_bits_strb;
	output wire m_axil_5_b_ready;
	input m_axil_5_b_valid;
	input [1:0] m_axil_5_b_bits_resp;
	wire _write_mux_io_sink_valid;
	wire [1:0] _write_mux_io_sink_bits_resp;
	wire _write_mux_io_select_ready;
	wire _write_demux_1_io_source_ready;
	wire _write_demux_1_io_select_ready;
	wire _write_demux_io_source_ready;
	wire _write_demux_io_select_ready;
	wire _write_portQueueB_io_enq_ready;
	wire _write_portQueueB_io_deq_valid;
	wire [2:0] _write_portQueueB_io_deq_bits;
	wire _write_portQueueW_io_enq_ready;
	wire _write_portQueueW_io_deq_valid;
	wire [2:0] _write_portQueueW_io_deq_bits;
	wire _read_mux_io_sink_valid;
	wire [63:0] _read_mux_io_sink_bits_data;
	wire [1:0] _read_mux_io_sink_bits_resp;
	wire _read_mux_io_select_ready;
	wire _read_demux_io_source_ready;
	wire _read_demux_io_select_ready;
	wire _read_portQueue_io_enq_ready;
	wire _read_portQueue_io_deq_valid;
	wire [2:0] _read_portQueue_io_deq_bits;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [11:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [11:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	reg read_eagerFork_regs_0;
	reg read_eagerFork_regs_1;
	reg read_eagerFork_regs_2;
	wire read_eagerFork_arPort_ready_qual1_0 = _read_demux_io_source_ready | read_eagerFork_regs_0;
	wire read_eagerFork_arPort_ready_qual1_1 = _read_demux_io_select_ready | read_eagerFork_regs_1;
	wire read_eagerFork_arPort_ready_qual1_2 = _read_portQueue_io_enq_ready | read_eagerFork_regs_2;
	wire read_result_ready = (read_eagerFork_arPort_ready_qual1_0 & read_eagerFork_arPort_ready_qual1_1) & read_eagerFork_arPort_ready_qual1_2;
	reg write_eagerFork_regs_0;
	reg write_eagerFork_regs_1;
	reg write_eagerFork_regs_2;
	reg write_eagerFork_regs_3;
	wire write_eagerFork_awPort_ready_qual1_0 = _write_demux_io_source_ready | write_eagerFork_regs_0;
	wire write_eagerFork_awPort_ready_qual1_1 = _write_demux_io_select_ready | write_eagerFork_regs_1;
	wire write_eagerFork_awPort_ready_qual1_2 = _write_portQueueW_io_enq_ready | write_eagerFork_regs_2;
	wire write_eagerFork_awPort_ready_qual1_3 = _write_portQueueB_io_enq_ready | write_eagerFork_regs_3;
	wire write_result_ready = ((write_eagerFork_awPort_ready_qual1_0 & write_eagerFork_awPort_ready_qual1_1) & write_eagerFork_awPort_ready_qual1_2) & write_eagerFork_awPort_ready_qual1_3;
	always @(posedge clock)
		if (reset) begin
			read_eagerFork_regs_0 <= 1'h0;
			read_eagerFork_regs_1 <= 1'h0;
			read_eagerFork_regs_2 <= 1'h0;
			write_eagerFork_regs_0 <= 1'h0;
			write_eagerFork_regs_1 <= 1'h0;
			write_eagerFork_regs_2 <= 1'h0;
			write_eagerFork_regs_3 <= 1'h0;
		end
		else begin
			read_eagerFork_regs_0 <= (read_eagerFork_arPort_ready_qual1_0 & _s_axil__sourceBuffer_io_deq_valid) & ~read_result_ready;
			read_eagerFork_regs_1 <= (read_eagerFork_arPort_ready_qual1_1 & _s_axil__sourceBuffer_io_deq_valid) & ~read_result_ready;
			read_eagerFork_regs_2 <= (read_eagerFork_arPort_ready_qual1_2 & _s_axil__sourceBuffer_io_deq_valid) & ~read_result_ready;
			write_eagerFork_regs_0 <= (write_eagerFork_awPort_ready_qual1_0 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
			write_eagerFork_regs_1 <= (write_eagerFork_awPort_ready_qual1_1 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
			write_eagerFork_regs_2 <= (write_eagerFork_awPort_ready_qual1_2 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
			write_eagerFork_regs_3 <= (write_eagerFork_awPort_ready_qual1_3 & _s_axil__sourceBuffer_1_io_deq_valid) & ~write_result_ready;
		end
	Queue2_AddressChannel s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axil_ar_ready),
		.io_enq_valid(s_axil_ar_valid),
		.io_enq_bits_addr(s_axil_ar_bits_addr),
		.io_enq_bits_prot(s_axil_ar_bits_prot),
		.io_deq_ready(read_result_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_read_mux_io_sink_valid),
		.io_enq_bits_data(_read_mux_io_sink_bits_data),
		.io_enq_bits_resp(_read_mux_io_sink_bits_resp),
		.io_deq_ready(s_axil_r_ready),
		.io_deq_valid(s_axil_r_valid),
		.io_deq_bits_data(s_axil_r_bits_data),
		.io_deq_bits_resp(s_axil_r_bits_resp)
	);
	Queue2_AddressChannel s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axil_aw_ready),
		.io_enq_valid(s_axil_aw_valid),
		.io_enq_bits_addr(s_axil_aw_bits_addr),
		.io_enq_bits_prot(s_axil_aw_bits_prot),
		.io_deq_ready(write_result_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(s_axil_w_ready),
		.io_enq_valid(s_axil_w_valid),
		.io_enq_bits_data(s_axil_w_bits_data),
		.io_enq_bits_strb(s_axil_w_bits_strb),
		.io_deq_ready(_write_demux_1_io_source_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_write_mux_io_sink_valid),
		.io_enq_bits_resp(_write_mux_io_sink_bits_resp),
		.io_deq_ready(s_axil_b_ready),
		.io_deq_valid(s_axil_b_valid),
		.io_deq_bits_resp(s_axil_b_bits_resp)
	);
	Queue8_UInt3 read_portQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_read_portQueue_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid & ~read_eagerFork_regs_2),
		.io_enq_bits(_s_axil__sourceBuffer_io_deq_bits_addr[8:6]),
		.io_deq_ready(_read_mux_io_select_ready),
		.io_deq_valid(_read_portQueue_io_deq_valid),
		.io_deq_bits(_read_portQueue_io_deq_bits)
	);
	elasticDemux read_demux(
		.io_source_ready(_read_demux_io_source_ready),
		.io_source_valid(_s_axil__sourceBuffer_io_deq_valid & ~read_eagerFork_regs_0),
		.io_source_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_source_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_sinks_0_ready(m_axil_0_ar_ready),
		.io_sinks_0_valid(m_axil_0_ar_valid),
		.io_sinks_0_bits_addr(m_axil_0_ar_bits_addr),
		.io_sinks_0_bits_prot(m_axil_0_ar_bits_prot),
		.io_sinks_1_ready(m_axil_1_ar_ready),
		.io_sinks_1_valid(m_axil_1_ar_valid),
		.io_sinks_1_bits_addr(m_axil_1_ar_bits_addr),
		.io_sinks_1_bits_prot(m_axil_1_ar_bits_prot),
		.io_sinks_2_ready(m_axil_2_ar_ready),
		.io_sinks_2_valid(m_axil_2_ar_valid),
		.io_sinks_2_bits_addr(m_axil_2_ar_bits_addr),
		.io_sinks_2_bits_prot(m_axil_2_ar_bits_prot),
		.io_sinks_3_ready(m_axil_3_ar_ready),
		.io_sinks_3_valid(m_axil_3_ar_valid),
		.io_sinks_3_bits_addr(m_axil_3_ar_bits_addr),
		.io_sinks_3_bits_prot(m_axil_3_ar_bits_prot),
		.io_sinks_4_ready(m_axil_4_ar_ready),
		.io_sinks_4_valid(m_axil_4_ar_valid),
		.io_sinks_4_bits_addr(m_axil_4_ar_bits_addr),
		.io_sinks_4_bits_prot(m_axil_4_ar_bits_prot),
		.io_sinks_5_ready(m_axil_5_ar_ready),
		.io_sinks_5_valid(m_axil_5_ar_valid),
		.io_sinks_5_bits_addr(m_axil_5_ar_bits_addr),
		.io_sinks_5_bits_prot(m_axil_5_ar_bits_prot),
		.io_select_ready(_read_demux_io_select_ready),
		.io_select_valid(_s_axil__sourceBuffer_io_deq_valid & ~read_eagerFork_regs_1),
		.io_select_bits(_s_axil__sourceBuffer_io_deq_bits_addr[8:6])
	);
	elasticMux read_mux(
		.io_sources_0_ready(m_axil_0_r_ready),
		.io_sources_0_valid(m_axil_0_r_valid),
		.io_sources_0_bits_data(m_axil_0_r_bits_data),
		.io_sources_0_bits_resp(m_axil_0_r_bits_resp),
		.io_sources_1_ready(m_axil_1_r_ready),
		.io_sources_1_valid(m_axil_1_r_valid),
		.io_sources_1_bits_data(m_axil_1_r_bits_data),
		.io_sources_1_bits_resp(m_axil_1_r_bits_resp),
		.io_sources_2_ready(m_axil_2_r_ready),
		.io_sources_2_valid(m_axil_2_r_valid),
		.io_sources_2_bits_data(m_axil_2_r_bits_data),
		.io_sources_2_bits_resp(m_axil_2_r_bits_resp),
		.io_sources_3_ready(m_axil_3_r_ready),
		.io_sources_3_valid(m_axil_3_r_valid),
		.io_sources_3_bits_data(m_axil_3_r_bits_data),
		.io_sources_3_bits_resp(m_axil_3_r_bits_resp),
		.io_sources_4_ready(m_axil_4_r_ready),
		.io_sources_4_valid(m_axil_4_r_valid),
		.io_sources_4_bits_data(m_axil_4_r_bits_data),
		.io_sources_4_bits_resp(m_axil_4_r_bits_resp),
		.io_sources_5_ready(m_axil_5_r_ready),
		.io_sources_5_valid(m_axil_5_r_valid),
		.io_sources_5_bits_data(m_axil_5_r_bits_data),
		.io_sources_5_bits_resp(m_axil_5_r_bits_resp),
		.io_sink_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_sink_valid(_read_mux_io_sink_valid),
		.io_sink_bits_data(_read_mux_io_sink_bits_data),
		.io_sink_bits_resp(_read_mux_io_sink_bits_resp),
		.io_select_ready(_read_mux_io_select_ready),
		.io_select_valid(_read_portQueue_io_deq_valid),
		.io_select_bits(_read_portQueue_io_deq_bits)
	);
	Queue8_UInt3 write_portQueueW(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueueW_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_2),
		.io_enq_bits(_s_axil__sourceBuffer_1_io_deq_bits_addr[8:6]),
		.io_deq_ready(_write_demux_1_io_select_ready),
		.io_deq_valid(_write_portQueueW_io_deq_valid),
		.io_deq_bits(_write_portQueueW_io_deq_bits)
	);
	Queue8_UInt3 write_portQueueB(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_write_portQueueB_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_3),
		.io_enq_bits(_s_axil__sourceBuffer_1_io_deq_bits_addr[8:6]),
		.io_deq_ready(_write_mux_io_select_ready),
		.io_deq_valid(_write_portQueueB_io_deq_valid),
		.io_deq_bits(_write_portQueueB_io_deq_bits)
	);
	elasticDemux write_demux(
		.io_source_ready(_write_demux_io_source_ready),
		.io_source_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_0),
		.io_source_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_source_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_sinks_0_ready(m_axil_0_aw_ready),
		.io_sinks_0_valid(m_axil_0_aw_valid),
		.io_sinks_0_bits_addr(m_axil_0_aw_bits_addr),
		.io_sinks_0_bits_prot(m_axil_0_aw_bits_prot),
		.io_sinks_1_ready(m_axil_1_aw_ready),
		.io_sinks_1_valid(m_axil_1_aw_valid),
		.io_sinks_1_bits_addr(m_axil_1_aw_bits_addr),
		.io_sinks_1_bits_prot(m_axil_1_aw_bits_prot),
		.io_sinks_2_ready(m_axil_2_aw_ready),
		.io_sinks_2_valid(m_axil_2_aw_valid),
		.io_sinks_2_bits_addr(m_axil_2_aw_bits_addr),
		.io_sinks_2_bits_prot(m_axil_2_aw_bits_prot),
		.io_sinks_3_ready(m_axil_3_aw_ready),
		.io_sinks_3_valid(m_axil_3_aw_valid),
		.io_sinks_3_bits_addr(m_axil_3_aw_bits_addr),
		.io_sinks_3_bits_prot(m_axil_3_aw_bits_prot),
		.io_sinks_4_ready(m_axil_4_aw_ready),
		.io_sinks_4_valid(m_axil_4_aw_valid),
		.io_sinks_4_bits_addr(m_axil_4_aw_bits_addr),
		.io_sinks_4_bits_prot(m_axil_4_aw_bits_prot),
		.io_sinks_5_ready(m_axil_5_aw_ready),
		.io_sinks_5_valid(m_axil_5_aw_valid),
		.io_sinks_5_bits_addr(m_axil_5_aw_bits_addr),
		.io_sinks_5_bits_prot(m_axil_5_aw_bits_prot),
		.io_select_ready(_write_demux_io_select_ready),
		.io_select_valid(_s_axil__sourceBuffer_1_io_deq_valid & ~write_eagerFork_regs_1),
		.io_select_bits(_s_axil__sourceBuffer_1_io_deq_bits_addr[8:6])
	);
	elasticDemux_2 write_demux_1(
		.io_source_ready(_write_demux_1_io_source_ready),
		.io_source_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_source_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_source_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_sinks_0_ready(m_axil_0_w_ready),
		.io_sinks_0_valid(m_axil_0_w_valid),
		.io_sinks_0_bits_data(m_axil_0_w_bits_data),
		.io_sinks_0_bits_strb(m_axil_0_w_bits_strb),
		.io_sinks_1_ready(m_axil_1_w_ready),
		.io_sinks_1_valid(m_axil_1_w_valid),
		.io_sinks_1_bits_data(m_axil_1_w_bits_data),
		.io_sinks_1_bits_strb(m_axil_1_w_bits_strb),
		.io_sinks_2_ready(m_axil_2_w_ready),
		.io_sinks_2_valid(m_axil_2_w_valid),
		.io_sinks_2_bits_data(m_axil_2_w_bits_data),
		.io_sinks_2_bits_strb(m_axil_2_w_bits_strb),
		.io_sinks_3_ready(m_axil_3_w_ready),
		.io_sinks_3_valid(m_axil_3_w_valid),
		.io_sinks_3_bits_data(m_axil_3_w_bits_data),
		.io_sinks_3_bits_strb(m_axil_3_w_bits_strb),
		.io_sinks_4_ready(m_axil_4_w_ready),
		.io_sinks_4_valid(m_axil_4_w_valid),
		.io_sinks_4_bits_data(m_axil_4_w_bits_data),
		.io_sinks_4_bits_strb(m_axil_4_w_bits_strb),
		.io_sinks_5_ready(m_axil_5_w_ready),
		.io_sinks_5_valid(m_axil_5_w_valid),
		.io_sinks_5_bits_data(m_axil_5_w_bits_data),
		.io_sinks_5_bits_strb(m_axil_5_w_bits_strb),
		.io_select_ready(_write_demux_1_io_select_ready),
		.io_select_valid(_write_portQueueW_io_deq_valid),
		.io_select_bits(_write_portQueueW_io_deq_bits)
	);
	elasticMux_1 write_mux(
		.io_sources_0_ready(m_axil_0_b_ready),
		.io_sources_0_valid(m_axil_0_b_valid),
		.io_sources_0_bits_resp(m_axil_0_b_bits_resp),
		.io_sources_1_ready(m_axil_1_b_ready),
		.io_sources_1_valid(m_axil_1_b_valid),
		.io_sources_1_bits_resp(m_axil_1_b_bits_resp),
		.io_sources_2_ready(m_axil_2_b_ready),
		.io_sources_2_valid(m_axil_2_b_valid),
		.io_sources_2_bits_resp(m_axil_2_b_bits_resp),
		.io_sources_3_ready(m_axil_3_b_ready),
		.io_sources_3_valid(m_axil_3_b_valid),
		.io_sources_3_bits_resp(m_axil_3_b_bits_resp),
		.io_sources_4_ready(m_axil_4_b_ready),
		.io_sources_4_valid(m_axil_4_b_valid),
		.io_sources_4_bits_resp(m_axil_4_b_bits_resp),
		.io_sources_5_ready(m_axil_5_b_ready),
		.io_sources_5_valid(m_axil_5_b_valid),
		.io_sources_5_bits_resp(m_axil_5_b_bits_resp),
		.io_sink_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_sink_valid(_write_mux_io_sink_valid),
		.io_sink_bits_resp(_write_mux_io_sink_bits_resp),
		.io_select_ready(_write_mux_io_select_ready),
		.io_select_valid(_write_portQueueB_io_deq_valid),
		.io_select_bits(_write_portQueueB_io_deq_bits)
	);
endmodule
module SchedulerNetworkDataUnit (
	clock,
	reset,
	io_taskIn,
	io_taskOut,
	io_validIn,
	io_validOut,
	io_connSS_availableTask_ready,
	io_connSS_availableTask_valid,
	io_connSS_availableTask_bits,
	io_connSS_qOutTask_ready,
	io_connSS_qOutTask_valid,
	io_connSS_qOutTask_bits,
	io_occupied
);
	input clock;
	input reset;
	input [255:0] io_taskIn;
	output wire [255:0] io_taskOut;
	input io_validIn;
	output wire io_validOut;
	input io_connSS_availableTask_ready;
	output wire io_connSS_availableTask_valid;
	output wire [255:0] io_connSS_availableTask_bits;
	output wire io_connSS_qOutTask_ready;
	input io_connSS_qOutTask_valid;
	input [255:0] io_connSS_qOutTask_bits;
	output wire io_occupied;
	reg [255:0] taskReg;
	reg validReg;
	wire io_connSS_availableTask_valid_0 = io_connSS_availableTask_ready & io_validIn;
	wire _GEN = io_connSS_qOutTask_valid & ~io_validIn;
	always @(posedge clock)
		if (reset) begin
			taskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			validReg <= 1'h0;
		end
		else begin
			taskReg <= (io_connSS_availableTask_valid_0 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : (_GEN ? io_connSS_qOutTask_bits : (io_validIn ? io_taskIn : 256'h0000000000000000000000000000000000000000000000000000000000000000)));
			validReg <= ~io_connSS_availableTask_valid_0 & (_GEN | io_validIn);
		end
	assign io_taskOut = taskReg;
	assign io_validOut = validReg;
	assign io_connSS_availableTask_valid = io_connSS_availableTask_valid_0;
	assign io_connSS_availableTask_bits = (io_connSS_availableTask_valid_0 ? io_taskIn : 256'h0000000000000000000000000000000000000000000000000000000000000000);
	assign io_connSS_qOutTask_ready = ~io_connSS_availableTask_valid_0 & _GEN;
	assign io_occupied = validReg;
endmodule
module SchedulerNetworkControlUnit (
	clock,
	reset,
	io_reqTaskIn,
	io_reqTaskOut,
	io_connSS_serveStealReq_valid,
	io_connSS_serveStealReq_ready,
	io_connSS_stealReq_valid,
	io_connSS_stealReq_ready
);
	input clock;
	input reset;
	input io_reqTaskIn;
	output wire io_reqTaskOut;
	input io_connSS_serveStealReq_valid;
	output wire io_connSS_serveStealReq_ready;
	input io_connSS_stealReq_valid;
	output wire io_connSS_stealReq_ready;
	reg stealReqReg;
	always @(posedge clock)
		if (reset)
			stealReqReg <= 1'h0;
		else
			stealReqReg <= io_reqTaskIn;
	assign io_reqTaskOut = io_connSS_stealReq_valid | (~io_connSS_serveStealReq_valid & stealReqReg);
	assign io_connSS_serveStealReq_ready = stealReqReg;
	assign io_connSS_stealReq_ready = ~stealReqReg;
endmodule
module SchedulerNetwork (
	clock,
	reset,
	io_connSS_0_ctrl_serveStealReq_valid,
	io_connSS_0_ctrl_serveStealReq_ready,
	io_connSS_0_data_availableTask_ready,
	io_connSS_0_data_availableTask_valid,
	io_connSS_0_data_availableTask_bits,
	io_connSS_0_data_qOutTask_ready,
	io_connSS_0_data_qOutTask_valid,
	io_connSS_0_data_qOutTask_bits,
	io_connSS_1_ctrl_serveStealReq_valid,
	io_connSS_1_ctrl_serveStealReq_ready,
	io_connSS_1_ctrl_stealReq_valid,
	io_connSS_1_ctrl_stealReq_ready,
	io_connSS_1_data_availableTask_ready,
	io_connSS_1_data_availableTask_valid,
	io_connSS_1_data_availableTask_bits,
	io_connSS_1_data_qOutTask_ready,
	io_connSS_1_data_qOutTask_valid,
	io_connSS_1_data_qOutTask_bits,
	io_connSS_2_ctrl_serveStealReq_valid,
	io_connSS_2_ctrl_serveStealReq_ready,
	io_connSS_2_ctrl_stealReq_valid,
	io_connSS_2_ctrl_stealReq_ready,
	io_connSS_2_data_availableTask_ready,
	io_connSS_2_data_availableTask_valid,
	io_connSS_2_data_availableTask_bits,
	io_connSS_2_data_qOutTask_ready,
	io_connSS_2_data_qOutTask_valid,
	io_connSS_2_data_qOutTask_bits,
	io_connSS_3_ctrl_serveStealReq_valid,
	io_connSS_3_ctrl_serveStealReq_ready,
	io_connSS_3_ctrl_stealReq_valid,
	io_connSS_3_ctrl_stealReq_ready,
	io_connSS_3_data_availableTask_ready,
	io_connSS_3_data_availableTask_valid,
	io_connSS_3_data_availableTask_bits,
	io_connSS_3_data_qOutTask_ready,
	io_connSS_3_data_qOutTask_valid,
	io_connSS_3_data_qOutTask_bits,
	io_connSS_4_ctrl_serveStealReq_valid,
	io_connSS_4_ctrl_serveStealReq_ready,
	io_connSS_4_ctrl_stealReq_valid,
	io_connSS_4_ctrl_stealReq_ready,
	io_connSS_4_data_availableTask_ready,
	io_connSS_4_data_availableTask_valid,
	io_connSS_4_data_availableTask_bits,
	io_connSS_4_data_qOutTask_ready,
	io_connSS_4_data_qOutTask_valid,
	io_connSS_4_data_qOutTask_bits,
	io_connSS_5_ctrl_serveStealReq_valid,
	io_connSS_5_ctrl_serveStealReq_ready,
	io_connSS_5_ctrl_stealReq_valid,
	io_connSS_5_ctrl_stealReq_ready,
	io_connSS_5_data_availableTask_ready,
	io_connSS_5_data_availableTask_valid,
	io_connSS_5_data_availableTask_bits,
	io_connSS_5_data_qOutTask_ready,
	io_connSS_5_data_qOutTask_valid,
	io_connSS_5_data_qOutTask_bits,
	io_connSS_6_ctrl_serveStealReq_valid,
	io_connSS_6_ctrl_serveStealReq_ready,
	io_connSS_6_ctrl_stealReq_valid,
	io_connSS_6_ctrl_stealReq_ready,
	io_connSS_6_data_availableTask_ready,
	io_connSS_6_data_availableTask_valid,
	io_connSS_6_data_availableTask_bits,
	io_connSS_6_data_qOutTask_ready,
	io_connSS_6_data_qOutTask_valid,
	io_connSS_6_data_qOutTask_bits,
	io_connSS_7_ctrl_serveStealReq_valid,
	io_connSS_7_ctrl_serveStealReq_ready,
	io_connSS_7_ctrl_stealReq_valid,
	io_connSS_7_ctrl_stealReq_ready,
	io_connSS_7_data_availableTask_ready,
	io_connSS_7_data_availableTask_valid,
	io_connSS_7_data_availableTask_bits,
	io_connSS_7_data_qOutTask_ready,
	io_connSS_7_data_qOutTask_valid,
	io_connSS_7_data_qOutTask_bits,
	io_connSS_8_ctrl_serveStealReq_valid,
	io_connSS_8_ctrl_serveStealReq_ready,
	io_connSS_8_ctrl_stealReq_valid,
	io_connSS_8_ctrl_stealReq_ready,
	io_connSS_8_data_availableTask_ready,
	io_connSS_8_data_availableTask_valid,
	io_connSS_8_data_availableTask_bits,
	io_connSS_8_data_qOutTask_ready,
	io_connSS_8_data_qOutTask_valid,
	io_connSS_8_data_qOutTask_bits,
	io_connSS_9_ctrl_serveStealReq_valid,
	io_connSS_9_ctrl_serveStealReq_ready,
	io_connSS_9_ctrl_stealReq_valid,
	io_connSS_9_ctrl_stealReq_ready,
	io_connSS_9_data_availableTask_ready,
	io_connSS_9_data_availableTask_valid,
	io_connSS_9_data_availableTask_bits,
	io_connSS_9_data_qOutTask_ready,
	io_connSS_9_data_qOutTask_valid,
	io_connSS_9_data_qOutTask_bits,
	io_connSS_10_ctrl_serveStealReq_valid,
	io_connSS_10_ctrl_serveStealReq_ready,
	io_connSS_10_ctrl_stealReq_valid,
	io_connSS_10_ctrl_stealReq_ready,
	io_connSS_10_data_availableTask_ready,
	io_connSS_10_data_availableTask_valid,
	io_connSS_10_data_availableTask_bits,
	io_connSS_10_data_qOutTask_ready,
	io_connSS_10_data_qOutTask_valid,
	io_connSS_10_data_qOutTask_bits,
	io_connSS_11_ctrl_serveStealReq_valid,
	io_connSS_11_ctrl_serveStealReq_ready,
	io_connSS_11_ctrl_stealReq_valid,
	io_connSS_11_ctrl_stealReq_ready,
	io_connSS_11_data_availableTask_ready,
	io_connSS_11_data_availableTask_valid,
	io_connSS_11_data_availableTask_bits,
	io_connSS_11_data_qOutTask_ready,
	io_connSS_11_data_qOutTask_valid,
	io_connSS_11_data_qOutTask_bits,
	io_connSS_12_ctrl_serveStealReq_valid,
	io_connSS_12_ctrl_serveStealReq_ready,
	io_connSS_12_ctrl_stealReq_valid,
	io_connSS_12_ctrl_stealReq_ready,
	io_connSS_12_data_availableTask_ready,
	io_connSS_12_data_availableTask_valid,
	io_connSS_12_data_availableTask_bits,
	io_connSS_12_data_qOutTask_ready,
	io_connSS_12_data_qOutTask_valid,
	io_connSS_12_data_qOutTask_bits,
	io_connSS_13_ctrl_serveStealReq_valid,
	io_connSS_13_ctrl_serveStealReq_ready,
	io_connSS_13_ctrl_stealReq_valid,
	io_connSS_13_ctrl_stealReq_ready,
	io_connSS_13_data_availableTask_ready,
	io_connSS_13_data_availableTask_valid,
	io_connSS_13_data_availableTask_bits,
	io_connSS_13_data_qOutTask_ready,
	io_connSS_13_data_qOutTask_valid,
	io_connSS_13_data_qOutTask_bits,
	io_connSS_14_ctrl_serveStealReq_valid,
	io_connSS_14_ctrl_serveStealReq_ready,
	io_connSS_14_ctrl_stealReq_valid,
	io_connSS_14_ctrl_stealReq_ready,
	io_connSS_14_data_availableTask_ready,
	io_connSS_14_data_availableTask_valid,
	io_connSS_14_data_availableTask_bits,
	io_connSS_14_data_qOutTask_ready,
	io_connSS_14_data_qOutTask_valid,
	io_connSS_14_data_qOutTask_bits,
	io_connSS_15_ctrl_serveStealReq_valid,
	io_connSS_15_ctrl_serveStealReq_ready,
	io_connSS_15_ctrl_stealReq_valid,
	io_connSS_15_ctrl_stealReq_ready,
	io_connSS_15_data_availableTask_ready,
	io_connSS_15_data_availableTask_valid,
	io_connSS_15_data_availableTask_bits,
	io_connSS_15_data_qOutTask_ready,
	io_connSS_15_data_qOutTask_valid,
	io_connSS_15_data_qOutTask_bits,
	io_connSS_16_ctrl_serveStealReq_valid,
	io_connSS_16_ctrl_serveStealReq_ready,
	io_connSS_16_ctrl_stealReq_valid,
	io_connSS_16_ctrl_stealReq_ready,
	io_connSS_16_data_availableTask_ready,
	io_connSS_16_data_availableTask_valid,
	io_connSS_16_data_availableTask_bits,
	io_connSS_16_data_qOutTask_ready,
	io_connSS_16_data_qOutTask_valid,
	io_connSS_16_data_qOutTask_bits,
	io_connSS_17_ctrl_serveStealReq_valid,
	io_connSS_17_ctrl_serveStealReq_ready,
	io_connSS_17_ctrl_stealReq_valid,
	io_connSS_17_ctrl_stealReq_ready,
	io_connSS_17_data_availableTask_ready,
	io_connSS_17_data_availableTask_valid,
	io_connSS_17_data_availableTask_bits,
	io_connSS_17_data_qOutTask_ready,
	io_connSS_17_data_qOutTask_valid,
	io_connSS_17_data_qOutTask_bits,
	io_connSS_18_ctrl_serveStealReq_valid,
	io_connSS_18_ctrl_serveStealReq_ready,
	io_connSS_18_ctrl_stealReq_valid,
	io_connSS_18_ctrl_stealReq_ready,
	io_connSS_18_data_availableTask_ready,
	io_connSS_18_data_availableTask_valid,
	io_connSS_18_data_availableTask_bits,
	io_connSS_18_data_qOutTask_ready,
	io_connSS_18_data_qOutTask_valid,
	io_connSS_18_data_qOutTask_bits,
	io_connSS_19_ctrl_serveStealReq_valid,
	io_connSS_19_ctrl_serveStealReq_ready,
	io_connSS_19_ctrl_stealReq_valid,
	io_connSS_19_ctrl_stealReq_ready,
	io_connSS_19_data_availableTask_ready,
	io_connSS_19_data_availableTask_valid,
	io_connSS_19_data_availableTask_bits,
	io_connSS_19_data_qOutTask_ready,
	io_connSS_19_data_qOutTask_valid,
	io_connSS_19_data_qOutTask_bits,
	io_connSS_20_ctrl_serveStealReq_valid,
	io_connSS_20_ctrl_serveStealReq_ready,
	io_connSS_20_ctrl_stealReq_valid,
	io_connSS_20_ctrl_stealReq_ready,
	io_connSS_20_data_availableTask_ready,
	io_connSS_20_data_availableTask_valid,
	io_connSS_20_data_availableTask_bits,
	io_connSS_20_data_qOutTask_ready,
	io_connSS_20_data_qOutTask_valid,
	io_connSS_20_data_qOutTask_bits,
	io_connSS_21_ctrl_serveStealReq_valid,
	io_connSS_21_ctrl_serveStealReq_ready,
	io_connSS_21_ctrl_stealReq_valid,
	io_connSS_21_ctrl_stealReq_ready,
	io_connSS_21_data_availableTask_ready,
	io_connSS_21_data_availableTask_valid,
	io_connSS_21_data_availableTask_bits,
	io_connSS_21_data_qOutTask_ready,
	io_connSS_21_data_qOutTask_valid,
	io_connSS_21_data_qOutTask_bits,
	io_connSS_22_ctrl_serveStealReq_valid,
	io_connSS_22_ctrl_serveStealReq_ready,
	io_connSS_22_ctrl_stealReq_valid,
	io_connSS_22_ctrl_stealReq_ready,
	io_connSS_22_data_availableTask_ready,
	io_connSS_22_data_availableTask_valid,
	io_connSS_22_data_availableTask_bits,
	io_connSS_22_data_qOutTask_ready,
	io_connSS_22_data_qOutTask_valid,
	io_connSS_22_data_qOutTask_bits,
	io_connSS_23_ctrl_serveStealReq_valid,
	io_connSS_23_ctrl_serveStealReq_ready,
	io_connSS_23_ctrl_stealReq_valid,
	io_connSS_23_ctrl_stealReq_ready,
	io_connSS_23_data_availableTask_ready,
	io_connSS_23_data_availableTask_valid,
	io_connSS_23_data_availableTask_bits,
	io_connSS_23_data_qOutTask_ready,
	io_connSS_23_data_qOutTask_valid,
	io_connSS_23_data_qOutTask_bits,
	io_connSS_24_ctrl_serveStealReq_valid,
	io_connSS_24_ctrl_serveStealReq_ready,
	io_connSS_24_ctrl_stealReq_valid,
	io_connSS_24_ctrl_stealReq_ready,
	io_connSS_24_data_availableTask_ready,
	io_connSS_24_data_availableTask_valid,
	io_connSS_24_data_availableTask_bits,
	io_connSS_24_data_qOutTask_ready,
	io_connSS_24_data_qOutTask_valid,
	io_connSS_24_data_qOutTask_bits,
	io_connSS_25_ctrl_serveStealReq_valid,
	io_connSS_25_ctrl_serveStealReq_ready,
	io_connSS_25_ctrl_stealReq_valid,
	io_connSS_25_ctrl_stealReq_ready,
	io_connSS_25_data_availableTask_ready,
	io_connSS_25_data_availableTask_valid,
	io_connSS_25_data_availableTask_bits,
	io_connSS_25_data_qOutTask_ready,
	io_connSS_25_data_qOutTask_valid,
	io_connSS_25_data_qOutTask_bits,
	io_connSS_26_ctrl_serveStealReq_valid,
	io_connSS_26_ctrl_serveStealReq_ready,
	io_connSS_26_ctrl_stealReq_valid,
	io_connSS_26_ctrl_stealReq_ready,
	io_connSS_26_data_availableTask_ready,
	io_connSS_26_data_availableTask_valid,
	io_connSS_26_data_availableTask_bits,
	io_connSS_26_data_qOutTask_ready,
	io_connSS_26_data_qOutTask_valid,
	io_connSS_26_data_qOutTask_bits,
	io_connSS_27_ctrl_serveStealReq_valid,
	io_connSS_27_ctrl_serveStealReq_ready,
	io_connSS_27_ctrl_stealReq_valid,
	io_connSS_27_ctrl_stealReq_ready,
	io_connSS_27_data_availableTask_ready,
	io_connSS_27_data_availableTask_valid,
	io_connSS_27_data_availableTask_bits,
	io_connSS_27_data_qOutTask_ready,
	io_connSS_27_data_qOutTask_valid,
	io_connSS_27_data_qOutTask_bits,
	io_connSS_28_ctrl_serveStealReq_valid,
	io_connSS_28_ctrl_serveStealReq_ready,
	io_connSS_28_ctrl_stealReq_valid,
	io_connSS_28_ctrl_stealReq_ready,
	io_connSS_28_data_availableTask_ready,
	io_connSS_28_data_availableTask_valid,
	io_connSS_28_data_availableTask_bits,
	io_connSS_28_data_qOutTask_ready,
	io_connSS_28_data_qOutTask_valid,
	io_connSS_28_data_qOutTask_bits,
	io_connSS_29_ctrl_serveStealReq_valid,
	io_connSS_29_ctrl_serveStealReq_ready,
	io_connSS_29_ctrl_stealReq_valid,
	io_connSS_29_ctrl_stealReq_ready,
	io_connSS_29_data_availableTask_ready,
	io_connSS_29_data_availableTask_valid,
	io_connSS_29_data_availableTask_bits,
	io_connSS_29_data_qOutTask_ready,
	io_connSS_29_data_qOutTask_valid,
	io_connSS_29_data_qOutTask_bits,
	io_connSS_30_ctrl_serveStealReq_valid,
	io_connSS_30_ctrl_serveStealReq_ready,
	io_connSS_30_ctrl_stealReq_valid,
	io_connSS_30_ctrl_stealReq_ready,
	io_connSS_30_data_availableTask_ready,
	io_connSS_30_data_availableTask_valid,
	io_connSS_30_data_availableTask_bits,
	io_connSS_30_data_qOutTask_ready,
	io_connSS_30_data_qOutTask_valid,
	io_connSS_30_data_qOutTask_bits,
	io_connSS_31_ctrl_serveStealReq_valid,
	io_connSS_31_ctrl_serveStealReq_ready,
	io_connSS_31_ctrl_stealReq_valid,
	io_connSS_31_ctrl_stealReq_ready,
	io_connSS_31_data_availableTask_ready,
	io_connSS_31_data_availableTask_valid,
	io_connSS_31_data_availableTask_bits,
	io_connSS_31_data_qOutTask_ready,
	io_connSS_31_data_qOutTask_valid,
	io_connSS_31_data_qOutTask_bits,
	io_connSS_32_ctrl_serveStealReq_valid,
	io_connSS_32_ctrl_serveStealReq_ready,
	io_connSS_32_ctrl_stealReq_valid,
	io_connSS_32_ctrl_stealReq_ready,
	io_connSS_32_data_availableTask_ready,
	io_connSS_32_data_availableTask_valid,
	io_connSS_32_data_availableTask_bits,
	io_connSS_32_data_qOutTask_ready,
	io_connSS_32_data_qOutTask_valid,
	io_connSS_32_data_qOutTask_bits,
	io_connSS_33_ctrl_serveStealReq_valid,
	io_connSS_33_ctrl_serveStealReq_ready,
	io_connSS_33_ctrl_stealReq_valid,
	io_connSS_33_ctrl_stealReq_ready,
	io_connSS_33_data_availableTask_ready,
	io_connSS_33_data_availableTask_valid,
	io_connSS_33_data_availableTask_bits,
	io_connSS_33_data_qOutTask_ready,
	io_connSS_33_data_qOutTask_valid,
	io_connSS_33_data_qOutTask_bits,
	io_connSS_34_ctrl_serveStealReq_valid,
	io_connSS_34_ctrl_serveStealReq_ready,
	io_connSS_34_ctrl_stealReq_valid,
	io_connSS_34_ctrl_stealReq_ready,
	io_connSS_34_data_availableTask_ready,
	io_connSS_34_data_availableTask_valid,
	io_connSS_34_data_availableTask_bits,
	io_connSS_34_data_qOutTask_ready,
	io_connSS_34_data_qOutTask_valid,
	io_connSS_34_data_qOutTask_bits,
	io_connSS_35_ctrl_serveStealReq_valid,
	io_connSS_35_ctrl_serveStealReq_ready,
	io_connSS_35_ctrl_stealReq_valid,
	io_connSS_35_ctrl_stealReq_ready,
	io_connSS_35_data_availableTask_ready,
	io_connSS_35_data_availableTask_valid,
	io_connSS_35_data_availableTask_bits,
	io_connSS_35_data_qOutTask_ready,
	io_connSS_35_data_qOutTask_valid,
	io_connSS_35_data_qOutTask_bits,
	io_connSS_36_ctrl_serveStealReq_valid,
	io_connSS_36_ctrl_serveStealReq_ready,
	io_connSS_36_ctrl_stealReq_valid,
	io_connSS_36_ctrl_stealReq_ready,
	io_connSS_36_data_availableTask_ready,
	io_connSS_36_data_availableTask_valid,
	io_connSS_36_data_availableTask_bits,
	io_connSS_36_data_qOutTask_ready,
	io_connSS_36_data_qOutTask_valid,
	io_connSS_36_data_qOutTask_bits,
	io_connSS_37_ctrl_serveStealReq_valid,
	io_connSS_37_ctrl_serveStealReq_ready,
	io_connSS_37_ctrl_stealReq_valid,
	io_connSS_37_ctrl_stealReq_ready,
	io_connSS_37_data_availableTask_ready,
	io_connSS_37_data_availableTask_valid,
	io_connSS_37_data_availableTask_bits,
	io_connSS_37_data_qOutTask_ready,
	io_connSS_37_data_qOutTask_valid,
	io_connSS_37_data_qOutTask_bits,
	io_connSS_38_ctrl_serveStealReq_valid,
	io_connSS_38_ctrl_serveStealReq_ready,
	io_connSS_38_ctrl_stealReq_valid,
	io_connSS_38_ctrl_stealReq_ready,
	io_connSS_38_data_availableTask_ready,
	io_connSS_38_data_availableTask_valid,
	io_connSS_38_data_availableTask_bits,
	io_connSS_38_data_qOutTask_ready,
	io_connSS_38_data_qOutTask_valid,
	io_connSS_38_data_qOutTask_bits,
	io_connSS_39_ctrl_serveStealReq_valid,
	io_connSS_39_ctrl_serveStealReq_ready,
	io_connSS_39_ctrl_stealReq_valid,
	io_connSS_39_ctrl_stealReq_ready,
	io_connSS_39_data_availableTask_ready,
	io_connSS_39_data_availableTask_valid,
	io_connSS_39_data_availableTask_bits,
	io_connSS_39_data_qOutTask_ready,
	io_connSS_39_data_qOutTask_valid,
	io_connSS_39_data_qOutTask_bits,
	io_connSS_40_ctrl_serveStealReq_valid,
	io_connSS_40_ctrl_serveStealReq_ready,
	io_connSS_40_ctrl_stealReq_valid,
	io_connSS_40_ctrl_stealReq_ready,
	io_connSS_40_data_availableTask_ready,
	io_connSS_40_data_availableTask_valid,
	io_connSS_40_data_availableTask_bits,
	io_connSS_40_data_qOutTask_ready,
	io_connSS_40_data_qOutTask_valid,
	io_connSS_40_data_qOutTask_bits,
	io_connSS_41_ctrl_serveStealReq_valid,
	io_connSS_41_ctrl_serveStealReq_ready,
	io_connSS_41_ctrl_stealReq_valid,
	io_connSS_41_ctrl_stealReq_ready,
	io_connSS_41_data_availableTask_ready,
	io_connSS_41_data_availableTask_valid,
	io_connSS_41_data_availableTask_bits,
	io_connSS_41_data_qOutTask_ready,
	io_connSS_41_data_qOutTask_valid,
	io_connSS_41_data_qOutTask_bits,
	io_connSS_42_ctrl_serveStealReq_valid,
	io_connSS_42_ctrl_serveStealReq_ready,
	io_connSS_42_ctrl_stealReq_valid,
	io_connSS_42_ctrl_stealReq_ready,
	io_connSS_42_data_availableTask_ready,
	io_connSS_42_data_availableTask_valid,
	io_connSS_42_data_availableTask_bits,
	io_connSS_42_data_qOutTask_ready,
	io_connSS_42_data_qOutTask_valid,
	io_connSS_42_data_qOutTask_bits,
	io_connSS_43_ctrl_serveStealReq_valid,
	io_connSS_43_ctrl_serveStealReq_ready,
	io_connSS_43_ctrl_stealReq_valid,
	io_connSS_43_ctrl_stealReq_ready,
	io_connSS_43_data_availableTask_ready,
	io_connSS_43_data_availableTask_valid,
	io_connSS_43_data_availableTask_bits,
	io_connSS_43_data_qOutTask_ready,
	io_connSS_43_data_qOutTask_valid,
	io_connSS_43_data_qOutTask_bits,
	io_connSS_44_ctrl_serveStealReq_valid,
	io_connSS_44_ctrl_serveStealReq_ready,
	io_connSS_44_ctrl_stealReq_valid,
	io_connSS_44_ctrl_stealReq_ready,
	io_connSS_44_data_availableTask_ready,
	io_connSS_44_data_availableTask_valid,
	io_connSS_44_data_availableTask_bits,
	io_connSS_44_data_qOutTask_ready,
	io_connSS_44_data_qOutTask_valid,
	io_connSS_44_data_qOutTask_bits,
	io_connSS_45_ctrl_serveStealReq_valid,
	io_connSS_45_ctrl_serveStealReq_ready,
	io_connSS_45_ctrl_stealReq_valid,
	io_connSS_45_ctrl_stealReq_ready,
	io_connSS_45_data_availableTask_ready,
	io_connSS_45_data_availableTask_valid,
	io_connSS_45_data_availableTask_bits,
	io_connSS_45_data_qOutTask_ready,
	io_connSS_45_data_qOutTask_valid,
	io_connSS_45_data_qOutTask_bits,
	io_connSS_46_ctrl_serveStealReq_valid,
	io_connSS_46_ctrl_serveStealReq_ready,
	io_connSS_46_ctrl_stealReq_valid,
	io_connSS_46_ctrl_stealReq_ready,
	io_connSS_46_data_availableTask_ready,
	io_connSS_46_data_availableTask_valid,
	io_connSS_46_data_availableTask_bits,
	io_connSS_46_data_qOutTask_ready,
	io_connSS_46_data_qOutTask_valid,
	io_connSS_46_data_qOutTask_bits,
	io_connSS_47_ctrl_serveStealReq_valid,
	io_connSS_47_ctrl_serveStealReq_ready,
	io_connSS_47_ctrl_stealReq_valid,
	io_connSS_47_ctrl_stealReq_ready,
	io_connSS_47_data_availableTask_ready,
	io_connSS_47_data_availableTask_valid,
	io_connSS_47_data_availableTask_bits,
	io_connSS_47_data_qOutTask_ready,
	io_connSS_47_data_qOutTask_valid,
	io_connSS_47_data_qOutTask_bits,
	io_connSS_48_ctrl_serveStealReq_valid,
	io_connSS_48_ctrl_serveStealReq_ready,
	io_connSS_48_ctrl_stealReq_valid,
	io_connSS_48_ctrl_stealReq_ready,
	io_connSS_48_data_availableTask_ready,
	io_connSS_48_data_availableTask_valid,
	io_connSS_48_data_availableTask_bits,
	io_connSS_48_data_qOutTask_ready,
	io_connSS_48_data_qOutTask_valid,
	io_connSS_48_data_qOutTask_bits,
	io_connSS_49_ctrl_serveStealReq_valid,
	io_connSS_49_ctrl_serveStealReq_ready,
	io_connSS_49_ctrl_stealReq_valid,
	io_connSS_49_ctrl_stealReq_ready,
	io_connSS_49_data_availableTask_ready,
	io_connSS_49_data_availableTask_valid,
	io_connSS_49_data_availableTask_bits,
	io_connSS_49_data_qOutTask_ready,
	io_connSS_49_data_qOutTask_valid,
	io_connSS_49_data_qOutTask_bits,
	io_connSS_50_ctrl_serveStealReq_valid,
	io_connSS_50_ctrl_serveStealReq_ready,
	io_connSS_50_ctrl_stealReq_valid,
	io_connSS_50_ctrl_stealReq_ready,
	io_connSS_50_data_availableTask_ready,
	io_connSS_50_data_availableTask_valid,
	io_connSS_50_data_availableTask_bits,
	io_connSS_50_data_qOutTask_ready,
	io_connSS_50_data_qOutTask_valid,
	io_connSS_50_data_qOutTask_bits,
	io_connSS_51_ctrl_serveStealReq_valid,
	io_connSS_51_ctrl_serveStealReq_ready,
	io_connSS_51_ctrl_stealReq_valid,
	io_connSS_51_ctrl_stealReq_ready,
	io_connSS_51_data_availableTask_ready,
	io_connSS_51_data_availableTask_valid,
	io_connSS_51_data_availableTask_bits,
	io_connSS_51_data_qOutTask_ready,
	io_connSS_51_data_qOutTask_valid,
	io_connSS_51_data_qOutTask_bits,
	io_connSS_52_ctrl_serveStealReq_valid,
	io_connSS_52_ctrl_serveStealReq_ready,
	io_connSS_52_ctrl_stealReq_valid,
	io_connSS_52_ctrl_stealReq_ready,
	io_connSS_52_data_availableTask_ready,
	io_connSS_52_data_availableTask_valid,
	io_connSS_52_data_availableTask_bits,
	io_connSS_52_data_qOutTask_ready,
	io_connSS_52_data_qOutTask_valid,
	io_connSS_52_data_qOutTask_bits,
	io_connSS_53_ctrl_serveStealReq_valid,
	io_connSS_53_ctrl_serveStealReq_ready,
	io_connSS_53_ctrl_stealReq_valid,
	io_connSS_53_ctrl_stealReq_ready,
	io_connSS_53_data_availableTask_ready,
	io_connSS_53_data_availableTask_valid,
	io_connSS_53_data_availableTask_bits,
	io_connSS_53_data_qOutTask_ready,
	io_connSS_53_data_qOutTask_valid,
	io_connSS_53_data_qOutTask_bits,
	io_connSS_54_ctrl_serveStealReq_valid,
	io_connSS_54_ctrl_serveStealReq_ready,
	io_connSS_54_ctrl_stealReq_valid,
	io_connSS_54_ctrl_stealReq_ready,
	io_connSS_54_data_availableTask_ready,
	io_connSS_54_data_availableTask_valid,
	io_connSS_54_data_availableTask_bits,
	io_connSS_54_data_qOutTask_ready,
	io_connSS_54_data_qOutTask_valid,
	io_connSS_54_data_qOutTask_bits,
	io_connSS_55_ctrl_serveStealReq_valid,
	io_connSS_55_ctrl_serveStealReq_ready,
	io_connSS_55_ctrl_stealReq_valid,
	io_connSS_55_ctrl_stealReq_ready,
	io_connSS_55_data_availableTask_ready,
	io_connSS_55_data_availableTask_valid,
	io_connSS_55_data_availableTask_bits,
	io_connSS_55_data_qOutTask_ready,
	io_connSS_55_data_qOutTask_valid,
	io_connSS_55_data_qOutTask_bits,
	io_connSS_56_ctrl_serveStealReq_valid,
	io_connSS_56_ctrl_serveStealReq_ready,
	io_connSS_56_ctrl_stealReq_valid,
	io_connSS_56_ctrl_stealReq_ready,
	io_connSS_56_data_availableTask_ready,
	io_connSS_56_data_availableTask_valid,
	io_connSS_56_data_availableTask_bits,
	io_connSS_56_data_qOutTask_ready,
	io_connSS_56_data_qOutTask_valid,
	io_connSS_56_data_qOutTask_bits,
	io_connSS_57_ctrl_serveStealReq_valid,
	io_connSS_57_ctrl_serveStealReq_ready,
	io_connSS_57_ctrl_stealReq_valid,
	io_connSS_57_ctrl_stealReq_ready,
	io_connSS_57_data_availableTask_ready,
	io_connSS_57_data_availableTask_valid,
	io_connSS_57_data_availableTask_bits,
	io_connSS_57_data_qOutTask_ready,
	io_connSS_57_data_qOutTask_valid,
	io_connSS_57_data_qOutTask_bits,
	io_connSS_58_ctrl_serveStealReq_valid,
	io_connSS_58_ctrl_serveStealReq_ready,
	io_connSS_58_ctrl_stealReq_valid,
	io_connSS_58_ctrl_stealReq_ready,
	io_connSS_58_data_availableTask_ready,
	io_connSS_58_data_availableTask_valid,
	io_connSS_58_data_availableTask_bits,
	io_connSS_58_data_qOutTask_ready,
	io_connSS_58_data_qOutTask_valid,
	io_connSS_58_data_qOutTask_bits,
	io_connSS_59_ctrl_serveStealReq_valid,
	io_connSS_59_ctrl_serveStealReq_ready,
	io_connSS_59_ctrl_stealReq_valid,
	io_connSS_59_ctrl_stealReq_ready,
	io_connSS_59_data_availableTask_ready,
	io_connSS_59_data_availableTask_valid,
	io_connSS_59_data_availableTask_bits,
	io_connSS_59_data_qOutTask_ready,
	io_connSS_59_data_qOutTask_valid,
	io_connSS_59_data_qOutTask_bits,
	io_connSS_60_ctrl_serveStealReq_valid,
	io_connSS_60_ctrl_serveStealReq_ready,
	io_connSS_60_ctrl_stealReq_valid,
	io_connSS_60_ctrl_stealReq_ready,
	io_connSS_60_data_availableTask_ready,
	io_connSS_60_data_availableTask_valid,
	io_connSS_60_data_availableTask_bits,
	io_connSS_60_data_qOutTask_ready,
	io_connSS_60_data_qOutTask_valid,
	io_connSS_60_data_qOutTask_bits,
	io_connSS_61_ctrl_serveStealReq_valid,
	io_connSS_61_ctrl_serveStealReq_ready,
	io_connSS_61_ctrl_stealReq_valid,
	io_connSS_61_ctrl_stealReq_ready,
	io_connSS_61_data_availableTask_ready,
	io_connSS_61_data_availableTask_valid,
	io_connSS_61_data_availableTask_bits,
	io_connSS_61_data_qOutTask_ready,
	io_connSS_61_data_qOutTask_valid,
	io_connSS_61_data_qOutTask_bits,
	io_connSS_62_ctrl_serveStealReq_valid,
	io_connSS_62_ctrl_serveStealReq_ready,
	io_connSS_62_ctrl_stealReq_valid,
	io_connSS_62_ctrl_stealReq_ready,
	io_connSS_62_data_availableTask_ready,
	io_connSS_62_data_availableTask_valid,
	io_connSS_62_data_availableTask_bits,
	io_connSS_62_data_qOutTask_ready,
	io_connSS_62_data_qOutTask_valid,
	io_connSS_62_data_qOutTask_bits,
	io_connSS_63_ctrl_serveStealReq_valid,
	io_connSS_63_ctrl_serveStealReq_ready,
	io_connSS_63_ctrl_stealReq_valid,
	io_connSS_63_ctrl_stealReq_ready,
	io_connSS_63_data_availableTask_ready,
	io_connSS_63_data_availableTask_valid,
	io_connSS_63_data_availableTask_bits,
	io_connSS_63_data_qOutTask_ready,
	io_connSS_63_data_qOutTask_valid,
	io_connSS_63_data_qOutTask_bits,
	io_connSS_64_ctrl_serveStealReq_valid,
	io_connSS_64_ctrl_serveStealReq_ready,
	io_connSS_64_ctrl_stealReq_valid,
	io_connSS_64_ctrl_stealReq_ready,
	io_connSS_64_data_availableTask_ready,
	io_connSS_64_data_availableTask_valid,
	io_connSS_64_data_availableTask_bits,
	io_connSS_64_data_qOutTask_ready,
	io_connSS_64_data_qOutTask_valid,
	io_connSS_64_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0
);
	input clock;
	input reset;
	input io_connSS_0_ctrl_serveStealReq_valid;
	output wire io_connSS_0_ctrl_serveStealReq_ready;
	input io_connSS_0_data_availableTask_ready;
	output wire io_connSS_0_data_availableTask_valid;
	output wire [255:0] io_connSS_0_data_availableTask_bits;
	output wire io_connSS_0_data_qOutTask_ready;
	input io_connSS_0_data_qOutTask_valid;
	input [255:0] io_connSS_0_data_qOutTask_bits;
	input io_connSS_1_ctrl_serveStealReq_valid;
	output wire io_connSS_1_ctrl_serveStealReq_ready;
	input io_connSS_1_ctrl_stealReq_valid;
	output wire io_connSS_1_ctrl_stealReq_ready;
	input io_connSS_1_data_availableTask_ready;
	output wire io_connSS_1_data_availableTask_valid;
	output wire [255:0] io_connSS_1_data_availableTask_bits;
	output wire io_connSS_1_data_qOutTask_ready;
	input io_connSS_1_data_qOutTask_valid;
	input [255:0] io_connSS_1_data_qOutTask_bits;
	input io_connSS_2_ctrl_serveStealReq_valid;
	output wire io_connSS_2_ctrl_serveStealReq_ready;
	input io_connSS_2_ctrl_stealReq_valid;
	output wire io_connSS_2_ctrl_stealReq_ready;
	input io_connSS_2_data_availableTask_ready;
	output wire io_connSS_2_data_availableTask_valid;
	output wire [255:0] io_connSS_2_data_availableTask_bits;
	output wire io_connSS_2_data_qOutTask_ready;
	input io_connSS_2_data_qOutTask_valid;
	input [255:0] io_connSS_2_data_qOutTask_bits;
	input io_connSS_3_ctrl_serveStealReq_valid;
	output wire io_connSS_3_ctrl_serveStealReq_ready;
	input io_connSS_3_ctrl_stealReq_valid;
	output wire io_connSS_3_ctrl_stealReq_ready;
	input io_connSS_3_data_availableTask_ready;
	output wire io_connSS_3_data_availableTask_valid;
	output wire [255:0] io_connSS_3_data_availableTask_bits;
	output wire io_connSS_3_data_qOutTask_ready;
	input io_connSS_3_data_qOutTask_valid;
	input [255:0] io_connSS_3_data_qOutTask_bits;
	input io_connSS_4_ctrl_serveStealReq_valid;
	output wire io_connSS_4_ctrl_serveStealReq_ready;
	input io_connSS_4_ctrl_stealReq_valid;
	output wire io_connSS_4_ctrl_stealReq_ready;
	input io_connSS_4_data_availableTask_ready;
	output wire io_connSS_4_data_availableTask_valid;
	output wire [255:0] io_connSS_4_data_availableTask_bits;
	output wire io_connSS_4_data_qOutTask_ready;
	input io_connSS_4_data_qOutTask_valid;
	input [255:0] io_connSS_4_data_qOutTask_bits;
	input io_connSS_5_ctrl_serveStealReq_valid;
	output wire io_connSS_5_ctrl_serveStealReq_ready;
	input io_connSS_5_ctrl_stealReq_valid;
	output wire io_connSS_5_ctrl_stealReq_ready;
	input io_connSS_5_data_availableTask_ready;
	output wire io_connSS_5_data_availableTask_valid;
	output wire [255:0] io_connSS_5_data_availableTask_bits;
	output wire io_connSS_5_data_qOutTask_ready;
	input io_connSS_5_data_qOutTask_valid;
	input [255:0] io_connSS_5_data_qOutTask_bits;
	input io_connSS_6_ctrl_serveStealReq_valid;
	output wire io_connSS_6_ctrl_serveStealReq_ready;
	input io_connSS_6_ctrl_stealReq_valid;
	output wire io_connSS_6_ctrl_stealReq_ready;
	input io_connSS_6_data_availableTask_ready;
	output wire io_connSS_6_data_availableTask_valid;
	output wire [255:0] io_connSS_6_data_availableTask_bits;
	output wire io_connSS_6_data_qOutTask_ready;
	input io_connSS_6_data_qOutTask_valid;
	input [255:0] io_connSS_6_data_qOutTask_bits;
	input io_connSS_7_ctrl_serveStealReq_valid;
	output wire io_connSS_7_ctrl_serveStealReq_ready;
	input io_connSS_7_ctrl_stealReq_valid;
	output wire io_connSS_7_ctrl_stealReq_ready;
	input io_connSS_7_data_availableTask_ready;
	output wire io_connSS_7_data_availableTask_valid;
	output wire [255:0] io_connSS_7_data_availableTask_bits;
	output wire io_connSS_7_data_qOutTask_ready;
	input io_connSS_7_data_qOutTask_valid;
	input [255:0] io_connSS_7_data_qOutTask_bits;
	input io_connSS_8_ctrl_serveStealReq_valid;
	output wire io_connSS_8_ctrl_serveStealReq_ready;
	input io_connSS_8_ctrl_stealReq_valid;
	output wire io_connSS_8_ctrl_stealReq_ready;
	input io_connSS_8_data_availableTask_ready;
	output wire io_connSS_8_data_availableTask_valid;
	output wire [255:0] io_connSS_8_data_availableTask_bits;
	output wire io_connSS_8_data_qOutTask_ready;
	input io_connSS_8_data_qOutTask_valid;
	input [255:0] io_connSS_8_data_qOutTask_bits;
	input io_connSS_9_ctrl_serveStealReq_valid;
	output wire io_connSS_9_ctrl_serveStealReq_ready;
	input io_connSS_9_ctrl_stealReq_valid;
	output wire io_connSS_9_ctrl_stealReq_ready;
	input io_connSS_9_data_availableTask_ready;
	output wire io_connSS_9_data_availableTask_valid;
	output wire [255:0] io_connSS_9_data_availableTask_bits;
	output wire io_connSS_9_data_qOutTask_ready;
	input io_connSS_9_data_qOutTask_valid;
	input [255:0] io_connSS_9_data_qOutTask_bits;
	input io_connSS_10_ctrl_serveStealReq_valid;
	output wire io_connSS_10_ctrl_serveStealReq_ready;
	input io_connSS_10_ctrl_stealReq_valid;
	output wire io_connSS_10_ctrl_stealReq_ready;
	input io_connSS_10_data_availableTask_ready;
	output wire io_connSS_10_data_availableTask_valid;
	output wire [255:0] io_connSS_10_data_availableTask_bits;
	output wire io_connSS_10_data_qOutTask_ready;
	input io_connSS_10_data_qOutTask_valid;
	input [255:0] io_connSS_10_data_qOutTask_bits;
	input io_connSS_11_ctrl_serveStealReq_valid;
	output wire io_connSS_11_ctrl_serveStealReq_ready;
	input io_connSS_11_ctrl_stealReq_valid;
	output wire io_connSS_11_ctrl_stealReq_ready;
	input io_connSS_11_data_availableTask_ready;
	output wire io_connSS_11_data_availableTask_valid;
	output wire [255:0] io_connSS_11_data_availableTask_bits;
	output wire io_connSS_11_data_qOutTask_ready;
	input io_connSS_11_data_qOutTask_valid;
	input [255:0] io_connSS_11_data_qOutTask_bits;
	input io_connSS_12_ctrl_serveStealReq_valid;
	output wire io_connSS_12_ctrl_serveStealReq_ready;
	input io_connSS_12_ctrl_stealReq_valid;
	output wire io_connSS_12_ctrl_stealReq_ready;
	input io_connSS_12_data_availableTask_ready;
	output wire io_connSS_12_data_availableTask_valid;
	output wire [255:0] io_connSS_12_data_availableTask_bits;
	output wire io_connSS_12_data_qOutTask_ready;
	input io_connSS_12_data_qOutTask_valid;
	input [255:0] io_connSS_12_data_qOutTask_bits;
	input io_connSS_13_ctrl_serveStealReq_valid;
	output wire io_connSS_13_ctrl_serveStealReq_ready;
	input io_connSS_13_ctrl_stealReq_valid;
	output wire io_connSS_13_ctrl_stealReq_ready;
	input io_connSS_13_data_availableTask_ready;
	output wire io_connSS_13_data_availableTask_valid;
	output wire [255:0] io_connSS_13_data_availableTask_bits;
	output wire io_connSS_13_data_qOutTask_ready;
	input io_connSS_13_data_qOutTask_valid;
	input [255:0] io_connSS_13_data_qOutTask_bits;
	input io_connSS_14_ctrl_serveStealReq_valid;
	output wire io_connSS_14_ctrl_serveStealReq_ready;
	input io_connSS_14_ctrl_stealReq_valid;
	output wire io_connSS_14_ctrl_stealReq_ready;
	input io_connSS_14_data_availableTask_ready;
	output wire io_connSS_14_data_availableTask_valid;
	output wire [255:0] io_connSS_14_data_availableTask_bits;
	output wire io_connSS_14_data_qOutTask_ready;
	input io_connSS_14_data_qOutTask_valid;
	input [255:0] io_connSS_14_data_qOutTask_bits;
	input io_connSS_15_ctrl_serveStealReq_valid;
	output wire io_connSS_15_ctrl_serveStealReq_ready;
	input io_connSS_15_ctrl_stealReq_valid;
	output wire io_connSS_15_ctrl_stealReq_ready;
	input io_connSS_15_data_availableTask_ready;
	output wire io_connSS_15_data_availableTask_valid;
	output wire [255:0] io_connSS_15_data_availableTask_bits;
	output wire io_connSS_15_data_qOutTask_ready;
	input io_connSS_15_data_qOutTask_valid;
	input [255:0] io_connSS_15_data_qOutTask_bits;
	input io_connSS_16_ctrl_serveStealReq_valid;
	output wire io_connSS_16_ctrl_serveStealReq_ready;
	input io_connSS_16_ctrl_stealReq_valid;
	output wire io_connSS_16_ctrl_stealReq_ready;
	input io_connSS_16_data_availableTask_ready;
	output wire io_connSS_16_data_availableTask_valid;
	output wire [255:0] io_connSS_16_data_availableTask_bits;
	output wire io_connSS_16_data_qOutTask_ready;
	input io_connSS_16_data_qOutTask_valid;
	input [255:0] io_connSS_16_data_qOutTask_bits;
	input io_connSS_17_ctrl_serveStealReq_valid;
	output wire io_connSS_17_ctrl_serveStealReq_ready;
	input io_connSS_17_ctrl_stealReq_valid;
	output wire io_connSS_17_ctrl_stealReq_ready;
	input io_connSS_17_data_availableTask_ready;
	output wire io_connSS_17_data_availableTask_valid;
	output wire [255:0] io_connSS_17_data_availableTask_bits;
	output wire io_connSS_17_data_qOutTask_ready;
	input io_connSS_17_data_qOutTask_valid;
	input [255:0] io_connSS_17_data_qOutTask_bits;
	input io_connSS_18_ctrl_serveStealReq_valid;
	output wire io_connSS_18_ctrl_serveStealReq_ready;
	input io_connSS_18_ctrl_stealReq_valid;
	output wire io_connSS_18_ctrl_stealReq_ready;
	input io_connSS_18_data_availableTask_ready;
	output wire io_connSS_18_data_availableTask_valid;
	output wire [255:0] io_connSS_18_data_availableTask_bits;
	output wire io_connSS_18_data_qOutTask_ready;
	input io_connSS_18_data_qOutTask_valid;
	input [255:0] io_connSS_18_data_qOutTask_bits;
	input io_connSS_19_ctrl_serveStealReq_valid;
	output wire io_connSS_19_ctrl_serveStealReq_ready;
	input io_connSS_19_ctrl_stealReq_valid;
	output wire io_connSS_19_ctrl_stealReq_ready;
	input io_connSS_19_data_availableTask_ready;
	output wire io_connSS_19_data_availableTask_valid;
	output wire [255:0] io_connSS_19_data_availableTask_bits;
	output wire io_connSS_19_data_qOutTask_ready;
	input io_connSS_19_data_qOutTask_valid;
	input [255:0] io_connSS_19_data_qOutTask_bits;
	input io_connSS_20_ctrl_serveStealReq_valid;
	output wire io_connSS_20_ctrl_serveStealReq_ready;
	input io_connSS_20_ctrl_stealReq_valid;
	output wire io_connSS_20_ctrl_stealReq_ready;
	input io_connSS_20_data_availableTask_ready;
	output wire io_connSS_20_data_availableTask_valid;
	output wire [255:0] io_connSS_20_data_availableTask_bits;
	output wire io_connSS_20_data_qOutTask_ready;
	input io_connSS_20_data_qOutTask_valid;
	input [255:0] io_connSS_20_data_qOutTask_bits;
	input io_connSS_21_ctrl_serveStealReq_valid;
	output wire io_connSS_21_ctrl_serveStealReq_ready;
	input io_connSS_21_ctrl_stealReq_valid;
	output wire io_connSS_21_ctrl_stealReq_ready;
	input io_connSS_21_data_availableTask_ready;
	output wire io_connSS_21_data_availableTask_valid;
	output wire [255:0] io_connSS_21_data_availableTask_bits;
	output wire io_connSS_21_data_qOutTask_ready;
	input io_connSS_21_data_qOutTask_valid;
	input [255:0] io_connSS_21_data_qOutTask_bits;
	input io_connSS_22_ctrl_serveStealReq_valid;
	output wire io_connSS_22_ctrl_serveStealReq_ready;
	input io_connSS_22_ctrl_stealReq_valid;
	output wire io_connSS_22_ctrl_stealReq_ready;
	input io_connSS_22_data_availableTask_ready;
	output wire io_connSS_22_data_availableTask_valid;
	output wire [255:0] io_connSS_22_data_availableTask_bits;
	output wire io_connSS_22_data_qOutTask_ready;
	input io_connSS_22_data_qOutTask_valid;
	input [255:0] io_connSS_22_data_qOutTask_bits;
	input io_connSS_23_ctrl_serveStealReq_valid;
	output wire io_connSS_23_ctrl_serveStealReq_ready;
	input io_connSS_23_ctrl_stealReq_valid;
	output wire io_connSS_23_ctrl_stealReq_ready;
	input io_connSS_23_data_availableTask_ready;
	output wire io_connSS_23_data_availableTask_valid;
	output wire [255:0] io_connSS_23_data_availableTask_bits;
	output wire io_connSS_23_data_qOutTask_ready;
	input io_connSS_23_data_qOutTask_valid;
	input [255:0] io_connSS_23_data_qOutTask_bits;
	input io_connSS_24_ctrl_serveStealReq_valid;
	output wire io_connSS_24_ctrl_serveStealReq_ready;
	input io_connSS_24_ctrl_stealReq_valid;
	output wire io_connSS_24_ctrl_stealReq_ready;
	input io_connSS_24_data_availableTask_ready;
	output wire io_connSS_24_data_availableTask_valid;
	output wire [255:0] io_connSS_24_data_availableTask_bits;
	output wire io_connSS_24_data_qOutTask_ready;
	input io_connSS_24_data_qOutTask_valid;
	input [255:0] io_connSS_24_data_qOutTask_bits;
	input io_connSS_25_ctrl_serveStealReq_valid;
	output wire io_connSS_25_ctrl_serveStealReq_ready;
	input io_connSS_25_ctrl_stealReq_valid;
	output wire io_connSS_25_ctrl_stealReq_ready;
	input io_connSS_25_data_availableTask_ready;
	output wire io_connSS_25_data_availableTask_valid;
	output wire [255:0] io_connSS_25_data_availableTask_bits;
	output wire io_connSS_25_data_qOutTask_ready;
	input io_connSS_25_data_qOutTask_valid;
	input [255:0] io_connSS_25_data_qOutTask_bits;
	input io_connSS_26_ctrl_serveStealReq_valid;
	output wire io_connSS_26_ctrl_serveStealReq_ready;
	input io_connSS_26_ctrl_stealReq_valid;
	output wire io_connSS_26_ctrl_stealReq_ready;
	input io_connSS_26_data_availableTask_ready;
	output wire io_connSS_26_data_availableTask_valid;
	output wire [255:0] io_connSS_26_data_availableTask_bits;
	output wire io_connSS_26_data_qOutTask_ready;
	input io_connSS_26_data_qOutTask_valid;
	input [255:0] io_connSS_26_data_qOutTask_bits;
	input io_connSS_27_ctrl_serveStealReq_valid;
	output wire io_connSS_27_ctrl_serveStealReq_ready;
	input io_connSS_27_ctrl_stealReq_valid;
	output wire io_connSS_27_ctrl_stealReq_ready;
	input io_connSS_27_data_availableTask_ready;
	output wire io_connSS_27_data_availableTask_valid;
	output wire [255:0] io_connSS_27_data_availableTask_bits;
	output wire io_connSS_27_data_qOutTask_ready;
	input io_connSS_27_data_qOutTask_valid;
	input [255:0] io_connSS_27_data_qOutTask_bits;
	input io_connSS_28_ctrl_serveStealReq_valid;
	output wire io_connSS_28_ctrl_serveStealReq_ready;
	input io_connSS_28_ctrl_stealReq_valid;
	output wire io_connSS_28_ctrl_stealReq_ready;
	input io_connSS_28_data_availableTask_ready;
	output wire io_connSS_28_data_availableTask_valid;
	output wire [255:0] io_connSS_28_data_availableTask_bits;
	output wire io_connSS_28_data_qOutTask_ready;
	input io_connSS_28_data_qOutTask_valid;
	input [255:0] io_connSS_28_data_qOutTask_bits;
	input io_connSS_29_ctrl_serveStealReq_valid;
	output wire io_connSS_29_ctrl_serveStealReq_ready;
	input io_connSS_29_ctrl_stealReq_valid;
	output wire io_connSS_29_ctrl_stealReq_ready;
	input io_connSS_29_data_availableTask_ready;
	output wire io_connSS_29_data_availableTask_valid;
	output wire [255:0] io_connSS_29_data_availableTask_bits;
	output wire io_connSS_29_data_qOutTask_ready;
	input io_connSS_29_data_qOutTask_valid;
	input [255:0] io_connSS_29_data_qOutTask_bits;
	input io_connSS_30_ctrl_serveStealReq_valid;
	output wire io_connSS_30_ctrl_serveStealReq_ready;
	input io_connSS_30_ctrl_stealReq_valid;
	output wire io_connSS_30_ctrl_stealReq_ready;
	input io_connSS_30_data_availableTask_ready;
	output wire io_connSS_30_data_availableTask_valid;
	output wire [255:0] io_connSS_30_data_availableTask_bits;
	output wire io_connSS_30_data_qOutTask_ready;
	input io_connSS_30_data_qOutTask_valid;
	input [255:0] io_connSS_30_data_qOutTask_bits;
	input io_connSS_31_ctrl_serveStealReq_valid;
	output wire io_connSS_31_ctrl_serveStealReq_ready;
	input io_connSS_31_ctrl_stealReq_valid;
	output wire io_connSS_31_ctrl_stealReq_ready;
	input io_connSS_31_data_availableTask_ready;
	output wire io_connSS_31_data_availableTask_valid;
	output wire [255:0] io_connSS_31_data_availableTask_bits;
	output wire io_connSS_31_data_qOutTask_ready;
	input io_connSS_31_data_qOutTask_valid;
	input [255:0] io_connSS_31_data_qOutTask_bits;
	input io_connSS_32_ctrl_serveStealReq_valid;
	output wire io_connSS_32_ctrl_serveStealReq_ready;
	input io_connSS_32_ctrl_stealReq_valid;
	output wire io_connSS_32_ctrl_stealReq_ready;
	input io_connSS_32_data_availableTask_ready;
	output wire io_connSS_32_data_availableTask_valid;
	output wire [255:0] io_connSS_32_data_availableTask_bits;
	output wire io_connSS_32_data_qOutTask_ready;
	input io_connSS_32_data_qOutTask_valid;
	input [255:0] io_connSS_32_data_qOutTask_bits;
	input io_connSS_33_ctrl_serveStealReq_valid;
	output wire io_connSS_33_ctrl_serveStealReq_ready;
	input io_connSS_33_ctrl_stealReq_valid;
	output wire io_connSS_33_ctrl_stealReq_ready;
	input io_connSS_33_data_availableTask_ready;
	output wire io_connSS_33_data_availableTask_valid;
	output wire [255:0] io_connSS_33_data_availableTask_bits;
	output wire io_connSS_33_data_qOutTask_ready;
	input io_connSS_33_data_qOutTask_valid;
	input [255:0] io_connSS_33_data_qOutTask_bits;
	input io_connSS_34_ctrl_serveStealReq_valid;
	output wire io_connSS_34_ctrl_serveStealReq_ready;
	input io_connSS_34_ctrl_stealReq_valid;
	output wire io_connSS_34_ctrl_stealReq_ready;
	input io_connSS_34_data_availableTask_ready;
	output wire io_connSS_34_data_availableTask_valid;
	output wire [255:0] io_connSS_34_data_availableTask_bits;
	output wire io_connSS_34_data_qOutTask_ready;
	input io_connSS_34_data_qOutTask_valid;
	input [255:0] io_connSS_34_data_qOutTask_bits;
	input io_connSS_35_ctrl_serveStealReq_valid;
	output wire io_connSS_35_ctrl_serveStealReq_ready;
	input io_connSS_35_ctrl_stealReq_valid;
	output wire io_connSS_35_ctrl_stealReq_ready;
	input io_connSS_35_data_availableTask_ready;
	output wire io_connSS_35_data_availableTask_valid;
	output wire [255:0] io_connSS_35_data_availableTask_bits;
	output wire io_connSS_35_data_qOutTask_ready;
	input io_connSS_35_data_qOutTask_valid;
	input [255:0] io_connSS_35_data_qOutTask_bits;
	input io_connSS_36_ctrl_serveStealReq_valid;
	output wire io_connSS_36_ctrl_serveStealReq_ready;
	input io_connSS_36_ctrl_stealReq_valid;
	output wire io_connSS_36_ctrl_stealReq_ready;
	input io_connSS_36_data_availableTask_ready;
	output wire io_connSS_36_data_availableTask_valid;
	output wire [255:0] io_connSS_36_data_availableTask_bits;
	output wire io_connSS_36_data_qOutTask_ready;
	input io_connSS_36_data_qOutTask_valid;
	input [255:0] io_connSS_36_data_qOutTask_bits;
	input io_connSS_37_ctrl_serveStealReq_valid;
	output wire io_connSS_37_ctrl_serveStealReq_ready;
	input io_connSS_37_ctrl_stealReq_valid;
	output wire io_connSS_37_ctrl_stealReq_ready;
	input io_connSS_37_data_availableTask_ready;
	output wire io_connSS_37_data_availableTask_valid;
	output wire [255:0] io_connSS_37_data_availableTask_bits;
	output wire io_connSS_37_data_qOutTask_ready;
	input io_connSS_37_data_qOutTask_valid;
	input [255:0] io_connSS_37_data_qOutTask_bits;
	input io_connSS_38_ctrl_serveStealReq_valid;
	output wire io_connSS_38_ctrl_serveStealReq_ready;
	input io_connSS_38_ctrl_stealReq_valid;
	output wire io_connSS_38_ctrl_stealReq_ready;
	input io_connSS_38_data_availableTask_ready;
	output wire io_connSS_38_data_availableTask_valid;
	output wire [255:0] io_connSS_38_data_availableTask_bits;
	output wire io_connSS_38_data_qOutTask_ready;
	input io_connSS_38_data_qOutTask_valid;
	input [255:0] io_connSS_38_data_qOutTask_bits;
	input io_connSS_39_ctrl_serveStealReq_valid;
	output wire io_connSS_39_ctrl_serveStealReq_ready;
	input io_connSS_39_ctrl_stealReq_valid;
	output wire io_connSS_39_ctrl_stealReq_ready;
	input io_connSS_39_data_availableTask_ready;
	output wire io_connSS_39_data_availableTask_valid;
	output wire [255:0] io_connSS_39_data_availableTask_bits;
	output wire io_connSS_39_data_qOutTask_ready;
	input io_connSS_39_data_qOutTask_valid;
	input [255:0] io_connSS_39_data_qOutTask_bits;
	input io_connSS_40_ctrl_serveStealReq_valid;
	output wire io_connSS_40_ctrl_serveStealReq_ready;
	input io_connSS_40_ctrl_stealReq_valid;
	output wire io_connSS_40_ctrl_stealReq_ready;
	input io_connSS_40_data_availableTask_ready;
	output wire io_connSS_40_data_availableTask_valid;
	output wire [255:0] io_connSS_40_data_availableTask_bits;
	output wire io_connSS_40_data_qOutTask_ready;
	input io_connSS_40_data_qOutTask_valid;
	input [255:0] io_connSS_40_data_qOutTask_bits;
	input io_connSS_41_ctrl_serveStealReq_valid;
	output wire io_connSS_41_ctrl_serveStealReq_ready;
	input io_connSS_41_ctrl_stealReq_valid;
	output wire io_connSS_41_ctrl_stealReq_ready;
	input io_connSS_41_data_availableTask_ready;
	output wire io_connSS_41_data_availableTask_valid;
	output wire [255:0] io_connSS_41_data_availableTask_bits;
	output wire io_connSS_41_data_qOutTask_ready;
	input io_connSS_41_data_qOutTask_valid;
	input [255:0] io_connSS_41_data_qOutTask_bits;
	input io_connSS_42_ctrl_serveStealReq_valid;
	output wire io_connSS_42_ctrl_serveStealReq_ready;
	input io_connSS_42_ctrl_stealReq_valid;
	output wire io_connSS_42_ctrl_stealReq_ready;
	input io_connSS_42_data_availableTask_ready;
	output wire io_connSS_42_data_availableTask_valid;
	output wire [255:0] io_connSS_42_data_availableTask_bits;
	output wire io_connSS_42_data_qOutTask_ready;
	input io_connSS_42_data_qOutTask_valid;
	input [255:0] io_connSS_42_data_qOutTask_bits;
	input io_connSS_43_ctrl_serveStealReq_valid;
	output wire io_connSS_43_ctrl_serveStealReq_ready;
	input io_connSS_43_ctrl_stealReq_valid;
	output wire io_connSS_43_ctrl_stealReq_ready;
	input io_connSS_43_data_availableTask_ready;
	output wire io_connSS_43_data_availableTask_valid;
	output wire [255:0] io_connSS_43_data_availableTask_bits;
	output wire io_connSS_43_data_qOutTask_ready;
	input io_connSS_43_data_qOutTask_valid;
	input [255:0] io_connSS_43_data_qOutTask_bits;
	input io_connSS_44_ctrl_serveStealReq_valid;
	output wire io_connSS_44_ctrl_serveStealReq_ready;
	input io_connSS_44_ctrl_stealReq_valid;
	output wire io_connSS_44_ctrl_stealReq_ready;
	input io_connSS_44_data_availableTask_ready;
	output wire io_connSS_44_data_availableTask_valid;
	output wire [255:0] io_connSS_44_data_availableTask_bits;
	output wire io_connSS_44_data_qOutTask_ready;
	input io_connSS_44_data_qOutTask_valid;
	input [255:0] io_connSS_44_data_qOutTask_bits;
	input io_connSS_45_ctrl_serveStealReq_valid;
	output wire io_connSS_45_ctrl_serveStealReq_ready;
	input io_connSS_45_ctrl_stealReq_valid;
	output wire io_connSS_45_ctrl_stealReq_ready;
	input io_connSS_45_data_availableTask_ready;
	output wire io_connSS_45_data_availableTask_valid;
	output wire [255:0] io_connSS_45_data_availableTask_bits;
	output wire io_connSS_45_data_qOutTask_ready;
	input io_connSS_45_data_qOutTask_valid;
	input [255:0] io_connSS_45_data_qOutTask_bits;
	input io_connSS_46_ctrl_serveStealReq_valid;
	output wire io_connSS_46_ctrl_serveStealReq_ready;
	input io_connSS_46_ctrl_stealReq_valid;
	output wire io_connSS_46_ctrl_stealReq_ready;
	input io_connSS_46_data_availableTask_ready;
	output wire io_connSS_46_data_availableTask_valid;
	output wire [255:0] io_connSS_46_data_availableTask_bits;
	output wire io_connSS_46_data_qOutTask_ready;
	input io_connSS_46_data_qOutTask_valid;
	input [255:0] io_connSS_46_data_qOutTask_bits;
	input io_connSS_47_ctrl_serveStealReq_valid;
	output wire io_connSS_47_ctrl_serveStealReq_ready;
	input io_connSS_47_ctrl_stealReq_valid;
	output wire io_connSS_47_ctrl_stealReq_ready;
	input io_connSS_47_data_availableTask_ready;
	output wire io_connSS_47_data_availableTask_valid;
	output wire [255:0] io_connSS_47_data_availableTask_bits;
	output wire io_connSS_47_data_qOutTask_ready;
	input io_connSS_47_data_qOutTask_valid;
	input [255:0] io_connSS_47_data_qOutTask_bits;
	input io_connSS_48_ctrl_serveStealReq_valid;
	output wire io_connSS_48_ctrl_serveStealReq_ready;
	input io_connSS_48_ctrl_stealReq_valid;
	output wire io_connSS_48_ctrl_stealReq_ready;
	input io_connSS_48_data_availableTask_ready;
	output wire io_connSS_48_data_availableTask_valid;
	output wire [255:0] io_connSS_48_data_availableTask_bits;
	output wire io_connSS_48_data_qOutTask_ready;
	input io_connSS_48_data_qOutTask_valid;
	input [255:0] io_connSS_48_data_qOutTask_bits;
	input io_connSS_49_ctrl_serveStealReq_valid;
	output wire io_connSS_49_ctrl_serveStealReq_ready;
	input io_connSS_49_ctrl_stealReq_valid;
	output wire io_connSS_49_ctrl_stealReq_ready;
	input io_connSS_49_data_availableTask_ready;
	output wire io_connSS_49_data_availableTask_valid;
	output wire [255:0] io_connSS_49_data_availableTask_bits;
	output wire io_connSS_49_data_qOutTask_ready;
	input io_connSS_49_data_qOutTask_valid;
	input [255:0] io_connSS_49_data_qOutTask_bits;
	input io_connSS_50_ctrl_serveStealReq_valid;
	output wire io_connSS_50_ctrl_serveStealReq_ready;
	input io_connSS_50_ctrl_stealReq_valid;
	output wire io_connSS_50_ctrl_stealReq_ready;
	input io_connSS_50_data_availableTask_ready;
	output wire io_connSS_50_data_availableTask_valid;
	output wire [255:0] io_connSS_50_data_availableTask_bits;
	output wire io_connSS_50_data_qOutTask_ready;
	input io_connSS_50_data_qOutTask_valid;
	input [255:0] io_connSS_50_data_qOutTask_bits;
	input io_connSS_51_ctrl_serveStealReq_valid;
	output wire io_connSS_51_ctrl_serveStealReq_ready;
	input io_connSS_51_ctrl_stealReq_valid;
	output wire io_connSS_51_ctrl_stealReq_ready;
	input io_connSS_51_data_availableTask_ready;
	output wire io_connSS_51_data_availableTask_valid;
	output wire [255:0] io_connSS_51_data_availableTask_bits;
	output wire io_connSS_51_data_qOutTask_ready;
	input io_connSS_51_data_qOutTask_valid;
	input [255:0] io_connSS_51_data_qOutTask_bits;
	input io_connSS_52_ctrl_serveStealReq_valid;
	output wire io_connSS_52_ctrl_serveStealReq_ready;
	input io_connSS_52_ctrl_stealReq_valid;
	output wire io_connSS_52_ctrl_stealReq_ready;
	input io_connSS_52_data_availableTask_ready;
	output wire io_connSS_52_data_availableTask_valid;
	output wire [255:0] io_connSS_52_data_availableTask_bits;
	output wire io_connSS_52_data_qOutTask_ready;
	input io_connSS_52_data_qOutTask_valid;
	input [255:0] io_connSS_52_data_qOutTask_bits;
	input io_connSS_53_ctrl_serveStealReq_valid;
	output wire io_connSS_53_ctrl_serveStealReq_ready;
	input io_connSS_53_ctrl_stealReq_valid;
	output wire io_connSS_53_ctrl_stealReq_ready;
	input io_connSS_53_data_availableTask_ready;
	output wire io_connSS_53_data_availableTask_valid;
	output wire [255:0] io_connSS_53_data_availableTask_bits;
	output wire io_connSS_53_data_qOutTask_ready;
	input io_connSS_53_data_qOutTask_valid;
	input [255:0] io_connSS_53_data_qOutTask_bits;
	input io_connSS_54_ctrl_serveStealReq_valid;
	output wire io_connSS_54_ctrl_serveStealReq_ready;
	input io_connSS_54_ctrl_stealReq_valid;
	output wire io_connSS_54_ctrl_stealReq_ready;
	input io_connSS_54_data_availableTask_ready;
	output wire io_connSS_54_data_availableTask_valid;
	output wire [255:0] io_connSS_54_data_availableTask_bits;
	output wire io_connSS_54_data_qOutTask_ready;
	input io_connSS_54_data_qOutTask_valid;
	input [255:0] io_connSS_54_data_qOutTask_bits;
	input io_connSS_55_ctrl_serveStealReq_valid;
	output wire io_connSS_55_ctrl_serveStealReq_ready;
	input io_connSS_55_ctrl_stealReq_valid;
	output wire io_connSS_55_ctrl_stealReq_ready;
	input io_connSS_55_data_availableTask_ready;
	output wire io_connSS_55_data_availableTask_valid;
	output wire [255:0] io_connSS_55_data_availableTask_bits;
	output wire io_connSS_55_data_qOutTask_ready;
	input io_connSS_55_data_qOutTask_valid;
	input [255:0] io_connSS_55_data_qOutTask_bits;
	input io_connSS_56_ctrl_serveStealReq_valid;
	output wire io_connSS_56_ctrl_serveStealReq_ready;
	input io_connSS_56_ctrl_stealReq_valid;
	output wire io_connSS_56_ctrl_stealReq_ready;
	input io_connSS_56_data_availableTask_ready;
	output wire io_connSS_56_data_availableTask_valid;
	output wire [255:0] io_connSS_56_data_availableTask_bits;
	output wire io_connSS_56_data_qOutTask_ready;
	input io_connSS_56_data_qOutTask_valid;
	input [255:0] io_connSS_56_data_qOutTask_bits;
	input io_connSS_57_ctrl_serveStealReq_valid;
	output wire io_connSS_57_ctrl_serveStealReq_ready;
	input io_connSS_57_ctrl_stealReq_valid;
	output wire io_connSS_57_ctrl_stealReq_ready;
	input io_connSS_57_data_availableTask_ready;
	output wire io_connSS_57_data_availableTask_valid;
	output wire [255:0] io_connSS_57_data_availableTask_bits;
	output wire io_connSS_57_data_qOutTask_ready;
	input io_connSS_57_data_qOutTask_valid;
	input [255:0] io_connSS_57_data_qOutTask_bits;
	input io_connSS_58_ctrl_serveStealReq_valid;
	output wire io_connSS_58_ctrl_serveStealReq_ready;
	input io_connSS_58_ctrl_stealReq_valid;
	output wire io_connSS_58_ctrl_stealReq_ready;
	input io_connSS_58_data_availableTask_ready;
	output wire io_connSS_58_data_availableTask_valid;
	output wire [255:0] io_connSS_58_data_availableTask_bits;
	output wire io_connSS_58_data_qOutTask_ready;
	input io_connSS_58_data_qOutTask_valid;
	input [255:0] io_connSS_58_data_qOutTask_bits;
	input io_connSS_59_ctrl_serveStealReq_valid;
	output wire io_connSS_59_ctrl_serveStealReq_ready;
	input io_connSS_59_ctrl_stealReq_valid;
	output wire io_connSS_59_ctrl_stealReq_ready;
	input io_connSS_59_data_availableTask_ready;
	output wire io_connSS_59_data_availableTask_valid;
	output wire [255:0] io_connSS_59_data_availableTask_bits;
	output wire io_connSS_59_data_qOutTask_ready;
	input io_connSS_59_data_qOutTask_valid;
	input [255:0] io_connSS_59_data_qOutTask_bits;
	input io_connSS_60_ctrl_serveStealReq_valid;
	output wire io_connSS_60_ctrl_serveStealReq_ready;
	input io_connSS_60_ctrl_stealReq_valid;
	output wire io_connSS_60_ctrl_stealReq_ready;
	input io_connSS_60_data_availableTask_ready;
	output wire io_connSS_60_data_availableTask_valid;
	output wire [255:0] io_connSS_60_data_availableTask_bits;
	output wire io_connSS_60_data_qOutTask_ready;
	input io_connSS_60_data_qOutTask_valid;
	input [255:0] io_connSS_60_data_qOutTask_bits;
	input io_connSS_61_ctrl_serveStealReq_valid;
	output wire io_connSS_61_ctrl_serveStealReq_ready;
	input io_connSS_61_ctrl_stealReq_valid;
	output wire io_connSS_61_ctrl_stealReq_ready;
	input io_connSS_61_data_availableTask_ready;
	output wire io_connSS_61_data_availableTask_valid;
	output wire [255:0] io_connSS_61_data_availableTask_bits;
	output wire io_connSS_61_data_qOutTask_ready;
	input io_connSS_61_data_qOutTask_valid;
	input [255:0] io_connSS_61_data_qOutTask_bits;
	input io_connSS_62_ctrl_serveStealReq_valid;
	output wire io_connSS_62_ctrl_serveStealReq_ready;
	input io_connSS_62_ctrl_stealReq_valid;
	output wire io_connSS_62_ctrl_stealReq_ready;
	input io_connSS_62_data_availableTask_ready;
	output wire io_connSS_62_data_availableTask_valid;
	output wire [255:0] io_connSS_62_data_availableTask_bits;
	output wire io_connSS_62_data_qOutTask_ready;
	input io_connSS_62_data_qOutTask_valid;
	input [255:0] io_connSS_62_data_qOutTask_bits;
	input io_connSS_63_ctrl_serveStealReq_valid;
	output wire io_connSS_63_ctrl_serveStealReq_ready;
	input io_connSS_63_ctrl_stealReq_valid;
	output wire io_connSS_63_ctrl_stealReq_ready;
	input io_connSS_63_data_availableTask_ready;
	output wire io_connSS_63_data_availableTask_valid;
	output wire [255:0] io_connSS_63_data_availableTask_bits;
	output wire io_connSS_63_data_qOutTask_ready;
	input io_connSS_63_data_qOutTask_valid;
	input [255:0] io_connSS_63_data_qOutTask_bits;
	input io_connSS_64_ctrl_serveStealReq_valid;
	output wire io_connSS_64_ctrl_serveStealReq_ready;
	input io_connSS_64_ctrl_stealReq_valid;
	output wire io_connSS_64_ctrl_stealReq_ready;
	input io_connSS_64_data_availableTask_ready;
	output wire io_connSS_64_data_availableTask_valid;
	output wire [255:0] io_connSS_64_data_availableTask_bits;
	output wire io_connSS_64_data_qOutTask_ready;
	input io_connSS_64_data_qOutTask_valid;
	input [255:0] io_connSS_64_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	wire _ctrlunits_64_io_reqTaskOut;
	wire _ctrlunits_63_io_reqTaskOut;
	wire _ctrlunits_62_io_reqTaskOut;
	wire _ctrlunits_61_io_reqTaskOut;
	wire _ctrlunits_60_io_reqTaskOut;
	wire _ctrlunits_59_io_reqTaskOut;
	wire _ctrlunits_58_io_reqTaskOut;
	wire _ctrlunits_57_io_reqTaskOut;
	wire _ctrlunits_56_io_reqTaskOut;
	wire _ctrlunits_55_io_reqTaskOut;
	wire _ctrlunits_54_io_reqTaskOut;
	wire _ctrlunits_53_io_reqTaskOut;
	wire _ctrlunits_52_io_reqTaskOut;
	wire _ctrlunits_51_io_reqTaskOut;
	wire _ctrlunits_50_io_reqTaskOut;
	wire _ctrlunits_49_io_reqTaskOut;
	wire _ctrlunits_48_io_reqTaskOut;
	wire _ctrlunits_47_io_reqTaskOut;
	wire _ctrlunits_46_io_reqTaskOut;
	wire _ctrlunits_45_io_reqTaskOut;
	wire _ctrlunits_44_io_reqTaskOut;
	wire _ctrlunits_43_io_reqTaskOut;
	wire _ctrlunits_42_io_reqTaskOut;
	wire _ctrlunits_41_io_reqTaskOut;
	wire _ctrlunits_40_io_reqTaskOut;
	wire _ctrlunits_39_io_reqTaskOut;
	wire _ctrlunits_38_io_reqTaskOut;
	wire _ctrlunits_37_io_reqTaskOut;
	wire _ctrlunits_36_io_reqTaskOut;
	wire _ctrlunits_35_io_reqTaskOut;
	wire _ctrlunits_34_io_reqTaskOut;
	wire _ctrlunits_33_io_reqTaskOut;
	wire _ctrlunits_32_io_reqTaskOut;
	wire _ctrlunits_31_io_reqTaskOut;
	wire _ctrlunits_30_io_reqTaskOut;
	wire _ctrlunits_29_io_reqTaskOut;
	wire _ctrlunits_28_io_reqTaskOut;
	wire _ctrlunits_27_io_reqTaskOut;
	wire _ctrlunits_26_io_reqTaskOut;
	wire _ctrlunits_25_io_reqTaskOut;
	wire _ctrlunits_24_io_reqTaskOut;
	wire _ctrlunits_23_io_reqTaskOut;
	wire _ctrlunits_22_io_reqTaskOut;
	wire _ctrlunits_21_io_reqTaskOut;
	wire _ctrlunits_20_io_reqTaskOut;
	wire _ctrlunits_19_io_reqTaskOut;
	wire _ctrlunits_18_io_reqTaskOut;
	wire _ctrlunits_17_io_reqTaskOut;
	wire _ctrlunits_16_io_reqTaskOut;
	wire _ctrlunits_15_io_reqTaskOut;
	wire _ctrlunits_14_io_reqTaskOut;
	wire _ctrlunits_13_io_reqTaskOut;
	wire _ctrlunits_12_io_reqTaskOut;
	wire _ctrlunits_11_io_reqTaskOut;
	wire _ctrlunits_10_io_reqTaskOut;
	wire _ctrlunits_9_io_reqTaskOut;
	wire _ctrlunits_8_io_reqTaskOut;
	wire _ctrlunits_7_io_reqTaskOut;
	wire _ctrlunits_6_io_reqTaskOut;
	wire _ctrlunits_5_io_reqTaskOut;
	wire _ctrlunits_4_io_reqTaskOut;
	wire _ctrlunits_3_io_reqTaskOut;
	wire _ctrlunits_2_io_reqTaskOut;
	wire _ctrlunits_1_io_reqTaskOut;
	wire _ctrlunits_0_io_reqTaskOut;
	wire [255:0] _dataUnits_64_io_taskOut;
	wire _dataUnits_64_io_validOut;
	wire [255:0] _dataUnits_63_io_taskOut;
	wire _dataUnits_63_io_validOut;
	wire [255:0] _dataUnits_62_io_taskOut;
	wire _dataUnits_62_io_validOut;
	wire [255:0] _dataUnits_61_io_taskOut;
	wire _dataUnits_61_io_validOut;
	wire [255:0] _dataUnits_60_io_taskOut;
	wire _dataUnits_60_io_validOut;
	wire [255:0] _dataUnits_59_io_taskOut;
	wire _dataUnits_59_io_validOut;
	wire [255:0] _dataUnits_58_io_taskOut;
	wire _dataUnits_58_io_validOut;
	wire [255:0] _dataUnits_57_io_taskOut;
	wire _dataUnits_57_io_validOut;
	wire [255:0] _dataUnits_56_io_taskOut;
	wire _dataUnits_56_io_validOut;
	wire [255:0] _dataUnits_55_io_taskOut;
	wire _dataUnits_55_io_validOut;
	wire [255:0] _dataUnits_54_io_taskOut;
	wire _dataUnits_54_io_validOut;
	wire [255:0] _dataUnits_53_io_taskOut;
	wire _dataUnits_53_io_validOut;
	wire [255:0] _dataUnits_52_io_taskOut;
	wire _dataUnits_52_io_validOut;
	wire [255:0] _dataUnits_51_io_taskOut;
	wire _dataUnits_51_io_validOut;
	wire [255:0] _dataUnits_50_io_taskOut;
	wire _dataUnits_50_io_validOut;
	wire [255:0] _dataUnits_49_io_taskOut;
	wire _dataUnits_49_io_validOut;
	wire [255:0] _dataUnits_48_io_taskOut;
	wire _dataUnits_48_io_validOut;
	wire [255:0] _dataUnits_47_io_taskOut;
	wire _dataUnits_47_io_validOut;
	wire [255:0] _dataUnits_46_io_taskOut;
	wire _dataUnits_46_io_validOut;
	wire [255:0] _dataUnits_45_io_taskOut;
	wire _dataUnits_45_io_validOut;
	wire [255:0] _dataUnits_44_io_taskOut;
	wire _dataUnits_44_io_validOut;
	wire [255:0] _dataUnits_43_io_taskOut;
	wire _dataUnits_43_io_validOut;
	wire [255:0] _dataUnits_42_io_taskOut;
	wire _dataUnits_42_io_validOut;
	wire [255:0] _dataUnits_41_io_taskOut;
	wire _dataUnits_41_io_validOut;
	wire [255:0] _dataUnits_40_io_taskOut;
	wire _dataUnits_40_io_validOut;
	wire [255:0] _dataUnits_39_io_taskOut;
	wire _dataUnits_39_io_validOut;
	wire [255:0] _dataUnits_38_io_taskOut;
	wire _dataUnits_38_io_validOut;
	wire [255:0] _dataUnits_37_io_taskOut;
	wire _dataUnits_37_io_validOut;
	wire [255:0] _dataUnits_36_io_taskOut;
	wire _dataUnits_36_io_validOut;
	wire [255:0] _dataUnits_35_io_taskOut;
	wire _dataUnits_35_io_validOut;
	wire [255:0] _dataUnits_34_io_taskOut;
	wire _dataUnits_34_io_validOut;
	wire [255:0] _dataUnits_33_io_taskOut;
	wire _dataUnits_33_io_validOut;
	wire [255:0] _dataUnits_32_io_taskOut;
	wire _dataUnits_32_io_validOut;
	wire [255:0] _dataUnits_31_io_taskOut;
	wire _dataUnits_31_io_validOut;
	wire [255:0] _dataUnits_30_io_taskOut;
	wire _dataUnits_30_io_validOut;
	wire [255:0] _dataUnits_29_io_taskOut;
	wire _dataUnits_29_io_validOut;
	wire [255:0] _dataUnits_28_io_taskOut;
	wire _dataUnits_28_io_validOut;
	wire [255:0] _dataUnits_27_io_taskOut;
	wire _dataUnits_27_io_validOut;
	wire [255:0] _dataUnits_26_io_taskOut;
	wire _dataUnits_26_io_validOut;
	wire [255:0] _dataUnits_25_io_taskOut;
	wire _dataUnits_25_io_validOut;
	wire [255:0] _dataUnits_24_io_taskOut;
	wire _dataUnits_24_io_validOut;
	wire [255:0] _dataUnits_23_io_taskOut;
	wire _dataUnits_23_io_validOut;
	wire [255:0] _dataUnits_22_io_taskOut;
	wire _dataUnits_22_io_validOut;
	wire [255:0] _dataUnits_21_io_taskOut;
	wire _dataUnits_21_io_validOut;
	wire [255:0] _dataUnits_20_io_taskOut;
	wire _dataUnits_20_io_validOut;
	wire [255:0] _dataUnits_19_io_taskOut;
	wire _dataUnits_19_io_validOut;
	wire [255:0] _dataUnits_18_io_taskOut;
	wire _dataUnits_18_io_validOut;
	wire [255:0] _dataUnits_17_io_taskOut;
	wire _dataUnits_17_io_validOut;
	wire [255:0] _dataUnits_16_io_taskOut;
	wire _dataUnits_16_io_validOut;
	wire [255:0] _dataUnits_15_io_taskOut;
	wire _dataUnits_15_io_validOut;
	wire [255:0] _dataUnits_14_io_taskOut;
	wire _dataUnits_14_io_validOut;
	wire [255:0] _dataUnits_13_io_taskOut;
	wire _dataUnits_13_io_validOut;
	wire [255:0] _dataUnits_12_io_taskOut;
	wire _dataUnits_12_io_validOut;
	wire [255:0] _dataUnits_11_io_taskOut;
	wire _dataUnits_11_io_validOut;
	wire [255:0] _dataUnits_10_io_taskOut;
	wire _dataUnits_10_io_validOut;
	wire [255:0] _dataUnits_9_io_taskOut;
	wire _dataUnits_9_io_validOut;
	wire [255:0] _dataUnits_8_io_taskOut;
	wire _dataUnits_8_io_validOut;
	wire [255:0] _dataUnits_7_io_taskOut;
	wire _dataUnits_7_io_validOut;
	wire [255:0] _dataUnits_6_io_taskOut;
	wire _dataUnits_6_io_validOut;
	wire [255:0] _dataUnits_5_io_taskOut;
	wire _dataUnits_5_io_validOut;
	wire [255:0] _dataUnits_4_io_taskOut;
	wire _dataUnits_4_io_validOut;
	wire [255:0] _dataUnits_3_io_taskOut;
	wire _dataUnits_3_io_validOut;
	wire [255:0] _dataUnits_2_io_taskOut;
	wire _dataUnits_2_io_validOut;
	wire [255:0] _dataUnits_1_io_taskOut;
	wire _dataUnits_1_io_validOut;
	wire [255:0] _dataUnits_0_io_taskOut;
	wire _dataUnits_0_io_validOut;
	SchedulerNetworkDataUnit dataUnits_0(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_64_io_taskOut),
		.io_taskOut(_dataUnits_0_io_taskOut),
		.io_validIn(_dataUnits_64_io_validOut),
		.io_validOut(_dataUnits_0_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_0_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_0_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_0_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_0_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_0_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_0_data_qOutTask_bits),
		.io_occupied(io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerNetworkDataUnit dataUnits_1(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_0_io_taskOut),
		.io_taskOut(_dataUnits_1_io_taskOut),
		.io_validIn(_dataUnits_0_io_validOut),
		.io_validOut(_dataUnits_1_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_1_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_1_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_1_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_1_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_1_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_1_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_2(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_1_io_taskOut),
		.io_taskOut(_dataUnits_2_io_taskOut),
		.io_validIn(_dataUnits_1_io_validOut),
		.io_validOut(_dataUnits_2_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_2_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_2_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_2_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_2_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_2_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_2_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_3(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_2_io_taskOut),
		.io_taskOut(_dataUnits_3_io_taskOut),
		.io_validIn(_dataUnits_2_io_validOut),
		.io_validOut(_dataUnits_3_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_3_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_3_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_3_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_3_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_3_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_3_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_4(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_3_io_taskOut),
		.io_taskOut(_dataUnits_4_io_taskOut),
		.io_validIn(_dataUnits_3_io_validOut),
		.io_validOut(_dataUnits_4_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_4_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_4_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_4_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_4_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_4_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_4_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_5(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_4_io_taskOut),
		.io_taskOut(_dataUnits_5_io_taskOut),
		.io_validIn(_dataUnits_4_io_validOut),
		.io_validOut(_dataUnits_5_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_5_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_5_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_5_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_5_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_5_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_5_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_6(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_5_io_taskOut),
		.io_taskOut(_dataUnits_6_io_taskOut),
		.io_validIn(_dataUnits_5_io_validOut),
		.io_validOut(_dataUnits_6_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_6_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_6_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_6_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_6_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_6_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_6_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_7(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_6_io_taskOut),
		.io_taskOut(_dataUnits_7_io_taskOut),
		.io_validIn(_dataUnits_6_io_validOut),
		.io_validOut(_dataUnits_7_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_7_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_7_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_7_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_7_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_7_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_7_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_8(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_7_io_taskOut),
		.io_taskOut(_dataUnits_8_io_taskOut),
		.io_validIn(_dataUnits_7_io_validOut),
		.io_validOut(_dataUnits_8_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_8_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_8_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_8_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_8_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_8_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_8_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_9(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_8_io_taskOut),
		.io_taskOut(_dataUnits_9_io_taskOut),
		.io_validIn(_dataUnits_8_io_validOut),
		.io_validOut(_dataUnits_9_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_9_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_9_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_9_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_9_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_9_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_9_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_10(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_9_io_taskOut),
		.io_taskOut(_dataUnits_10_io_taskOut),
		.io_validIn(_dataUnits_9_io_validOut),
		.io_validOut(_dataUnits_10_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_10_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_10_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_10_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_10_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_10_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_10_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_11(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_10_io_taskOut),
		.io_taskOut(_dataUnits_11_io_taskOut),
		.io_validIn(_dataUnits_10_io_validOut),
		.io_validOut(_dataUnits_11_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_11_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_11_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_11_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_11_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_11_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_11_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_12(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_11_io_taskOut),
		.io_taskOut(_dataUnits_12_io_taskOut),
		.io_validIn(_dataUnits_11_io_validOut),
		.io_validOut(_dataUnits_12_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_12_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_12_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_12_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_12_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_12_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_12_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_13(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_12_io_taskOut),
		.io_taskOut(_dataUnits_13_io_taskOut),
		.io_validIn(_dataUnits_12_io_validOut),
		.io_validOut(_dataUnits_13_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_13_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_13_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_13_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_13_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_13_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_13_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_14(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_13_io_taskOut),
		.io_taskOut(_dataUnits_14_io_taskOut),
		.io_validIn(_dataUnits_13_io_validOut),
		.io_validOut(_dataUnits_14_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_14_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_14_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_14_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_14_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_14_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_14_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_15(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_14_io_taskOut),
		.io_taskOut(_dataUnits_15_io_taskOut),
		.io_validIn(_dataUnits_14_io_validOut),
		.io_validOut(_dataUnits_15_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_15_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_15_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_15_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_15_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_15_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_15_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_16(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_15_io_taskOut),
		.io_taskOut(_dataUnits_16_io_taskOut),
		.io_validIn(_dataUnits_15_io_validOut),
		.io_validOut(_dataUnits_16_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_16_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_16_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_16_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_16_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_16_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_16_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_17(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_16_io_taskOut),
		.io_taskOut(_dataUnits_17_io_taskOut),
		.io_validIn(_dataUnits_16_io_validOut),
		.io_validOut(_dataUnits_17_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_17_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_17_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_17_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_17_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_17_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_17_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_18(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_17_io_taskOut),
		.io_taskOut(_dataUnits_18_io_taskOut),
		.io_validIn(_dataUnits_17_io_validOut),
		.io_validOut(_dataUnits_18_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_18_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_18_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_18_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_18_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_18_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_18_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_19(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_18_io_taskOut),
		.io_taskOut(_dataUnits_19_io_taskOut),
		.io_validIn(_dataUnits_18_io_validOut),
		.io_validOut(_dataUnits_19_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_19_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_19_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_19_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_19_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_19_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_19_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_20(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_19_io_taskOut),
		.io_taskOut(_dataUnits_20_io_taskOut),
		.io_validIn(_dataUnits_19_io_validOut),
		.io_validOut(_dataUnits_20_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_20_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_20_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_20_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_20_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_20_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_20_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_21(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_20_io_taskOut),
		.io_taskOut(_dataUnits_21_io_taskOut),
		.io_validIn(_dataUnits_20_io_validOut),
		.io_validOut(_dataUnits_21_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_21_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_21_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_21_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_21_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_21_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_21_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_22(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_21_io_taskOut),
		.io_taskOut(_dataUnits_22_io_taskOut),
		.io_validIn(_dataUnits_21_io_validOut),
		.io_validOut(_dataUnits_22_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_22_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_22_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_22_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_22_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_22_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_22_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_23(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_22_io_taskOut),
		.io_taskOut(_dataUnits_23_io_taskOut),
		.io_validIn(_dataUnits_22_io_validOut),
		.io_validOut(_dataUnits_23_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_23_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_23_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_23_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_23_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_23_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_23_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_24(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_23_io_taskOut),
		.io_taskOut(_dataUnits_24_io_taskOut),
		.io_validIn(_dataUnits_23_io_validOut),
		.io_validOut(_dataUnits_24_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_24_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_24_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_24_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_24_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_24_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_24_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_25(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_24_io_taskOut),
		.io_taskOut(_dataUnits_25_io_taskOut),
		.io_validIn(_dataUnits_24_io_validOut),
		.io_validOut(_dataUnits_25_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_25_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_25_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_25_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_25_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_25_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_25_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_26(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_25_io_taskOut),
		.io_taskOut(_dataUnits_26_io_taskOut),
		.io_validIn(_dataUnits_25_io_validOut),
		.io_validOut(_dataUnits_26_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_26_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_26_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_26_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_26_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_26_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_26_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_27(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_26_io_taskOut),
		.io_taskOut(_dataUnits_27_io_taskOut),
		.io_validIn(_dataUnits_26_io_validOut),
		.io_validOut(_dataUnits_27_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_27_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_27_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_27_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_27_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_27_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_27_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_28(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_27_io_taskOut),
		.io_taskOut(_dataUnits_28_io_taskOut),
		.io_validIn(_dataUnits_27_io_validOut),
		.io_validOut(_dataUnits_28_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_28_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_28_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_28_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_28_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_28_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_28_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_29(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_28_io_taskOut),
		.io_taskOut(_dataUnits_29_io_taskOut),
		.io_validIn(_dataUnits_28_io_validOut),
		.io_validOut(_dataUnits_29_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_29_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_29_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_29_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_29_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_29_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_29_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_30(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_29_io_taskOut),
		.io_taskOut(_dataUnits_30_io_taskOut),
		.io_validIn(_dataUnits_29_io_validOut),
		.io_validOut(_dataUnits_30_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_30_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_30_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_30_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_30_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_30_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_30_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_31(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_30_io_taskOut),
		.io_taskOut(_dataUnits_31_io_taskOut),
		.io_validIn(_dataUnits_30_io_validOut),
		.io_validOut(_dataUnits_31_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_31_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_31_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_31_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_31_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_31_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_31_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_32(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_31_io_taskOut),
		.io_taskOut(_dataUnits_32_io_taskOut),
		.io_validIn(_dataUnits_31_io_validOut),
		.io_validOut(_dataUnits_32_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_32_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_32_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_32_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_32_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_32_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_32_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_33(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_32_io_taskOut),
		.io_taskOut(_dataUnits_33_io_taskOut),
		.io_validIn(_dataUnits_32_io_validOut),
		.io_validOut(_dataUnits_33_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_33_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_33_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_33_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_33_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_33_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_33_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_34(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_33_io_taskOut),
		.io_taskOut(_dataUnits_34_io_taskOut),
		.io_validIn(_dataUnits_33_io_validOut),
		.io_validOut(_dataUnits_34_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_34_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_34_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_34_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_34_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_34_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_34_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_35(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_34_io_taskOut),
		.io_taskOut(_dataUnits_35_io_taskOut),
		.io_validIn(_dataUnits_34_io_validOut),
		.io_validOut(_dataUnits_35_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_35_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_35_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_35_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_35_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_35_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_35_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_36(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_35_io_taskOut),
		.io_taskOut(_dataUnits_36_io_taskOut),
		.io_validIn(_dataUnits_35_io_validOut),
		.io_validOut(_dataUnits_36_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_36_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_36_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_36_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_36_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_36_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_36_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_37(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_36_io_taskOut),
		.io_taskOut(_dataUnits_37_io_taskOut),
		.io_validIn(_dataUnits_36_io_validOut),
		.io_validOut(_dataUnits_37_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_37_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_37_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_37_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_37_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_37_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_37_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_38(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_37_io_taskOut),
		.io_taskOut(_dataUnits_38_io_taskOut),
		.io_validIn(_dataUnits_37_io_validOut),
		.io_validOut(_dataUnits_38_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_38_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_38_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_38_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_38_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_38_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_38_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_39(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_38_io_taskOut),
		.io_taskOut(_dataUnits_39_io_taskOut),
		.io_validIn(_dataUnits_38_io_validOut),
		.io_validOut(_dataUnits_39_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_39_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_39_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_39_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_39_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_39_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_39_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_40(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_39_io_taskOut),
		.io_taskOut(_dataUnits_40_io_taskOut),
		.io_validIn(_dataUnits_39_io_validOut),
		.io_validOut(_dataUnits_40_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_40_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_40_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_40_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_40_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_40_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_40_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_41(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_40_io_taskOut),
		.io_taskOut(_dataUnits_41_io_taskOut),
		.io_validIn(_dataUnits_40_io_validOut),
		.io_validOut(_dataUnits_41_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_41_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_41_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_41_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_41_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_41_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_41_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_42(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_41_io_taskOut),
		.io_taskOut(_dataUnits_42_io_taskOut),
		.io_validIn(_dataUnits_41_io_validOut),
		.io_validOut(_dataUnits_42_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_42_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_42_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_42_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_42_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_42_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_42_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_43(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_42_io_taskOut),
		.io_taskOut(_dataUnits_43_io_taskOut),
		.io_validIn(_dataUnits_42_io_validOut),
		.io_validOut(_dataUnits_43_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_43_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_43_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_43_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_43_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_43_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_43_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_44(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_43_io_taskOut),
		.io_taskOut(_dataUnits_44_io_taskOut),
		.io_validIn(_dataUnits_43_io_validOut),
		.io_validOut(_dataUnits_44_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_44_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_44_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_44_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_44_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_44_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_44_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_45(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_44_io_taskOut),
		.io_taskOut(_dataUnits_45_io_taskOut),
		.io_validIn(_dataUnits_44_io_validOut),
		.io_validOut(_dataUnits_45_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_45_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_45_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_45_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_45_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_45_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_45_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_46(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_45_io_taskOut),
		.io_taskOut(_dataUnits_46_io_taskOut),
		.io_validIn(_dataUnits_45_io_validOut),
		.io_validOut(_dataUnits_46_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_46_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_46_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_46_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_46_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_46_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_46_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_47(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_46_io_taskOut),
		.io_taskOut(_dataUnits_47_io_taskOut),
		.io_validIn(_dataUnits_46_io_validOut),
		.io_validOut(_dataUnits_47_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_47_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_47_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_47_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_47_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_47_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_47_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_48(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_47_io_taskOut),
		.io_taskOut(_dataUnits_48_io_taskOut),
		.io_validIn(_dataUnits_47_io_validOut),
		.io_validOut(_dataUnits_48_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_48_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_48_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_48_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_48_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_48_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_48_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_49(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_48_io_taskOut),
		.io_taskOut(_dataUnits_49_io_taskOut),
		.io_validIn(_dataUnits_48_io_validOut),
		.io_validOut(_dataUnits_49_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_49_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_49_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_49_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_49_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_49_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_49_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_50(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_49_io_taskOut),
		.io_taskOut(_dataUnits_50_io_taskOut),
		.io_validIn(_dataUnits_49_io_validOut),
		.io_validOut(_dataUnits_50_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_50_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_50_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_50_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_50_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_50_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_50_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_51(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_50_io_taskOut),
		.io_taskOut(_dataUnits_51_io_taskOut),
		.io_validIn(_dataUnits_50_io_validOut),
		.io_validOut(_dataUnits_51_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_51_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_51_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_51_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_51_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_51_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_51_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_52(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_51_io_taskOut),
		.io_taskOut(_dataUnits_52_io_taskOut),
		.io_validIn(_dataUnits_51_io_validOut),
		.io_validOut(_dataUnits_52_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_52_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_52_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_52_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_52_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_52_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_52_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_53(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_52_io_taskOut),
		.io_taskOut(_dataUnits_53_io_taskOut),
		.io_validIn(_dataUnits_52_io_validOut),
		.io_validOut(_dataUnits_53_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_53_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_53_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_53_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_53_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_53_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_53_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_54(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_53_io_taskOut),
		.io_taskOut(_dataUnits_54_io_taskOut),
		.io_validIn(_dataUnits_53_io_validOut),
		.io_validOut(_dataUnits_54_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_54_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_54_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_54_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_54_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_54_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_54_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_55(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_54_io_taskOut),
		.io_taskOut(_dataUnits_55_io_taskOut),
		.io_validIn(_dataUnits_54_io_validOut),
		.io_validOut(_dataUnits_55_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_55_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_55_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_55_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_55_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_55_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_55_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_56(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_55_io_taskOut),
		.io_taskOut(_dataUnits_56_io_taskOut),
		.io_validIn(_dataUnits_55_io_validOut),
		.io_validOut(_dataUnits_56_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_56_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_56_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_56_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_56_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_56_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_56_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_57(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_56_io_taskOut),
		.io_taskOut(_dataUnits_57_io_taskOut),
		.io_validIn(_dataUnits_56_io_validOut),
		.io_validOut(_dataUnits_57_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_57_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_57_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_57_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_57_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_57_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_57_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_58(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_57_io_taskOut),
		.io_taskOut(_dataUnits_58_io_taskOut),
		.io_validIn(_dataUnits_57_io_validOut),
		.io_validOut(_dataUnits_58_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_58_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_58_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_58_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_58_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_58_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_58_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_59(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_58_io_taskOut),
		.io_taskOut(_dataUnits_59_io_taskOut),
		.io_validIn(_dataUnits_58_io_validOut),
		.io_validOut(_dataUnits_59_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_59_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_59_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_59_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_59_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_59_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_59_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_60(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_59_io_taskOut),
		.io_taskOut(_dataUnits_60_io_taskOut),
		.io_validIn(_dataUnits_59_io_validOut),
		.io_validOut(_dataUnits_60_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_60_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_60_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_60_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_60_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_60_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_60_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_61(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_60_io_taskOut),
		.io_taskOut(_dataUnits_61_io_taskOut),
		.io_validIn(_dataUnits_60_io_validOut),
		.io_validOut(_dataUnits_61_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_61_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_61_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_61_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_61_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_61_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_61_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_62(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_61_io_taskOut),
		.io_taskOut(_dataUnits_62_io_taskOut),
		.io_validIn(_dataUnits_61_io_validOut),
		.io_validOut(_dataUnits_62_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_62_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_62_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_62_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_62_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_62_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_62_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_63(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_62_io_taskOut),
		.io_taskOut(_dataUnits_63_io_taskOut),
		.io_validIn(_dataUnits_62_io_validOut),
		.io_validOut(_dataUnits_63_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_63_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_63_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_63_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_63_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_63_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_63_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit dataUnits_64(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_63_io_taskOut),
		.io_taskOut(_dataUnits_64_io_taskOut),
		.io_validIn(_dataUnits_63_io_validOut),
		.io_validOut(_dataUnits_64_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_64_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_64_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_64_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_64_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_64_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_64_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkControlUnit ctrlunits_0(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_1_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_0_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_0_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_0_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_1(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_2_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_1_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_1_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_1_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_1_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_1_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_2(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_3_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_2_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_2_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_2_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_2_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_2_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_3(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_4_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_3_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_3_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_3_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_3_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_3_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_4(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_5_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_4_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_4_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_4_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_4_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_4_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_5(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_6_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_5_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_5_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_5_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_5_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_5_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_6(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_7_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_6_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_6_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_6_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_6_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_6_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_7(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_8_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_7_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_7_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_7_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_7_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_7_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_8(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_9_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_8_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_8_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_8_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_8_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_8_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_9(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_10_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_9_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_9_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_9_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_9_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_9_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_10(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_11_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_10_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_10_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_10_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_10_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_10_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_11(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_12_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_11_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_11_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_11_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_11_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_11_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_12(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_13_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_12_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_12_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_12_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_12_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_12_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_13(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_14_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_13_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_13_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_13_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_13_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_13_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_14(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_15_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_14_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_14_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_14_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_14_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_14_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_15(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_16_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_15_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_15_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_15_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_15_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_15_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_16(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_17_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_16_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_16_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_16_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_16_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_16_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_17(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_18_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_17_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_17_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_17_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_17_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_18(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_19_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_18_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_18_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_18_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_18_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_19(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_20_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_19_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_19_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_19_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_19_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_20(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_21_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_20_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_20_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_20_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_20_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_21(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_22_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_21_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_21_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_21_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_21_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_22(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_23_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_22_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_22_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_22_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_22_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_23(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_24_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_23_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_23_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_23_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_23_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_24(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_25_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_24_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_24_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_24_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_24_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_25(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_26_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_25_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_25_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_25_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_25_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_26(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_27_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_26_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_26_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_26_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_26_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_27(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_28_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_27_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_27_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_27_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_27_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_28(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_29_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_28_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_28_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_28_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_28_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_29(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_30_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_29_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_29_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_29_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_29_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_30(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_31_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_30_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_30_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_30_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_30_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_31(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_32_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_31_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_31_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_31_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_31_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_32(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_33_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_32_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_32_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_32_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_32_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_33(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_34_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_33_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_33_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_33_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_33_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_33_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_34(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_35_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_34_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_34_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_34_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_34_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_34_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_35(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_36_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_35_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_35_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_35_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_35_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_35_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_36(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_37_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_36_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_36_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_36_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_36_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_36_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_37(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_38_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_37_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_37_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_37_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_37_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_37_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_38(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_39_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_38_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_38_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_38_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_38_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_38_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_39(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_40_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_39_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_39_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_39_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_39_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_39_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_40(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_41_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_40_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_40_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_40_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_40_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_40_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_41(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_42_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_41_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_41_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_41_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_41_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_41_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_42(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_43_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_42_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_42_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_42_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_42_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_42_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_43(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_44_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_43_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_43_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_43_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_43_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_43_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_44(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_45_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_44_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_44_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_44_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_44_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_44_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_45(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_46_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_45_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_45_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_45_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_45_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_45_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_46(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_47_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_46_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_46_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_46_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_46_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_46_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_47(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_48_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_47_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_47_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_47_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_47_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_47_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_48(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_49_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_48_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_48_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_48_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_48_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_48_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_49(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_50_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_49_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_49_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_49_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_49_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_49_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_50(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_51_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_50_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_50_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_50_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_50_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_50_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_51(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_52_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_51_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_51_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_51_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_51_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_51_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_52(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_53_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_52_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_52_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_52_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_52_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_52_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_53(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_54_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_53_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_53_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_53_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_53_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_53_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_54(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_55_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_54_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_54_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_54_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_54_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_54_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_55(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_56_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_55_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_55_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_55_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_55_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_55_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_56(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_57_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_56_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_56_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_56_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_56_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_56_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_57(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_58_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_57_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_57_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_57_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_57_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_57_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_58(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_59_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_58_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_58_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_58_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_58_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_58_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_59(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_60_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_59_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_59_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_59_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_59_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_59_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_60(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_61_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_60_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_60_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_60_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_60_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_60_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_61(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_62_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_61_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_61_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_61_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_61_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_61_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_62(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_63_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_62_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_62_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_62_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_62_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_62_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_63(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_64_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_63_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_63_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_63_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_63_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_63_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_64(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_0_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_64_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_64_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_64_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_64_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_64_ctrl_stealReq_ready)
	);
endmodule
module SchedulerClient (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_ctrl_stealReq_valid,
	io_connNetwork_ctrl_stealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_connQ_currLength,
	io_connQ_push_ready,
	io_connQ_push_valid,
	io_connQ_push_bits,
	io_connQ_pop_ready,
	io_connQ_pop_valid,
	io_connQ_pop_bits
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_ctrl_stealReq_valid;
	input io_connNetwork_ctrl_stealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [255:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [255:0] io_connNetwork_data_qOutTask_bits;
	input [7:0] io_connQ_currLength;
	input io_connQ_push_ready;
	output wire io_connQ_push_valid;
	output wire [255:0] io_connQ_push_bits;
	output wire io_connQ_pop_ready;
	input io_connQ_pop_valid;
	input [255:0] io_connQ_pop_bits;
	reg [2:0] stateReg;
	reg [255:0] stolenTaskReg;
	reg [255:0] giveTaskReg;
	reg [1:0] taskRequestCount;
	reg [31:0] tasksGivenAwayCount;
	reg [31:0] requestKilledCount;
	reg [31:0] requestFullCount;
	wire _GEN = stateReg == 3'h0;
	wire _GEN_0 = stateReg == 3'h1;
	wire _GEN_1 = io_connNetwork_ctrl_stealReq_ready & (taskRequestCount == 2'h1);
	wire _GEN_2 = io_connNetwork_ctrl_stealReq_ready & (taskRequestCount == 2'h2);
	wire _GEN_3 = _GEN_2 | (|io_connQ_currLength[7:2]);
	wire _GEN_4 = _GEN_1 | _GEN_3;
	wire _GEN_5 = stateReg == 3'h2;
	wire _GEN_6 = _GEN | _GEN_0;
	wire _GEN_7 = stateReg == 3'h3;
	wire _GEN_8 = (_GEN | _GEN_0) | _GEN_5;
	wire _GEN_9 = stateReg == 3'h4;
	wire _GEN_10 = stateReg == 3'h5;
	wire _GEN_11 = (_GEN_5 | _GEN_7) | _GEN_9;
	wire _GEN_12 = (_GEN | _GEN_0) | _GEN_11;
	wire _GEN_13 = stateReg == 3'h6;
	wire _GEN_14 = ((_GEN_5 | _GEN_7) | _GEN_9) | _GEN_10;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 3'h0;
			stolenTaskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			giveTaskReg <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			taskRequestCount <= 2'h1;
			tasksGivenAwayCount <= 32'h00000000;
			requestKilledCount <= 32'h00000041;
			requestFullCount <= 32'h00000041;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_15;
			reg _GEN_16;
			reg _GEN_17;
			reg _GEN_18;
			reg _GEN_19;
			reg [31:0] _GEN_20;
			reg _GEN_21;
			reg _GEN_22;
			reg _GEN_23;
			reg [1:0] _GEN_24;
			reg [23:0] _GEN_25;
			reg [15:0] _GEN_26;
			reg [255:0] _GEN_27;
			_GEN_16 = io_connQ_currLength > 8'h59;
			_GEN_20 = (_GEN_11 | ~(_GEN_10 & io_connNetwork_data_qOutTask_ready) ? tasksGivenAwayCount : tasksGivenAwayCount + 32'h00000001);
			_GEN_27 = {_GEN_20, _GEN_20, _GEN_20, tasksGivenAwayCount, tasksGivenAwayCount, tasksGivenAwayCount, (_GEN_4 | ~(|tasksGivenAwayCount) ? tasksGivenAwayCount : tasksGivenAwayCount - 32'h00000001), tasksGivenAwayCount};
			_GEN_15 = io_connQ_currLength < 8'h04;
			_GEN_17 = requestKilledCount == 32'h00000000;
			_GEN_18 = io_connQ_currLength > 8'h58;
			_GEN_19 = io_connQ_currLength == 8'h00;
			_GEN_21 = _GEN_16 | (io_connNetwork_ctrl_serveStealReq_ready & |io_connQ_currLength[7:2]);
			_GEN_22 = _GEN_15 & io_connNetwork_ctrl_serveStealReq_ready;
			_GEN_23 = _GEN_22 | _GEN_15;
			_GEN_24 = ((_GEN_14 | ~_GEN_13) | _GEN_21 ? taskRequestCount : (_GEN_22 ? 2'h2 : (_GEN_15 ? 2'h1 : taskRequestCount)));
			_GEN_25 = {stateReg, (_GEN_21 ? 3'h4 : (_GEN_23 ? 3'h1 : 3'h6)), (io_connNetwork_data_qOutTask_ready ? 3'h0 : 3'h5), (io_connQ_pop_valid ? 3'h5 : (_GEN_19 ? 3'h1 : 3'h4)), (io_connQ_push_ready ? 3'h0 : (_GEN_18 ? 3'h5 : 3'h3)), (io_connNetwork_data_availableTask_valid ? 3'h3 : (|io_connQ_currLength[7:2] ? 3'h0 : (_GEN_17 ? 3'h1 : 3'h2))), (_GEN_1 ? 3'h2 : (_GEN_2 ? 3'h1 : (|io_connQ_currLength[7:2] ? 3'h6 : (|tasksGivenAwayCount | (requestFullCount == 32'h00000000) ? 3'h2 : 3'h1)))), (_GEN_15 ? 3'h1 : (_GEN_16 ? 3'h4 : (io_connQ_currLength > 8'h04 ? 3'h6 : 3'h0)))};
			stateReg <= _GEN_25[stateReg * 3+:3];
			if (_GEN_6 | ~(_GEN_5 & io_connNetwork_data_availableTask_valid))
				;
			else
				stolenTaskReg <= io_connNetwork_data_availableTask_bits;
			if (~_GEN_8) begin
				if (_GEN_7) begin
					if (io_connQ_push_ready | ~_GEN_18)
						;
					else
						giveTaskReg <= stolenTaskReg;
				end
				else if (_GEN_9 & io_connQ_pop_valid)
					giveTaskReg <= io_connQ_pop_bits;
			end
			_GEN_26 = {_GEN_24, _GEN_24, taskRequestCount, taskRequestCount, taskRequestCount, taskRequestCount, (_GEN_1 | ~_GEN_2 ? taskRequestCount : 2'h1), taskRequestCount};
			taskRequestCount <= _GEN_26[stateReg * 2+:2];
			tasksGivenAwayCount <= _GEN_27[stateReg * 32+:32];
			if (_GEN) begin
				if (_GEN_15)
					requestFullCount <= 32'h00000041;
			end
			else if (_GEN_0) begin
				if (_GEN_1 | ~(_GEN_3 | ~(|tasksGivenAwayCount)))
					requestKilledCount <= 32'h00000041;
				if (io_connNetwork_ctrl_serveStealReq_ready)
					requestFullCount <= requestFullCount - 32'h00000001;
				else
					requestFullCount <= 32'h00000041;
			end
			else begin
				if (_GEN_5) begin
					if (io_connNetwork_ctrl_serveStealReq_ready)
						requestKilledCount <= 32'h00000041;
					else
						requestKilledCount <= requestKilledCount - 32'h00000001;
				end
				if ((_GEN_5 ? (io_connNetwork_data_availableTask_valid | (|io_connQ_currLength[7:2])) | ~_GEN_17 : _GEN_7 | (_GEN_9 ? io_connQ_pop_valid | ~_GEN_19 : ((_GEN_10 | ~_GEN_13) | _GEN_21) | ~_GEN_23)))
					;
				else
					requestFullCount <= 32'h00000041;
			end
		end
	assign io_connNetwork_ctrl_serveStealReq_valid = ~_GEN & (_GEN_0 ? ~_GEN_4 & |tasksGivenAwayCount : ~_GEN_14 & _GEN_13);
	assign io_connNetwork_ctrl_stealReq_valid = ~_GEN & _GEN_0;
	assign io_connNetwork_data_availableTask_ready = ~_GEN_6 & _GEN_5;
	assign io_connNetwork_data_qOutTask_valid = ~_GEN_12 & _GEN_10;
	assign io_connNetwork_data_qOutTask_bits = (_GEN_12 | ~_GEN_10 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : giveTaskReg);
	assign io_connQ_push_valid = ~_GEN_8 & _GEN_7;
	assign io_connQ_push_bits = (_GEN_8 | ~_GEN_7 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : stolenTaskReg);
	assign io_connQ_pop_ready = ~(((_GEN | _GEN_0) | _GEN_5) | _GEN_7) & _GEN_9;
endmodule
module hw_deque (
	clock,
	reset,
	io_connVec_0_push_ready,
	io_connVec_0_push_valid,
	io_connVec_0_push_bits,
	io_connVec_0_pop_ready,
	io_connVec_0_pop_valid,
	io_connVec_1_currLength,
	io_connVec_1_push_ready,
	io_connVec_1_push_valid,
	io_connVec_1_push_bits,
	io_connVec_1_pop_ready,
	io_connVec_1_pop_valid,
	io_connVec_1_pop_bits
);
	input clock;
	input reset;
	output wire io_connVec_0_push_ready;
	input io_connVec_0_push_valid;
	input [255:0] io_connVec_0_push_bits;
	input io_connVec_0_pop_ready;
	output wire io_connVec_0_pop_valid;
	output wire [8:0] io_connVec_1_currLength;
	output wire io_connVec_1_push_ready;
	input io_connVec_1_push_valid;
	input [255:0] io_connVec_1_push_bits;
	input io_connVec_1_pop_ready;
	output wire io_connVec_1_pop_valid;
	output wire [255:0] io_connVec_1_pop_bits;
	wire [255:0] _bramMem_b_dout;
	reg [8:0] sideReg_0;
	reg [8:0] sideReg_1;
	reg readLatency_0;
	reg readLatency_1;
	reg writeLatency_0;
	reg writeLatency_1;
	reg [2:0] stateRegs_0;
	reg [2:0] stateRegs_1;
	wire _GEN = stateRegs_0 == 3'h0;
	wire _GEN_0 = stateRegs_1 == 3'h0;
	wire _GEN_1 = stateRegs_0 == 3'h1;
	wire _GEN_2 = stateRegs_0 == 3'h2;
	wire _GEN_3 = sideReg_0 == 9'h081;
	wire _GEN_4 = stateRegs_0 == 3'h4;
	wire [8:0] _bramMem_io_a_addr_T_2 = sideReg_0 + 9'h001;
	wire _GEN_5 = (_GEN | _GEN_1) | _GEN_2;
	wire _GEN_6 = stateRegs_0 == 3'h3;
	wire _GEN_7 = stateRegs_1 == 3'h1;
	wire _GEN_8 = stateRegs_1 == 3'h2;
	wire _GEN_9 = sideReg_1 == 9'h000;
	wire _GEN_10 = stateRegs_1 == 3'h4;
	wire [8:0] _bramMem_io_b_addr_T_6 = sideReg_1 - 9'h001;
	wire _GEN_11 = (_GEN_0 | _GEN_7) | _GEN_8;
	wire _GEN_12 = stateRegs_1 == 3'h3;
	wire [8:0] currLen = (sideReg_0 > sideReg_1 ? ((sideReg_1 + 9'h082) - sideReg_0) - 9'h001 : (sideReg_1 - sideReg_0) - 9'h001);
	always @(posedge clock)
		if (reset) begin
			sideReg_0 <= 9'h000;
			sideReg_1 <= 9'h001;
			readLatency_0 <= 1'h0;
			readLatency_1 <= 1'h0;
			writeLatency_0 <= 1'h0;
			writeLatency_1 <= 1'h0;
			stateRegs_0 <= 3'h0;
			stateRegs_1 <= 3'h0;
		end
		else begin : sv2v_autoblock_1
			reg [23:0] _GEN_13;
			reg [23:0] _GEN_14;
			_GEN_13 = {stateRegs_0, stateRegs_0, stateRegs_0, 6'h00, (readLatency_0 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_0, 1'h1, ((io_connVec_0_pop_ready & |currLen[8:1]) | ((io_connVec_0_pop_ready & _GEN_0) & |currLen) ? 3'h2 : {2'h0, io_connVec_0_push_valid & (currLen < 9'h082)})};
			_GEN_14 = {stateRegs_1, stateRegs_1, stateRegs_1, 6'h00, (readLatency_1 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_1, 1'h1, (io_connVec_1_push_valid & (currLen < 9'h081) ? 3'h1 : {1'h0, (io_connVec_1_pop_ready & |currLen[8:1]) | (((io_connVec_1_pop_ready & ~io_connVec_0_pop_ready) & |currLen) & (stateRegs_0 != 3'h4)), 1'h0})};
			if (~_GEN_5) begin
				if (_GEN_4) begin
					if (_GEN_3)
						sideReg_0 <= 9'h000;
					else
						sideReg_0 <= _bramMem_io_a_addr_T_2;
				end
				else if (_GEN_6) begin
					if (sideReg_0 == 9'h000)
						sideReg_0 <= 9'h081;
					else
						sideReg_0 <= sideReg_0 - 9'h001;
				end
			end
			if (~_GEN_11) begin
				if (_GEN_10) begin
					if (_GEN_9)
						sideReg_1 <= 9'h081;
					else
						sideReg_1 <= _bramMem_io_b_addr_T_6;
				end
				else if (_GEN_12) begin
					if (sideReg_1 == 9'h081)
						sideReg_1 <= 9'h000;
					else
						sideReg_1 <= sideReg_1 + 9'h001;
				end
			end
			readLatency_0 <= (((_GEN | _GEN_1) | ~_GEN_2) | (readLatency_0 - 1'h1)) & readLatency_0;
			readLatency_1 <= (((_GEN_0 | _GEN_7) | ~_GEN_8) | (readLatency_1 - 1'h1)) & readLatency_1;
			writeLatency_0 <= ((_GEN | ~_GEN_1) | (writeLatency_0 - 1'h1)) & writeLatency_0;
			writeLatency_1 <= ((_GEN_0 | ~_GEN_7) | (writeLatency_1 - 1'h1)) & writeLatency_1;
			stateRegs_0 <= _GEN_13[stateRegs_0 * 3+:3];
			stateRegs_1 <= _GEN_14[stateRegs_1 * 3+:3];
		end
	DualPortBRAM #(
		.ADDR(11),
		.DATA(256)
	) bramMem(
		.clk(clock),
		.rst(reset),
		.a_addr((_GEN ? 11'h7ff : (_GEN_1 ? {2'h0, sideReg_0} : (_GEN_2 ? (_GEN_3 ? 11'h000 : {2'h0, sideReg_0 + 9'h001}) : (_GEN_4 ? (_GEN_3 ? 11'h000 : {2'h0, _bramMem_io_a_addr_T_2}) : 11'h7ff))))),
		.a_din(io_connVec_0_push_bits),
		.a_wr(~_GEN & _GEN_1),
		.a_dout(),
		.b_addr((_GEN_0 ? 11'h7ff : (_GEN_7 ? {2'h0, sideReg_1} : (_GEN_8 ? (_GEN_9 ? 11'h081 : {2'h0, sideReg_1 - 9'h001}) : (_GEN_10 ? (_GEN_9 ? 11'h081 : {2'h0, _bramMem_io_b_addr_T_6}) : 11'h7ff))))),
		.b_din(io_connVec_1_push_bits),
		.b_wr(~_GEN_0 & _GEN_7),
		.b_dout(_bramMem_b_dout)
	);
	assign io_connVec_0_push_ready = ~(((_GEN | _GEN_1) | _GEN_2) | _GEN_4) & _GEN_6;
	assign io_connVec_0_pop_valid = ~_GEN_5 & _GEN_4;
	assign io_connVec_1_currLength = currLen;
	assign io_connVec_1_push_ready = ~(((_GEN_0 | _GEN_7) | _GEN_8) | _GEN_10) & _GEN_12;
	assign io_connVec_1_pop_valid = ~_GEN_11 & _GEN_10;
	assign io_connVec_1_pop_bits = (_GEN_11 | ~_GEN_10 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : _bramMem_b_dout);
endmodule
module SchedulerLocalNetwork (
	clock,
	reset,
	io_connPE_0_push_ready,
	io_connPE_0_push_valid,
	io_connPE_0_push_bits,
	io_connPE_0_pop_ready,
	io_connPE_0_pop_valid,
	io_connPE_1_push_ready,
	io_connPE_1_push_valid,
	io_connPE_1_push_bits,
	io_connPE_1_pop_ready,
	io_connPE_1_pop_valid,
	io_connPE_2_push_ready,
	io_connPE_2_push_valid,
	io_connPE_2_push_bits,
	io_connPE_2_pop_ready,
	io_connPE_2_pop_valid,
	io_connPE_3_push_ready,
	io_connPE_3_push_valid,
	io_connPE_3_push_bits,
	io_connPE_3_pop_ready,
	io_connPE_3_pop_valid,
	io_connPE_4_push_ready,
	io_connPE_4_push_valid,
	io_connPE_4_push_bits,
	io_connPE_4_pop_ready,
	io_connPE_4_pop_valid,
	io_connPE_5_push_ready,
	io_connPE_5_push_valid,
	io_connPE_5_push_bits,
	io_connPE_5_pop_ready,
	io_connPE_5_pop_valid,
	io_connPE_6_push_ready,
	io_connPE_6_push_valid,
	io_connPE_6_push_bits,
	io_connPE_6_pop_ready,
	io_connPE_6_pop_valid,
	io_connPE_7_push_ready,
	io_connPE_7_push_valid,
	io_connPE_7_push_bits,
	io_connPE_7_pop_ready,
	io_connPE_7_pop_valid,
	io_connPE_8_push_ready,
	io_connPE_8_push_valid,
	io_connPE_8_push_bits,
	io_connPE_8_pop_ready,
	io_connPE_8_pop_valid,
	io_connPE_9_push_ready,
	io_connPE_9_push_valid,
	io_connPE_9_push_bits,
	io_connPE_9_pop_ready,
	io_connPE_9_pop_valid,
	io_connPE_10_push_ready,
	io_connPE_10_push_valid,
	io_connPE_10_push_bits,
	io_connPE_10_pop_ready,
	io_connPE_10_pop_valid,
	io_connPE_11_push_ready,
	io_connPE_11_push_valid,
	io_connPE_11_push_bits,
	io_connPE_11_pop_ready,
	io_connPE_11_pop_valid,
	io_connPE_12_push_ready,
	io_connPE_12_push_valid,
	io_connPE_12_push_bits,
	io_connPE_12_pop_ready,
	io_connPE_12_pop_valid,
	io_connPE_13_push_ready,
	io_connPE_13_push_valid,
	io_connPE_13_push_bits,
	io_connPE_13_pop_ready,
	io_connPE_13_pop_valid,
	io_connPE_14_push_ready,
	io_connPE_14_push_valid,
	io_connPE_14_push_bits,
	io_connPE_14_pop_ready,
	io_connPE_14_pop_valid,
	io_connPE_15_push_ready,
	io_connPE_15_push_valid,
	io_connPE_15_push_bits,
	io_connPE_15_pop_ready,
	io_connPE_15_pop_valid,
	io_connPE_16_push_ready,
	io_connPE_16_push_valid,
	io_connPE_16_push_bits,
	io_connPE_16_pop_ready,
	io_connPE_16_pop_valid,
	io_connPE_17_push_ready,
	io_connPE_17_push_valid,
	io_connPE_17_push_bits,
	io_connPE_17_pop_ready,
	io_connPE_17_pop_valid,
	io_connPE_18_push_ready,
	io_connPE_18_push_valid,
	io_connPE_18_push_bits,
	io_connPE_18_pop_ready,
	io_connPE_18_pop_valid,
	io_connPE_19_push_ready,
	io_connPE_19_push_valid,
	io_connPE_19_push_bits,
	io_connPE_19_pop_ready,
	io_connPE_19_pop_valid,
	io_connPE_20_push_ready,
	io_connPE_20_push_valid,
	io_connPE_20_push_bits,
	io_connPE_20_pop_ready,
	io_connPE_20_pop_valid,
	io_connPE_21_push_ready,
	io_connPE_21_push_valid,
	io_connPE_21_push_bits,
	io_connPE_21_pop_ready,
	io_connPE_21_pop_valid,
	io_connPE_22_push_ready,
	io_connPE_22_push_valid,
	io_connPE_22_push_bits,
	io_connPE_22_pop_ready,
	io_connPE_22_pop_valid,
	io_connPE_23_push_ready,
	io_connPE_23_push_valid,
	io_connPE_23_push_bits,
	io_connPE_23_pop_ready,
	io_connPE_23_pop_valid,
	io_connPE_24_push_ready,
	io_connPE_24_push_valid,
	io_connPE_24_push_bits,
	io_connPE_24_pop_ready,
	io_connPE_24_pop_valid,
	io_connPE_25_push_ready,
	io_connPE_25_push_valid,
	io_connPE_25_push_bits,
	io_connPE_25_pop_ready,
	io_connPE_25_pop_valid,
	io_connPE_26_push_ready,
	io_connPE_26_push_valid,
	io_connPE_26_push_bits,
	io_connPE_26_pop_ready,
	io_connPE_26_pop_valid,
	io_connPE_27_push_ready,
	io_connPE_27_push_valid,
	io_connPE_27_push_bits,
	io_connPE_27_pop_ready,
	io_connPE_27_pop_valid,
	io_connPE_28_push_ready,
	io_connPE_28_push_valid,
	io_connPE_28_push_bits,
	io_connPE_28_pop_ready,
	io_connPE_28_pop_valid,
	io_connPE_29_push_ready,
	io_connPE_29_push_valid,
	io_connPE_29_push_bits,
	io_connPE_29_pop_ready,
	io_connPE_29_pop_valid,
	io_connPE_30_push_ready,
	io_connPE_30_push_valid,
	io_connPE_30_push_bits,
	io_connPE_30_pop_ready,
	io_connPE_30_pop_valid,
	io_connPE_31_push_ready,
	io_connPE_31_push_valid,
	io_connPE_31_push_bits,
	io_connPE_31_pop_ready,
	io_connPE_31_pop_valid,
	io_connPE_32_push_ready,
	io_connPE_32_push_valid,
	io_connPE_32_push_bits,
	io_connPE_32_pop_ready,
	io_connPE_32_pop_valid,
	io_connPE_33_push_ready,
	io_connPE_33_push_valid,
	io_connPE_33_push_bits,
	io_connPE_33_pop_ready,
	io_connPE_33_pop_valid,
	io_connPE_34_push_ready,
	io_connPE_34_push_valid,
	io_connPE_34_push_bits,
	io_connPE_34_pop_ready,
	io_connPE_34_pop_valid,
	io_connPE_35_push_ready,
	io_connPE_35_push_valid,
	io_connPE_35_push_bits,
	io_connPE_35_pop_ready,
	io_connPE_35_pop_valid,
	io_connPE_36_push_ready,
	io_connPE_36_push_valid,
	io_connPE_36_push_bits,
	io_connPE_36_pop_ready,
	io_connPE_36_pop_valid,
	io_connPE_37_push_ready,
	io_connPE_37_push_valid,
	io_connPE_37_push_bits,
	io_connPE_37_pop_ready,
	io_connPE_37_pop_valid,
	io_connPE_38_push_ready,
	io_connPE_38_push_valid,
	io_connPE_38_push_bits,
	io_connPE_38_pop_ready,
	io_connPE_38_pop_valid,
	io_connPE_39_push_ready,
	io_connPE_39_push_valid,
	io_connPE_39_push_bits,
	io_connPE_39_pop_ready,
	io_connPE_39_pop_valid,
	io_connPE_40_push_ready,
	io_connPE_40_push_valid,
	io_connPE_40_push_bits,
	io_connPE_40_pop_ready,
	io_connPE_40_pop_valid,
	io_connPE_41_push_ready,
	io_connPE_41_push_valid,
	io_connPE_41_push_bits,
	io_connPE_41_pop_ready,
	io_connPE_41_pop_valid,
	io_connPE_42_push_ready,
	io_connPE_42_push_valid,
	io_connPE_42_push_bits,
	io_connPE_42_pop_ready,
	io_connPE_42_pop_valid,
	io_connPE_43_push_ready,
	io_connPE_43_push_valid,
	io_connPE_43_push_bits,
	io_connPE_43_pop_ready,
	io_connPE_43_pop_valid,
	io_connPE_44_push_ready,
	io_connPE_44_push_valid,
	io_connPE_44_push_bits,
	io_connPE_44_pop_ready,
	io_connPE_44_pop_valid,
	io_connPE_45_push_ready,
	io_connPE_45_push_valid,
	io_connPE_45_push_bits,
	io_connPE_45_pop_ready,
	io_connPE_45_pop_valid,
	io_connPE_46_push_ready,
	io_connPE_46_push_valid,
	io_connPE_46_push_bits,
	io_connPE_46_pop_ready,
	io_connPE_46_pop_valid,
	io_connPE_47_push_ready,
	io_connPE_47_push_valid,
	io_connPE_47_push_bits,
	io_connPE_47_pop_ready,
	io_connPE_47_pop_valid,
	io_connPE_48_push_ready,
	io_connPE_48_push_valid,
	io_connPE_48_push_bits,
	io_connPE_48_pop_ready,
	io_connPE_48_pop_valid,
	io_connPE_49_push_ready,
	io_connPE_49_push_valid,
	io_connPE_49_push_bits,
	io_connPE_49_pop_ready,
	io_connPE_49_pop_valid,
	io_connPE_50_push_ready,
	io_connPE_50_push_valid,
	io_connPE_50_push_bits,
	io_connPE_50_pop_ready,
	io_connPE_50_pop_valid,
	io_connPE_51_push_ready,
	io_connPE_51_push_valid,
	io_connPE_51_push_bits,
	io_connPE_51_pop_ready,
	io_connPE_51_pop_valid,
	io_connPE_52_push_ready,
	io_connPE_52_push_valid,
	io_connPE_52_push_bits,
	io_connPE_52_pop_ready,
	io_connPE_52_pop_valid,
	io_connPE_53_push_ready,
	io_connPE_53_push_valid,
	io_connPE_53_push_bits,
	io_connPE_53_pop_ready,
	io_connPE_53_pop_valid,
	io_connPE_54_push_ready,
	io_connPE_54_push_valid,
	io_connPE_54_push_bits,
	io_connPE_54_pop_ready,
	io_connPE_54_pop_valid,
	io_connPE_55_push_ready,
	io_connPE_55_push_valid,
	io_connPE_55_push_bits,
	io_connPE_55_pop_ready,
	io_connPE_55_pop_valid,
	io_connPE_56_push_ready,
	io_connPE_56_push_valid,
	io_connPE_56_push_bits,
	io_connPE_56_pop_ready,
	io_connPE_56_pop_valid,
	io_connPE_57_push_ready,
	io_connPE_57_push_valid,
	io_connPE_57_push_bits,
	io_connPE_57_pop_ready,
	io_connPE_57_pop_valid,
	io_connPE_58_push_ready,
	io_connPE_58_push_valid,
	io_connPE_58_push_bits,
	io_connPE_58_pop_ready,
	io_connPE_58_pop_valid,
	io_connPE_59_push_ready,
	io_connPE_59_push_valid,
	io_connPE_59_push_bits,
	io_connPE_59_pop_ready,
	io_connPE_59_pop_valid,
	io_connPE_60_push_ready,
	io_connPE_60_push_valid,
	io_connPE_60_push_bits,
	io_connPE_60_pop_ready,
	io_connPE_60_pop_valid,
	io_connPE_61_push_ready,
	io_connPE_61_push_valid,
	io_connPE_61_push_bits,
	io_connPE_61_pop_ready,
	io_connPE_61_pop_valid,
	io_connPE_62_push_ready,
	io_connPE_62_push_valid,
	io_connPE_62_push_bits,
	io_connPE_62_pop_ready,
	io_connPE_62_pop_valid,
	io_connPE_63_push_ready,
	io_connPE_63_push_valid,
	io_connPE_63_push_bits,
	io_connPE_63_pop_ready,
	io_connPE_63_pop_valid,
	io_connVSS_0_ctrl_serveStealReq_valid,
	io_connVSS_0_ctrl_serveStealReq_ready,
	io_connVSS_0_data_availableTask_ready,
	io_connVSS_0_data_availableTask_valid,
	io_connVSS_0_data_availableTask_bits,
	io_connVSS_0_data_qOutTask_ready,
	io_connVSS_0_data_qOutTask_valid,
	io_connVSS_0_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0
);
	input clock;
	input reset;
	output wire io_connPE_0_push_ready;
	input io_connPE_0_push_valid;
	input [255:0] io_connPE_0_push_bits;
	input io_connPE_0_pop_ready;
	output wire io_connPE_0_pop_valid;
	output wire io_connPE_1_push_ready;
	input io_connPE_1_push_valid;
	input [255:0] io_connPE_1_push_bits;
	input io_connPE_1_pop_ready;
	output wire io_connPE_1_pop_valid;
	output wire io_connPE_2_push_ready;
	input io_connPE_2_push_valid;
	input [255:0] io_connPE_2_push_bits;
	input io_connPE_2_pop_ready;
	output wire io_connPE_2_pop_valid;
	output wire io_connPE_3_push_ready;
	input io_connPE_3_push_valid;
	input [255:0] io_connPE_3_push_bits;
	input io_connPE_3_pop_ready;
	output wire io_connPE_3_pop_valid;
	output wire io_connPE_4_push_ready;
	input io_connPE_4_push_valid;
	input [255:0] io_connPE_4_push_bits;
	input io_connPE_4_pop_ready;
	output wire io_connPE_4_pop_valid;
	output wire io_connPE_5_push_ready;
	input io_connPE_5_push_valid;
	input [255:0] io_connPE_5_push_bits;
	input io_connPE_5_pop_ready;
	output wire io_connPE_5_pop_valid;
	output wire io_connPE_6_push_ready;
	input io_connPE_6_push_valid;
	input [255:0] io_connPE_6_push_bits;
	input io_connPE_6_pop_ready;
	output wire io_connPE_6_pop_valid;
	output wire io_connPE_7_push_ready;
	input io_connPE_7_push_valid;
	input [255:0] io_connPE_7_push_bits;
	input io_connPE_7_pop_ready;
	output wire io_connPE_7_pop_valid;
	output wire io_connPE_8_push_ready;
	input io_connPE_8_push_valid;
	input [255:0] io_connPE_8_push_bits;
	input io_connPE_8_pop_ready;
	output wire io_connPE_8_pop_valid;
	output wire io_connPE_9_push_ready;
	input io_connPE_9_push_valid;
	input [255:0] io_connPE_9_push_bits;
	input io_connPE_9_pop_ready;
	output wire io_connPE_9_pop_valid;
	output wire io_connPE_10_push_ready;
	input io_connPE_10_push_valid;
	input [255:0] io_connPE_10_push_bits;
	input io_connPE_10_pop_ready;
	output wire io_connPE_10_pop_valid;
	output wire io_connPE_11_push_ready;
	input io_connPE_11_push_valid;
	input [255:0] io_connPE_11_push_bits;
	input io_connPE_11_pop_ready;
	output wire io_connPE_11_pop_valid;
	output wire io_connPE_12_push_ready;
	input io_connPE_12_push_valid;
	input [255:0] io_connPE_12_push_bits;
	input io_connPE_12_pop_ready;
	output wire io_connPE_12_pop_valid;
	output wire io_connPE_13_push_ready;
	input io_connPE_13_push_valid;
	input [255:0] io_connPE_13_push_bits;
	input io_connPE_13_pop_ready;
	output wire io_connPE_13_pop_valid;
	output wire io_connPE_14_push_ready;
	input io_connPE_14_push_valid;
	input [255:0] io_connPE_14_push_bits;
	input io_connPE_14_pop_ready;
	output wire io_connPE_14_pop_valid;
	output wire io_connPE_15_push_ready;
	input io_connPE_15_push_valid;
	input [255:0] io_connPE_15_push_bits;
	input io_connPE_15_pop_ready;
	output wire io_connPE_15_pop_valid;
	output wire io_connPE_16_push_ready;
	input io_connPE_16_push_valid;
	input [255:0] io_connPE_16_push_bits;
	input io_connPE_16_pop_ready;
	output wire io_connPE_16_pop_valid;
	output wire io_connPE_17_push_ready;
	input io_connPE_17_push_valid;
	input [255:0] io_connPE_17_push_bits;
	input io_connPE_17_pop_ready;
	output wire io_connPE_17_pop_valid;
	output wire io_connPE_18_push_ready;
	input io_connPE_18_push_valid;
	input [255:0] io_connPE_18_push_bits;
	input io_connPE_18_pop_ready;
	output wire io_connPE_18_pop_valid;
	output wire io_connPE_19_push_ready;
	input io_connPE_19_push_valid;
	input [255:0] io_connPE_19_push_bits;
	input io_connPE_19_pop_ready;
	output wire io_connPE_19_pop_valid;
	output wire io_connPE_20_push_ready;
	input io_connPE_20_push_valid;
	input [255:0] io_connPE_20_push_bits;
	input io_connPE_20_pop_ready;
	output wire io_connPE_20_pop_valid;
	output wire io_connPE_21_push_ready;
	input io_connPE_21_push_valid;
	input [255:0] io_connPE_21_push_bits;
	input io_connPE_21_pop_ready;
	output wire io_connPE_21_pop_valid;
	output wire io_connPE_22_push_ready;
	input io_connPE_22_push_valid;
	input [255:0] io_connPE_22_push_bits;
	input io_connPE_22_pop_ready;
	output wire io_connPE_22_pop_valid;
	output wire io_connPE_23_push_ready;
	input io_connPE_23_push_valid;
	input [255:0] io_connPE_23_push_bits;
	input io_connPE_23_pop_ready;
	output wire io_connPE_23_pop_valid;
	output wire io_connPE_24_push_ready;
	input io_connPE_24_push_valid;
	input [255:0] io_connPE_24_push_bits;
	input io_connPE_24_pop_ready;
	output wire io_connPE_24_pop_valid;
	output wire io_connPE_25_push_ready;
	input io_connPE_25_push_valid;
	input [255:0] io_connPE_25_push_bits;
	input io_connPE_25_pop_ready;
	output wire io_connPE_25_pop_valid;
	output wire io_connPE_26_push_ready;
	input io_connPE_26_push_valid;
	input [255:0] io_connPE_26_push_bits;
	input io_connPE_26_pop_ready;
	output wire io_connPE_26_pop_valid;
	output wire io_connPE_27_push_ready;
	input io_connPE_27_push_valid;
	input [255:0] io_connPE_27_push_bits;
	input io_connPE_27_pop_ready;
	output wire io_connPE_27_pop_valid;
	output wire io_connPE_28_push_ready;
	input io_connPE_28_push_valid;
	input [255:0] io_connPE_28_push_bits;
	input io_connPE_28_pop_ready;
	output wire io_connPE_28_pop_valid;
	output wire io_connPE_29_push_ready;
	input io_connPE_29_push_valid;
	input [255:0] io_connPE_29_push_bits;
	input io_connPE_29_pop_ready;
	output wire io_connPE_29_pop_valid;
	output wire io_connPE_30_push_ready;
	input io_connPE_30_push_valid;
	input [255:0] io_connPE_30_push_bits;
	input io_connPE_30_pop_ready;
	output wire io_connPE_30_pop_valid;
	output wire io_connPE_31_push_ready;
	input io_connPE_31_push_valid;
	input [255:0] io_connPE_31_push_bits;
	input io_connPE_31_pop_ready;
	output wire io_connPE_31_pop_valid;
	output wire io_connPE_32_push_ready;
	input io_connPE_32_push_valid;
	input [255:0] io_connPE_32_push_bits;
	input io_connPE_32_pop_ready;
	output wire io_connPE_32_pop_valid;
	output wire io_connPE_33_push_ready;
	input io_connPE_33_push_valid;
	input [255:0] io_connPE_33_push_bits;
	input io_connPE_33_pop_ready;
	output wire io_connPE_33_pop_valid;
	output wire io_connPE_34_push_ready;
	input io_connPE_34_push_valid;
	input [255:0] io_connPE_34_push_bits;
	input io_connPE_34_pop_ready;
	output wire io_connPE_34_pop_valid;
	output wire io_connPE_35_push_ready;
	input io_connPE_35_push_valid;
	input [255:0] io_connPE_35_push_bits;
	input io_connPE_35_pop_ready;
	output wire io_connPE_35_pop_valid;
	output wire io_connPE_36_push_ready;
	input io_connPE_36_push_valid;
	input [255:0] io_connPE_36_push_bits;
	input io_connPE_36_pop_ready;
	output wire io_connPE_36_pop_valid;
	output wire io_connPE_37_push_ready;
	input io_connPE_37_push_valid;
	input [255:0] io_connPE_37_push_bits;
	input io_connPE_37_pop_ready;
	output wire io_connPE_37_pop_valid;
	output wire io_connPE_38_push_ready;
	input io_connPE_38_push_valid;
	input [255:0] io_connPE_38_push_bits;
	input io_connPE_38_pop_ready;
	output wire io_connPE_38_pop_valid;
	output wire io_connPE_39_push_ready;
	input io_connPE_39_push_valid;
	input [255:0] io_connPE_39_push_bits;
	input io_connPE_39_pop_ready;
	output wire io_connPE_39_pop_valid;
	output wire io_connPE_40_push_ready;
	input io_connPE_40_push_valid;
	input [255:0] io_connPE_40_push_bits;
	input io_connPE_40_pop_ready;
	output wire io_connPE_40_pop_valid;
	output wire io_connPE_41_push_ready;
	input io_connPE_41_push_valid;
	input [255:0] io_connPE_41_push_bits;
	input io_connPE_41_pop_ready;
	output wire io_connPE_41_pop_valid;
	output wire io_connPE_42_push_ready;
	input io_connPE_42_push_valid;
	input [255:0] io_connPE_42_push_bits;
	input io_connPE_42_pop_ready;
	output wire io_connPE_42_pop_valid;
	output wire io_connPE_43_push_ready;
	input io_connPE_43_push_valid;
	input [255:0] io_connPE_43_push_bits;
	input io_connPE_43_pop_ready;
	output wire io_connPE_43_pop_valid;
	output wire io_connPE_44_push_ready;
	input io_connPE_44_push_valid;
	input [255:0] io_connPE_44_push_bits;
	input io_connPE_44_pop_ready;
	output wire io_connPE_44_pop_valid;
	output wire io_connPE_45_push_ready;
	input io_connPE_45_push_valid;
	input [255:0] io_connPE_45_push_bits;
	input io_connPE_45_pop_ready;
	output wire io_connPE_45_pop_valid;
	output wire io_connPE_46_push_ready;
	input io_connPE_46_push_valid;
	input [255:0] io_connPE_46_push_bits;
	input io_connPE_46_pop_ready;
	output wire io_connPE_46_pop_valid;
	output wire io_connPE_47_push_ready;
	input io_connPE_47_push_valid;
	input [255:0] io_connPE_47_push_bits;
	input io_connPE_47_pop_ready;
	output wire io_connPE_47_pop_valid;
	output wire io_connPE_48_push_ready;
	input io_connPE_48_push_valid;
	input [255:0] io_connPE_48_push_bits;
	input io_connPE_48_pop_ready;
	output wire io_connPE_48_pop_valid;
	output wire io_connPE_49_push_ready;
	input io_connPE_49_push_valid;
	input [255:0] io_connPE_49_push_bits;
	input io_connPE_49_pop_ready;
	output wire io_connPE_49_pop_valid;
	output wire io_connPE_50_push_ready;
	input io_connPE_50_push_valid;
	input [255:0] io_connPE_50_push_bits;
	input io_connPE_50_pop_ready;
	output wire io_connPE_50_pop_valid;
	output wire io_connPE_51_push_ready;
	input io_connPE_51_push_valid;
	input [255:0] io_connPE_51_push_bits;
	input io_connPE_51_pop_ready;
	output wire io_connPE_51_pop_valid;
	output wire io_connPE_52_push_ready;
	input io_connPE_52_push_valid;
	input [255:0] io_connPE_52_push_bits;
	input io_connPE_52_pop_ready;
	output wire io_connPE_52_pop_valid;
	output wire io_connPE_53_push_ready;
	input io_connPE_53_push_valid;
	input [255:0] io_connPE_53_push_bits;
	input io_connPE_53_pop_ready;
	output wire io_connPE_53_pop_valid;
	output wire io_connPE_54_push_ready;
	input io_connPE_54_push_valid;
	input [255:0] io_connPE_54_push_bits;
	input io_connPE_54_pop_ready;
	output wire io_connPE_54_pop_valid;
	output wire io_connPE_55_push_ready;
	input io_connPE_55_push_valid;
	input [255:0] io_connPE_55_push_bits;
	input io_connPE_55_pop_ready;
	output wire io_connPE_55_pop_valid;
	output wire io_connPE_56_push_ready;
	input io_connPE_56_push_valid;
	input [255:0] io_connPE_56_push_bits;
	input io_connPE_56_pop_ready;
	output wire io_connPE_56_pop_valid;
	output wire io_connPE_57_push_ready;
	input io_connPE_57_push_valid;
	input [255:0] io_connPE_57_push_bits;
	input io_connPE_57_pop_ready;
	output wire io_connPE_57_pop_valid;
	output wire io_connPE_58_push_ready;
	input io_connPE_58_push_valid;
	input [255:0] io_connPE_58_push_bits;
	input io_connPE_58_pop_ready;
	output wire io_connPE_58_pop_valid;
	output wire io_connPE_59_push_ready;
	input io_connPE_59_push_valid;
	input [255:0] io_connPE_59_push_bits;
	input io_connPE_59_pop_ready;
	output wire io_connPE_59_pop_valid;
	output wire io_connPE_60_push_ready;
	input io_connPE_60_push_valid;
	input [255:0] io_connPE_60_push_bits;
	input io_connPE_60_pop_ready;
	output wire io_connPE_60_pop_valid;
	output wire io_connPE_61_push_ready;
	input io_connPE_61_push_valid;
	input [255:0] io_connPE_61_push_bits;
	input io_connPE_61_pop_ready;
	output wire io_connPE_61_pop_valid;
	output wire io_connPE_62_push_ready;
	input io_connPE_62_push_valid;
	input [255:0] io_connPE_62_push_bits;
	input io_connPE_62_pop_ready;
	output wire io_connPE_62_pop_valid;
	output wire io_connPE_63_push_ready;
	input io_connPE_63_push_valid;
	input [255:0] io_connPE_63_push_bits;
	input io_connPE_63_pop_ready;
	output wire io_connPE_63_pop_valid;
	input io_connVSS_0_ctrl_serveStealReq_valid;
	output wire io_connVSS_0_ctrl_serveStealReq_ready;
	input io_connVSS_0_data_availableTask_ready;
	output wire io_connVSS_0_data_availableTask_valid;
	output wire [255:0] io_connVSS_0_data_availableTask_bits;
	output wire io_connVSS_0_data_qOutTask_ready;
	input io_connVSS_0_data_qOutTask_valid;
	input [255:0] io_connVSS_0_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	wire [8:0] _taskQueues_63_io_connVec_1_currLength;
	wire _taskQueues_63_io_connVec_1_push_ready;
	wire _taskQueues_63_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_63_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_62_io_connVec_1_currLength;
	wire _taskQueues_62_io_connVec_1_push_ready;
	wire _taskQueues_62_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_62_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_61_io_connVec_1_currLength;
	wire _taskQueues_61_io_connVec_1_push_ready;
	wire _taskQueues_61_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_61_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_60_io_connVec_1_currLength;
	wire _taskQueues_60_io_connVec_1_push_ready;
	wire _taskQueues_60_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_60_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_59_io_connVec_1_currLength;
	wire _taskQueues_59_io_connVec_1_push_ready;
	wire _taskQueues_59_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_59_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_58_io_connVec_1_currLength;
	wire _taskQueues_58_io_connVec_1_push_ready;
	wire _taskQueues_58_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_58_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_57_io_connVec_1_currLength;
	wire _taskQueues_57_io_connVec_1_push_ready;
	wire _taskQueues_57_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_57_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_56_io_connVec_1_currLength;
	wire _taskQueues_56_io_connVec_1_push_ready;
	wire _taskQueues_56_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_56_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_55_io_connVec_1_currLength;
	wire _taskQueues_55_io_connVec_1_push_ready;
	wire _taskQueues_55_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_55_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_54_io_connVec_1_currLength;
	wire _taskQueues_54_io_connVec_1_push_ready;
	wire _taskQueues_54_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_54_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_53_io_connVec_1_currLength;
	wire _taskQueues_53_io_connVec_1_push_ready;
	wire _taskQueues_53_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_53_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_52_io_connVec_1_currLength;
	wire _taskQueues_52_io_connVec_1_push_ready;
	wire _taskQueues_52_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_52_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_51_io_connVec_1_currLength;
	wire _taskQueues_51_io_connVec_1_push_ready;
	wire _taskQueues_51_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_51_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_50_io_connVec_1_currLength;
	wire _taskQueues_50_io_connVec_1_push_ready;
	wire _taskQueues_50_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_50_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_49_io_connVec_1_currLength;
	wire _taskQueues_49_io_connVec_1_push_ready;
	wire _taskQueues_49_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_49_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_48_io_connVec_1_currLength;
	wire _taskQueues_48_io_connVec_1_push_ready;
	wire _taskQueues_48_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_48_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_47_io_connVec_1_currLength;
	wire _taskQueues_47_io_connVec_1_push_ready;
	wire _taskQueues_47_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_47_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_46_io_connVec_1_currLength;
	wire _taskQueues_46_io_connVec_1_push_ready;
	wire _taskQueues_46_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_46_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_45_io_connVec_1_currLength;
	wire _taskQueues_45_io_connVec_1_push_ready;
	wire _taskQueues_45_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_45_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_44_io_connVec_1_currLength;
	wire _taskQueues_44_io_connVec_1_push_ready;
	wire _taskQueues_44_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_44_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_43_io_connVec_1_currLength;
	wire _taskQueues_43_io_connVec_1_push_ready;
	wire _taskQueues_43_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_43_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_42_io_connVec_1_currLength;
	wire _taskQueues_42_io_connVec_1_push_ready;
	wire _taskQueues_42_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_42_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_41_io_connVec_1_currLength;
	wire _taskQueues_41_io_connVec_1_push_ready;
	wire _taskQueues_41_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_41_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_40_io_connVec_1_currLength;
	wire _taskQueues_40_io_connVec_1_push_ready;
	wire _taskQueues_40_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_40_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_39_io_connVec_1_currLength;
	wire _taskQueues_39_io_connVec_1_push_ready;
	wire _taskQueues_39_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_39_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_38_io_connVec_1_currLength;
	wire _taskQueues_38_io_connVec_1_push_ready;
	wire _taskQueues_38_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_38_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_37_io_connVec_1_currLength;
	wire _taskQueues_37_io_connVec_1_push_ready;
	wire _taskQueues_37_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_37_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_36_io_connVec_1_currLength;
	wire _taskQueues_36_io_connVec_1_push_ready;
	wire _taskQueues_36_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_36_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_35_io_connVec_1_currLength;
	wire _taskQueues_35_io_connVec_1_push_ready;
	wire _taskQueues_35_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_35_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_34_io_connVec_1_currLength;
	wire _taskQueues_34_io_connVec_1_push_ready;
	wire _taskQueues_34_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_34_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_33_io_connVec_1_currLength;
	wire _taskQueues_33_io_connVec_1_push_ready;
	wire _taskQueues_33_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_33_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_32_io_connVec_1_currLength;
	wire _taskQueues_32_io_connVec_1_push_ready;
	wire _taskQueues_32_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_32_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_31_io_connVec_1_currLength;
	wire _taskQueues_31_io_connVec_1_push_ready;
	wire _taskQueues_31_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_31_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_30_io_connVec_1_currLength;
	wire _taskQueues_30_io_connVec_1_push_ready;
	wire _taskQueues_30_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_30_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_29_io_connVec_1_currLength;
	wire _taskQueues_29_io_connVec_1_push_ready;
	wire _taskQueues_29_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_29_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_28_io_connVec_1_currLength;
	wire _taskQueues_28_io_connVec_1_push_ready;
	wire _taskQueues_28_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_28_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_27_io_connVec_1_currLength;
	wire _taskQueues_27_io_connVec_1_push_ready;
	wire _taskQueues_27_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_27_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_26_io_connVec_1_currLength;
	wire _taskQueues_26_io_connVec_1_push_ready;
	wire _taskQueues_26_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_26_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_25_io_connVec_1_currLength;
	wire _taskQueues_25_io_connVec_1_push_ready;
	wire _taskQueues_25_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_25_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_24_io_connVec_1_currLength;
	wire _taskQueues_24_io_connVec_1_push_ready;
	wire _taskQueues_24_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_24_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_23_io_connVec_1_currLength;
	wire _taskQueues_23_io_connVec_1_push_ready;
	wire _taskQueues_23_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_23_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_22_io_connVec_1_currLength;
	wire _taskQueues_22_io_connVec_1_push_ready;
	wire _taskQueues_22_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_22_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_21_io_connVec_1_currLength;
	wire _taskQueues_21_io_connVec_1_push_ready;
	wire _taskQueues_21_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_21_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_20_io_connVec_1_currLength;
	wire _taskQueues_20_io_connVec_1_push_ready;
	wire _taskQueues_20_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_20_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_19_io_connVec_1_currLength;
	wire _taskQueues_19_io_connVec_1_push_ready;
	wire _taskQueues_19_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_19_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_18_io_connVec_1_currLength;
	wire _taskQueues_18_io_connVec_1_push_ready;
	wire _taskQueues_18_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_18_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_17_io_connVec_1_currLength;
	wire _taskQueues_17_io_connVec_1_push_ready;
	wire _taskQueues_17_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_17_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_16_io_connVec_1_currLength;
	wire _taskQueues_16_io_connVec_1_push_ready;
	wire _taskQueues_16_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_16_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_15_io_connVec_1_currLength;
	wire _taskQueues_15_io_connVec_1_push_ready;
	wire _taskQueues_15_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_15_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_14_io_connVec_1_currLength;
	wire _taskQueues_14_io_connVec_1_push_ready;
	wire _taskQueues_14_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_14_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_13_io_connVec_1_currLength;
	wire _taskQueues_13_io_connVec_1_push_ready;
	wire _taskQueues_13_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_13_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_12_io_connVec_1_currLength;
	wire _taskQueues_12_io_connVec_1_push_ready;
	wire _taskQueues_12_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_12_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_11_io_connVec_1_currLength;
	wire _taskQueues_11_io_connVec_1_push_ready;
	wire _taskQueues_11_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_11_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_10_io_connVec_1_currLength;
	wire _taskQueues_10_io_connVec_1_push_ready;
	wire _taskQueues_10_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_10_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_9_io_connVec_1_currLength;
	wire _taskQueues_9_io_connVec_1_push_ready;
	wire _taskQueues_9_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_9_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_8_io_connVec_1_currLength;
	wire _taskQueues_8_io_connVec_1_push_ready;
	wire _taskQueues_8_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_8_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_7_io_connVec_1_currLength;
	wire _taskQueues_7_io_connVec_1_push_ready;
	wire _taskQueues_7_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_7_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_6_io_connVec_1_currLength;
	wire _taskQueues_6_io_connVec_1_push_ready;
	wire _taskQueues_6_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_6_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_5_io_connVec_1_currLength;
	wire _taskQueues_5_io_connVec_1_push_ready;
	wire _taskQueues_5_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_5_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_4_io_connVec_1_currLength;
	wire _taskQueues_4_io_connVec_1_push_ready;
	wire _taskQueues_4_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_4_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_3_io_connVec_1_currLength;
	wire _taskQueues_3_io_connVec_1_push_ready;
	wire _taskQueues_3_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_3_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_2_io_connVec_1_currLength;
	wire _taskQueues_2_io_connVec_1_push_ready;
	wire _taskQueues_2_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_2_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_1_io_connVec_1_currLength;
	wire _taskQueues_1_io_connVec_1_push_ready;
	wire _taskQueues_1_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_1_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_0_io_connVec_1_currLength;
	wire _taskQueues_0_io_connVec_1_push_ready;
	wire _taskQueues_0_io_connVec_1_pop_valid;
	wire [255:0] _taskQueues_0_io_connVec_1_pop_bits;
	wire _stealServers_63_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_63_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_63_io_connNetwork_data_availableTask_ready;
	wire _stealServers_63_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_63_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_63_io_connQ_push_valid;
	wire [255:0] _stealServers_63_io_connQ_push_bits;
	wire _stealServers_63_io_connQ_pop_ready;
	wire _stealServers_62_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_62_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_62_io_connNetwork_data_availableTask_ready;
	wire _stealServers_62_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_62_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_62_io_connQ_push_valid;
	wire [255:0] _stealServers_62_io_connQ_push_bits;
	wire _stealServers_62_io_connQ_pop_ready;
	wire _stealServers_61_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_61_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_61_io_connNetwork_data_availableTask_ready;
	wire _stealServers_61_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_61_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_61_io_connQ_push_valid;
	wire [255:0] _stealServers_61_io_connQ_push_bits;
	wire _stealServers_61_io_connQ_pop_ready;
	wire _stealServers_60_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_60_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_60_io_connNetwork_data_availableTask_ready;
	wire _stealServers_60_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_60_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_60_io_connQ_push_valid;
	wire [255:0] _stealServers_60_io_connQ_push_bits;
	wire _stealServers_60_io_connQ_pop_ready;
	wire _stealServers_59_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_59_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_59_io_connNetwork_data_availableTask_ready;
	wire _stealServers_59_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_59_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_59_io_connQ_push_valid;
	wire [255:0] _stealServers_59_io_connQ_push_bits;
	wire _stealServers_59_io_connQ_pop_ready;
	wire _stealServers_58_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_58_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_58_io_connNetwork_data_availableTask_ready;
	wire _stealServers_58_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_58_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_58_io_connQ_push_valid;
	wire [255:0] _stealServers_58_io_connQ_push_bits;
	wire _stealServers_58_io_connQ_pop_ready;
	wire _stealServers_57_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_57_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_57_io_connNetwork_data_availableTask_ready;
	wire _stealServers_57_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_57_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_57_io_connQ_push_valid;
	wire [255:0] _stealServers_57_io_connQ_push_bits;
	wire _stealServers_57_io_connQ_pop_ready;
	wire _stealServers_56_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_56_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_56_io_connNetwork_data_availableTask_ready;
	wire _stealServers_56_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_56_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_56_io_connQ_push_valid;
	wire [255:0] _stealServers_56_io_connQ_push_bits;
	wire _stealServers_56_io_connQ_pop_ready;
	wire _stealServers_55_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_55_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_55_io_connNetwork_data_availableTask_ready;
	wire _stealServers_55_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_55_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_55_io_connQ_push_valid;
	wire [255:0] _stealServers_55_io_connQ_push_bits;
	wire _stealServers_55_io_connQ_pop_ready;
	wire _stealServers_54_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_54_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_54_io_connNetwork_data_availableTask_ready;
	wire _stealServers_54_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_54_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_54_io_connQ_push_valid;
	wire [255:0] _stealServers_54_io_connQ_push_bits;
	wire _stealServers_54_io_connQ_pop_ready;
	wire _stealServers_53_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_53_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_53_io_connNetwork_data_availableTask_ready;
	wire _stealServers_53_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_53_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_53_io_connQ_push_valid;
	wire [255:0] _stealServers_53_io_connQ_push_bits;
	wire _stealServers_53_io_connQ_pop_ready;
	wire _stealServers_52_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_52_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_52_io_connNetwork_data_availableTask_ready;
	wire _stealServers_52_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_52_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_52_io_connQ_push_valid;
	wire [255:0] _stealServers_52_io_connQ_push_bits;
	wire _stealServers_52_io_connQ_pop_ready;
	wire _stealServers_51_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_51_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_51_io_connNetwork_data_availableTask_ready;
	wire _stealServers_51_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_51_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_51_io_connQ_push_valid;
	wire [255:0] _stealServers_51_io_connQ_push_bits;
	wire _stealServers_51_io_connQ_pop_ready;
	wire _stealServers_50_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_50_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_50_io_connNetwork_data_availableTask_ready;
	wire _stealServers_50_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_50_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_50_io_connQ_push_valid;
	wire [255:0] _stealServers_50_io_connQ_push_bits;
	wire _stealServers_50_io_connQ_pop_ready;
	wire _stealServers_49_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_49_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_49_io_connNetwork_data_availableTask_ready;
	wire _stealServers_49_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_49_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_49_io_connQ_push_valid;
	wire [255:0] _stealServers_49_io_connQ_push_bits;
	wire _stealServers_49_io_connQ_pop_ready;
	wire _stealServers_48_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_48_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_48_io_connNetwork_data_availableTask_ready;
	wire _stealServers_48_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_48_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_48_io_connQ_push_valid;
	wire [255:0] _stealServers_48_io_connQ_push_bits;
	wire _stealServers_48_io_connQ_pop_ready;
	wire _stealServers_47_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_47_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_47_io_connNetwork_data_availableTask_ready;
	wire _stealServers_47_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_47_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_47_io_connQ_push_valid;
	wire [255:0] _stealServers_47_io_connQ_push_bits;
	wire _stealServers_47_io_connQ_pop_ready;
	wire _stealServers_46_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_46_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_46_io_connNetwork_data_availableTask_ready;
	wire _stealServers_46_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_46_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_46_io_connQ_push_valid;
	wire [255:0] _stealServers_46_io_connQ_push_bits;
	wire _stealServers_46_io_connQ_pop_ready;
	wire _stealServers_45_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_45_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_45_io_connNetwork_data_availableTask_ready;
	wire _stealServers_45_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_45_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_45_io_connQ_push_valid;
	wire [255:0] _stealServers_45_io_connQ_push_bits;
	wire _stealServers_45_io_connQ_pop_ready;
	wire _stealServers_44_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_44_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_44_io_connNetwork_data_availableTask_ready;
	wire _stealServers_44_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_44_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_44_io_connQ_push_valid;
	wire [255:0] _stealServers_44_io_connQ_push_bits;
	wire _stealServers_44_io_connQ_pop_ready;
	wire _stealServers_43_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_43_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_43_io_connNetwork_data_availableTask_ready;
	wire _stealServers_43_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_43_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_43_io_connQ_push_valid;
	wire [255:0] _stealServers_43_io_connQ_push_bits;
	wire _stealServers_43_io_connQ_pop_ready;
	wire _stealServers_42_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_42_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_42_io_connNetwork_data_availableTask_ready;
	wire _stealServers_42_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_42_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_42_io_connQ_push_valid;
	wire [255:0] _stealServers_42_io_connQ_push_bits;
	wire _stealServers_42_io_connQ_pop_ready;
	wire _stealServers_41_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_41_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_41_io_connNetwork_data_availableTask_ready;
	wire _stealServers_41_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_41_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_41_io_connQ_push_valid;
	wire [255:0] _stealServers_41_io_connQ_push_bits;
	wire _stealServers_41_io_connQ_pop_ready;
	wire _stealServers_40_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_40_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_40_io_connNetwork_data_availableTask_ready;
	wire _stealServers_40_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_40_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_40_io_connQ_push_valid;
	wire [255:0] _stealServers_40_io_connQ_push_bits;
	wire _stealServers_40_io_connQ_pop_ready;
	wire _stealServers_39_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_39_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_39_io_connNetwork_data_availableTask_ready;
	wire _stealServers_39_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_39_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_39_io_connQ_push_valid;
	wire [255:0] _stealServers_39_io_connQ_push_bits;
	wire _stealServers_39_io_connQ_pop_ready;
	wire _stealServers_38_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_38_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_38_io_connNetwork_data_availableTask_ready;
	wire _stealServers_38_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_38_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_38_io_connQ_push_valid;
	wire [255:0] _stealServers_38_io_connQ_push_bits;
	wire _stealServers_38_io_connQ_pop_ready;
	wire _stealServers_37_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_37_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_37_io_connNetwork_data_availableTask_ready;
	wire _stealServers_37_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_37_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_37_io_connQ_push_valid;
	wire [255:0] _stealServers_37_io_connQ_push_bits;
	wire _stealServers_37_io_connQ_pop_ready;
	wire _stealServers_36_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_36_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_36_io_connNetwork_data_availableTask_ready;
	wire _stealServers_36_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_36_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_36_io_connQ_push_valid;
	wire [255:0] _stealServers_36_io_connQ_push_bits;
	wire _stealServers_36_io_connQ_pop_ready;
	wire _stealServers_35_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_35_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_35_io_connNetwork_data_availableTask_ready;
	wire _stealServers_35_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_35_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_35_io_connQ_push_valid;
	wire [255:0] _stealServers_35_io_connQ_push_bits;
	wire _stealServers_35_io_connQ_pop_ready;
	wire _stealServers_34_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_34_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_34_io_connNetwork_data_availableTask_ready;
	wire _stealServers_34_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_34_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_34_io_connQ_push_valid;
	wire [255:0] _stealServers_34_io_connQ_push_bits;
	wire _stealServers_34_io_connQ_pop_ready;
	wire _stealServers_33_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_33_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_33_io_connNetwork_data_availableTask_ready;
	wire _stealServers_33_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_33_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_33_io_connQ_push_valid;
	wire [255:0] _stealServers_33_io_connQ_push_bits;
	wire _stealServers_33_io_connQ_pop_ready;
	wire _stealServers_32_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_32_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_32_io_connNetwork_data_availableTask_ready;
	wire _stealServers_32_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_32_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_32_io_connQ_push_valid;
	wire [255:0] _stealServers_32_io_connQ_push_bits;
	wire _stealServers_32_io_connQ_pop_ready;
	wire _stealServers_31_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_31_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_31_io_connNetwork_data_availableTask_ready;
	wire _stealServers_31_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_31_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_31_io_connQ_push_valid;
	wire [255:0] _stealServers_31_io_connQ_push_bits;
	wire _stealServers_31_io_connQ_pop_ready;
	wire _stealServers_30_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_30_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_30_io_connNetwork_data_availableTask_ready;
	wire _stealServers_30_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_30_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_30_io_connQ_push_valid;
	wire [255:0] _stealServers_30_io_connQ_push_bits;
	wire _stealServers_30_io_connQ_pop_ready;
	wire _stealServers_29_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_29_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_29_io_connNetwork_data_availableTask_ready;
	wire _stealServers_29_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_29_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_29_io_connQ_push_valid;
	wire [255:0] _stealServers_29_io_connQ_push_bits;
	wire _stealServers_29_io_connQ_pop_ready;
	wire _stealServers_28_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_28_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_28_io_connNetwork_data_availableTask_ready;
	wire _stealServers_28_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_28_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_28_io_connQ_push_valid;
	wire [255:0] _stealServers_28_io_connQ_push_bits;
	wire _stealServers_28_io_connQ_pop_ready;
	wire _stealServers_27_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_27_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_27_io_connNetwork_data_availableTask_ready;
	wire _stealServers_27_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_27_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_27_io_connQ_push_valid;
	wire [255:0] _stealServers_27_io_connQ_push_bits;
	wire _stealServers_27_io_connQ_pop_ready;
	wire _stealServers_26_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_26_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_26_io_connNetwork_data_availableTask_ready;
	wire _stealServers_26_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_26_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_26_io_connQ_push_valid;
	wire [255:0] _stealServers_26_io_connQ_push_bits;
	wire _stealServers_26_io_connQ_pop_ready;
	wire _stealServers_25_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_25_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_25_io_connNetwork_data_availableTask_ready;
	wire _stealServers_25_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_25_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_25_io_connQ_push_valid;
	wire [255:0] _stealServers_25_io_connQ_push_bits;
	wire _stealServers_25_io_connQ_pop_ready;
	wire _stealServers_24_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_24_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_24_io_connNetwork_data_availableTask_ready;
	wire _stealServers_24_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_24_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_24_io_connQ_push_valid;
	wire [255:0] _stealServers_24_io_connQ_push_bits;
	wire _stealServers_24_io_connQ_pop_ready;
	wire _stealServers_23_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_23_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_23_io_connNetwork_data_availableTask_ready;
	wire _stealServers_23_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_23_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_23_io_connQ_push_valid;
	wire [255:0] _stealServers_23_io_connQ_push_bits;
	wire _stealServers_23_io_connQ_pop_ready;
	wire _stealServers_22_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_22_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_22_io_connNetwork_data_availableTask_ready;
	wire _stealServers_22_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_22_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_22_io_connQ_push_valid;
	wire [255:0] _stealServers_22_io_connQ_push_bits;
	wire _stealServers_22_io_connQ_pop_ready;
	wire _stealServers_21_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_21_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_21_io_connNetwork_data_availableTask_ready;
	wire _stealServers_21_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_21_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_21_io_connQ_push_valid;
	wire [255:0] _stealServers_21_io_connQ_push_bits;
	wire _stealServers_21_io_connQ_pop_ready;
	wire _stealServers_20_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_20_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_20_io_connNetwork_data_availableTask_ready;
	wire _stealServers_20_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_20_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_20_io_connQ_push_valid;
	wire [255:0] _stealServers_20_io_connQ_push_bits;
	wire _stealServers_20_io_connQ_pop_ready;
	wire _stealServers_19_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_19_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_19_io_connNetwork_data_availableTask_ready;
	wire _stealServers_19_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_19_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_19_io_connQ_push_valid;
	wire [255:0] _stealServers_19_io_connQ_push_bits;
	wire _stealServers_19_io_connQ_pop_ready;
	wire _stealServers_18_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_18_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_18_io_connNetwork_data_availableTask_ready;
	wire _stealServers_18_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_18_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_18_io_connQ_push_valid;
	wire [255:0] _stealServers_18_io_connQ_push_bits;
	wire _stealServers_18_io_connQ_pop_ready;
	wire _stealServers_17_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_17_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_17_io_connNetwork_data_availableTask_ready;
	wire _stealServers_17_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_17_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_17_io_connQ_push_valid;
	wire [255:0] _stealServers_17_io_connQ_push_bits;
	wire _stealServers_17_io_connQ_pop_ready;
	wire _stealServers_16_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_16_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_16_io_connNetwork_data_availableTask_ready;
	wire _stealServers_16_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_16_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_16_io_connQ_push_valid;
	wire [255:0] _stealServers_16_io_connQ_push_bits;
	wire _stealServers_16_io_connQ_pop_ready;
	wire _stealServers_15_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_15_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_15_io_connNetwork_data_availableTask_ready;
	wire _stealServers_15_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_15_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_15_io_connQ_push_valid;
	wire [255:0] _stealServers_15_io_connQ_push_bits;
	wire _stealServers_15_io_connQ_pop_ready;
	wire _stealServers_14_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_14_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_14_io_connNetwork_data_availableTask_ready;
	wire _stealServers_14_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_14_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_14_io_connQ_push_valid;
	wire [255:0] _stealServers_14_io_connQ_push_bits;
	wire _stealServers_14_io_connQ_pop_ready;
	wire _stealServers_13_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_13_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_13_io_connNetwork_data_availableTask_ready;
	wire _stealServers_13_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_13_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_13_io_connQ_push_valid;
	wire [255:0] _stealServers_13_io_connQ_push_bits;
	wire _stealServers_13_io_connQ_pop_ready;
	wire _stealServers_12_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_12_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_12_io_connNetwork_data_availableTask_ready;
	wire _stealServers_12_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_12_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_12_io_connQ_push_valid;
	wire [255:0] _stealServers_12_io_connQ_push_bits;
	wire _stealServers_12_io_connQ_pop_ready;
	wire _stealServers_11_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_11_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_11_io_connNetwork_data_availableTask_ready;
	wire _stealServers_11_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_11_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_11_io_connQ_push_valid;
	wire [255:0] _stealServers_11_io_connQ_push_bits;
	wire _stealServers_11_io_connQ_pop_ready;
	wire _stealServers_10_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_10_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_10_io_connNetwork_data_availableTask_ready;
	wire _stealServers_10_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_10_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_10_io_connQ_push_valid;
	wire [255:0] _stealServers_10_io_connQ_push_bits;
	wire _stealServers_10_io_connQ_pop_ready;
	wire _stealServers_9_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_9_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_9_io_connNetwork_data_availableTask_ready;
	wire _stealServers_9_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_9_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_9_io_connQ_push_valid;
	wire [255:0] _stealServers_9_io_connQ_push_bits;
	wire _stealServers_9_io_connQ_pop_ready;
	wire _stealServers_8_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_8_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_8_io_connNetwork_data_availableTask_ready;
	wire _stealServers_8_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_8_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_8_io_connQ_push_valid;
	wire [255:0] _stealServers_8_io_connQ_push_bits;
	wire _stealServers_8_io_connQ_pop_ready;
	wire _stealServers_7_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_7_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_7_io_connNetwork_data_availableTask_ready;
	wire _stealServers_7_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_7_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_7_io_connQ_push_valid;
	wire [255:0] _stealServers_7_io_connQ_push_bits;
	wire _stealServers_7_io_connQ_pop_ready;
	wire _stealServers_6_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_6_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_6_io_connNetwork_data_availableTask_ready;
	wire _stealServers_6_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_6_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_6_io_connQ_push_valid;
	wire [255:0] _stealServers_6_io_connQ_push_bits;
	wire _stealServers_6_io_connQ_pop_ready;
	wire _stealServers_5_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_5_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_5_io_connNetwork_data_availableTask_ready;
	wire _stealServers_5_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_5_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_5_io_connQ_push_valid;
	wire [255:0] _stealServers_5_io_connQ_push_bits;
	wire _stealServers_5_io_connQ_pop_ready;
	wire _stealServers_4_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_4_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_4_io_connNetwork_data_availableTask_ready;
	wire _stealServers_4_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_4_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_4_io_connQ_push_valid;
	wire [255:0] _stealServers_4_io_connQ_push_bits;
	wire _stealServers_4_io_connQ_pop_ready;
	wire _stealServers_3_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_3_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_3_io_connNetwork_data_availableTask_ready;
	wire _stealServers_3_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_3_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_3_io_connQ_push_valid;
	wire [255:0] _stealServers_3_io_connQ_push_bits;
	wire _stealServers_3_io_connQ_pop_ready;
	wire _stealServers_2_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_2_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_2_io_connNetwork_data_availableTask_ready;
	wire _stealServers_2_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_2_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_2_io_connQ_push_valid;
	wire [255:0] _stealServers_2_io_connQ_push_bits;
	wire _stealServers_2_io_connQ_pop_ready;
	wire _stealServers_1_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_1_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_1_io_connNetwork_data_availableTask_ready;
	wire _stealServers_1_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_1_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_1_io_connQ_push_valid;
	wire [255:0] _stealServers_1_io_connQ_push_bits;
	wire _stealServers_1_io_connQ_pop_ready;
	wire _stealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_0_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_0_io_connNetwork_data_availableTask_ready;
	wire _stealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _stealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_0_io_connQ_push_valid;
	wire [255:0] _stealServers_0_io_connQ_push_bits;
	wire _stealServers_0_io_connQ_pop_ready;
	wire _stealNet_io_connSS_1_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_1_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_1_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_1_data_availableTask_bits;
	wire _stealNet_io_connSS_1_data_qOutTask_ready;
	wire _stealNet_io_connSS_2_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_2_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_2_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_2_data_availableTask_bits;
	wire _stealNet_io_connSS_2_data_qOutTask_ready;
	wire _stealNet_io_connSS_3_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_3_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_3_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_3_data_availableTask_bits;
	wire _stealNet_io_connSS_3_data_qOutTask_ready;
	wire _stealNet_io_connSS_4_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_4_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_4_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_4_data_availableTask_bits;
	wire _stealNet_io_connSS_4_data_qOutTask_ready;
	wire _stealNet_io_connSS_5_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_5_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_5_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_5_data_availableTask_bits;
	wire _stealNet_io_connSS_5_data_qOutTask_ready;
	wire _stealNet_io_connSS_6_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_6_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_6_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_6_data_availableTask_bits;
	wire _stealNet_io_connSS_6_data_qOutTask_ready;
	wire _stealNet_io_connSS_7_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_7_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_7_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_7_data_availableTask_bits;
	wire _stealNet_io_connSS_7_data_qOutTask_ready;
	wire _stealNet_io_connSS_8_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_8_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_8_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_8_data_availableTask_bits;
	wire _stealNet_io_connSS_8_data_qOutTask_ready;
	wire _stealNet_io_connSS_9_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_9_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_9_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_9_data_availableTask_bits;
	wire _stealNet_io_connSS_9_data_qOutTask_ready;
	wire _stealNet_io_connSS_10_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_10_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_10_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_10_data_availableTask_bits;
	wire _stealNet_io_connSS_10_data_qOutTask_ready;
	wire _stealNet_io_connSS_11_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_11_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_11_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_11_data_availableTask_bits;
	wire _stealNet_io_connSS_11_data_qOutTask_ready;
	wire _stealNet_io_connSS_12_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_12_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_12_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_12_data_availableTask_bits;
	wire _stealNet_io_connSS_12_data_qOutTask_ready;
	wire _stealNet_io_connSS_13_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_13_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_13_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_13_data_availableTask_bits;
	wire _stealNet_io_connSS_13_data_qOutTask_ready;
	wire _stealNet_io_connSS_14_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_14_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_14_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_14_data_availableTask_bits;
	wire _stealNet_io_connSS_14_data_qOutTask_ready;
	wire _stealNet_io_connSS_15_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_15_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_15_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_15_data_availableTask_bits;
	wire _stealNet_io_connSS_15_data_qOutTask_ready;
	wire _stealNet_io_connSS_16_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_16_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_16_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_16_data_availableTask_bits;
	wire _stealNet_io_connSS_16_data_qOutTask_ready;
	wire _stealNet_io_connSS_17_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_17_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_17_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_17_data_availableTask_bits;
	wire _stealNet_io_connSS_17_data_qOutTask_ready;
	wire _stealNet_io_connSS_18_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_18_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_18_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_18_data_availableTask_bits;
	wire _stealNet_io_connSS_18_data_qOutTask_ready;
	wire _stealNet_io_connSS_19_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_19_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_19_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_19_data_availableTask_bits;
	wire _stealNet_io_connSS_19_data_qOutTask_ready;
	wire _stealNet_io_connSS_20_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_20_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_20_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_20_data_availableTask_bits;
	wire _stealNet_io_connSS_20_data_qOutTask_ready;
	wire _stealNet_io_connSS_21_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_21_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_21_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_21_data_availableTask_bits;
	wire _stealNet_io_connSS_21_data_qOutTask_ready;
	wire _stealNet_io_connSS_22_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_22_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_22_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_22_data_availableTask_bits;
	wire _stealNet_io_connSS_22_data_qOutTask_ready;
	wire _stealNet_io_connSS_23_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_23_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_23_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_23_data_availableTask_bits;
	wire _stealNet_io_connSS_23_data_qOutTask_ready;
	wire _stealNet_io_connSS_24_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_24_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_24_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_24_data_availableTask_bits;
	wire _stealNet_io_connSS_24_data_qOutTask_ready;
	wire _stealNet_io_connSS_25_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_25_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_25_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_25_data_availableTask_bits;
	wire _stealNet_io_connSS_25_data_qOutTask_ready;
	wire _stealNet_io_connSS_26_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_26_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_26_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_26_data_availableTask_bits;
	wire _stealNet_io_connSS_26_data_qOutTask_ready;
	wire _stealNet_io_connSS_27_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_27_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_27_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_27_data_availableTask_bits;
	wire _stealNet_io_connSS_27_data_qOutTask_ready;
	wire _stealNet_io_connSS_28_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_28_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_28_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_28_data_availableTask_bits;
	wire _stealNet_io_connSS_28_data_qOutTask_ready;
	wire _stealNet_io_connSS_29_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_29_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_29_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_29_data_availableTask_bits;
	wire _stealNet_io_connSS_29_data_qOutTask_ready;
	wire _stealNet_io_connSS_30_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_30_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_30_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_30_data_availableTask_bits;
	wire _stealNet_io_connSS_30_data_qOutTask_ready;
	wire _stealNet_io_connSS_31_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_31_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_31_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_31_data_availableTask_bits;
	wire _stealNet_io_connSS_31_data_qOutTask_ready;
	wire _stealNet_io_connSS_32_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_32_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_32_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_32_data_availableTask_bits;
	wire _stealNet_io_connSS_32_data_qOutTask_ready;
	wire _stealNet_io_connSS_33_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_33_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_33_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_33_data_availableTask_bits;
	wire _stealNet_io_connSS_33_data_qOutTask_ready;
	wire _stealNet_io_connSS_34_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_34_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_34_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_34_data_availableTask_bits;
	wire _stealNet_io_connSS_34_data_qOutTask_ready;
	wire _stealNet_io_connSS_35_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_35_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_35_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_35_data_availableTask_bits;
	wire _stealNet_io_connSS_35_data_qOutTask_ready;
	wire _stealNet_io_connSS_36_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_36_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_36_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_36_data_availableTask_bits;
	wire _stealNet_io_connSS_36_data_qOutTask_ready;
	wire _stealNet_io_connSS_37_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_37_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_37_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_37_data_availableTask_bits;
	wire _stealNet_io_connSS_37_data_qOutTask_ready;
	wire _stealNet_io_connSS_38_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_38_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_38_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_38_data_availableTask_bits;
	wire _stealNet_io_connSS_38_data_qOutTask_ready;
	wire _stealNet_io_connSS_39_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_39_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_39_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_39_data_availableTask_bits;
	wire _stealNet_io_connSS_39_data_qOutTask_ready;
	wire _stealNet_io_connSS_40_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_40_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_40_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_40_data_availableTask_bits;
	wire _stealNet_io_connSS_40_data_qOutTask_ready;
	wire _stealNet_io_connSS_41_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_41_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_41_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_41_data_availableTask_bits;
	wire _stealNet_io_connSS_41_data_qOutTask_ready;
	wire _stealNet_io_connSS_42_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_42_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_42_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_42_data_availableTask_bits;
	wire _stealNet_io_connSS_42_data_qOutTask_ready;
	wire _stealNet_io_connSS_43_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_43_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_43_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_43_data_availableTask_bits;
	wire _stealNet_io_connSS_43_data_qOutTask_ready;
	wire _stealNet_io_connSS_44_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_44_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_44_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_44_data_availableTask_bits;
	wire _stealNet_io_connSS_44_data_qOutTask_ready;
	wire _stealNet_io_connSS_45_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_45_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_45_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_45_data_availableTask_bits;
	wire _stealNet_io_connSS_45_data_qOutTask_ready;
	wire _stealNet_io_connSS_46_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_46_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_46_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_46_data_availableTask_bits;
	wire _stealNet_io_connSS_46_data_qOutTask_ready;
	wire _stealNet_io_connSS_47_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_47_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_47_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_47_data_availableTask_bits;
	wire _stealNet_io_connSS_47_data_qOutTask_ready;
	wire _stealNet_io_connSS_48_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_48_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_48_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_48_data_availableTask_bits;
	wire _stealNet_io_connSS_48_data_qOutTask_ready;
	wire _stealNet_io_connSS_49_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_49_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_49_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_49_data_availableTask_bits;
	wire _stealNet_io_connSS_49_data_qOutTask_ready;
	wire _stealNet_io_connSS_50_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_50_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_50_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_50_data_availableTask_bits;
	wire _stealNet_io_connSS_50_data_qOutTask_ready;
	wire _stealNet_io_connSS_51_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_51_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_51_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_51_data_availableTask_bits;
	wire _stealNet_io_connSS_51_data_qOutTask_ready;
	wire _stealNet_io_connSS_52_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_52_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_52_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_52_data_availableTask_bits;
	wire _stealNet_io_connSS_52_data_qOutTask_ready;
	wire _stealNet_io_connSS_53_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_53_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_53_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_53_data_availableTask_bits;
	wire _stealNet_io_connSS_53_data_qOutTask_ready;
	wire _stealNet_io_connSS_54_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_54_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_54_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_54_data_availableTask_bits;
	wire _stealNet_io_connSS_54_data_qOutTask_ready;
	wire _stealNet_io_connSS_55_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_55_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_55_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_55_data_availableTask_bits;
	wire _stealNet_io_connSS_55_data_qOutTask_ready;
	wire _stealNet_io_connSS_56_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_56_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_56_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_56_data_availableTask_bits;
	wire _stealNet_io_connSS_56_data_qOutTask_ready;
	wire _stealNet_io_connSS_57_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_57_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_57_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_57_data_availableTask_bits;
	wire _stealNet_io_connSS_57_data_qOutTask_ready;
	wire _stealNet_io_connSS_58_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_58_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_58_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_58_data_availableTask_bits;
	wire _stealNet_io_connSS_58_data_qOutTask_ready;
	wire _stealNet_io_connSS_59_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_59_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_59_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_59_data_availableTask_bits;
	wire _stealNet_io_connSS_59_data_qOutTask_ready;
	wire _stealNet_io_connSS_60_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_60_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_60_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_60_data_availableTask_bits;
	wire _stealNet_io_connSS_60_data_qOutTask_ready;
	wire _stealNet_io_connSS_61_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_61_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_61_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_61_data_availableTask_bits;
	wire _stealNet_io_connSS_61_data_qOutTask_ready;
	wire _stealNet_io_connSS_62_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_62_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_62_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_62_data_availableTask_bits;
	wire _stealNet_io_connSS_62_data_qOutTask_ready;
	wire _stealNet_io_connSS_63_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_63_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_63_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_63_data_availableTask_bits;
	wire _stealNet_io_connSS_63_data_qOutTask_ready;
	wire _stealNet_io_connSS_64_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_64_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_64_data_availableTask_valid;
	wire [255:0] _stealNet_io_connSS_64_data_availableTask_bits;
	wire _stealNet_io_connSS_64_data_qOutTask_ready;
	SchedulerNetwork stealNet(
		.clock(clock),
		.reset(reset),
		.io_connSS_0_ctrl_serveStealReq_valid(io_connVSS_0_ctrl_serveStealReq_valid),
		.io_connSS_0_ctrl_serveStealReq_ready(io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connSS_0_data_availableTask_ready(io_connVSS_0_data_availableTask_ready),
		.io_connSS_0_data_availableTask_valid(io_connVSS_0_data_availableTask_valid),
		.io_connSS_0_data_availableTask_bits(io_connVSS_0_data_availableTask_bits),
		.io_connSS_0_data_qOutTask_ready(io_connVSS_0_data_qOutTask_ready),
		.io_connSS_0_data_qOutTask_valid(io_connVSS_0_data_qOutTask_valid),
		.io_connSS_0_data_qOutTask_bits(io_connVSS_0_data_qOutTask_bits),
		.io_connSS_1_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_1_ctrl_serveStealReq_ready(_stealNet_io_connSS_1_ctrl_serveStealReq_ready),
		.io_connSS_1_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_1_ctrl_stealReq_ready(_stealNet_io_connSS_1_ctrl_stealReq_ready),
		.io_connSS_1_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connSS_1_data_availableTask_valid(_stealNet_io_connSS_1_data_availableTask_valid),
		.io_connSS_1_data_availableTask_bits(_stealNet_io_connSS_1_data_availableTask_bits),
		.io_connSS_1_data_qOutTask_ready(_stealNet_io_connSS_1_data_qOutTask_ready),
		.io_connSS_1_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connSS_1_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connSS_2_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_2_ctrl_serveStealReq_ready(_stealNet_io_connSS_2_ctrl_serveStealReq_ready),
		.io_connSS_2_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_2_ctrl_stealReq_ready(_stealNet_io_connSS_2_ctrl_stealReq_ready),
		.io_connSS_2_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connSS_2_data_availableTask_valid(_stealNet_io_connSS_2_data_availableTask_valid),
		.io_connSS_2_data_availableTask_bits(_stealNet_io_connSS_2_data_availableTask_bits),
		.io_connSS_2_data_qOutTask_ready(_stealNet_io_connSS_2_data_qOutTask_ready),
		.io_connSS_2_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connSS_2_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connSS_3_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_3_ctrl_serveStealReq_ready(_stealNet_io_connSS_3_ctrl_serveStealReq_ready),
		.io_connSS_3_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_3_ctrl_stealReq_ready(_stealNet_io_connSS_3_ctrl_stealReq_ready),
		.io_connSS_3_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connSS_3_data_availableTask_valid(_stealNet_io_connSS_3_data_availableTask_valid),
		.io_connSS_3_data_availableTask_bits(_stealNet_io_connSS_3_data_availableTask_bits),
		.io_connSS_3_data_qOutTask_ready(_stealNet_io_connSS_3_data_qOutTask_ready),
		.io_connSS_3_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connSS_3_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connSS_4_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_4_ctrl_serveStealReq_ready(_stealNet_io_connSS_4_ctrl_serveStealReq_ready),
		.io_connSS_4_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_4_ctrl_stealReq_ready(_stealNet_io_connSS_4_ctrl_stealReq_ready),
		.io_connSS_4_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connSS_4_data_availableTask_valid(_stealNet_io_connSS_4_data_availableTask_valid),
		.io_connSS_4_data_availableTask_bits(_stealNet_io_connSS_4_data_availableTask_bits),
		.io_connSS_4_data_qOutTask_ready(_stealNet_io_connSS_4_data_qOutTask_ready),
		.io_connSS_4_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connSS_4_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connSS_5_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_5_ctrl_serveStealReq_ready(_stealNet_io_connSS_5_ctrl_serveStealReq_ready),
		.io_connSS_5_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_5_ctrl_stealReq_ready(_stealNet_io_connSS_5_ctrl_stealReq_ready),
		.io_connSS_5_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connSS_5_data_availableTask_valid(_stealNet_io_connSS_5_data_availableTask_valid),
		.io_connSS_5_data_availableTask_bits(_stealNet_io_connSS_5_data_availableTask_bits),
		.io_connSS_5_data_qOutTask_ready(_stealNet_io_connSS_5_data_qOutTask_ready),
		.io_connSS_5_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connSS_5_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connSS_6_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_6_ctrl_serveStealReq_ready(_stealNet_io_connSS_6_ctrl_serveStealReq_ready),
		.io_connSS_6_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_6_ctrl_stealReq_ready(_stealNet_io_connSS_6_ctrl_stealReq_ready),
		.io_connSS_6_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connSS_6_data_availableTask_valid(_stealNet_io_connSS_6_data_availableTask_valid),
		.io_connSS_6_data_availableTask_bits(_stealNet_io_connSS_6_data_availableTask_bits),
		.io_connSS_6_data_qOutTask_ready(_stealNet_io_connSS_6_data_qOutTask_ready),
		.io_connSS_6_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connSS_6_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connSS_7_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_7_ctrl_serveStealReq_ready(_stealNet_io_connSS_7_ctrl_serveStealReq_ready),
		.io_connSS_7_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_7_ctrl_stealReq_ready(_stealNet_io_connSS_7_ctrl_stealReq_ready),
		.io_connSS_7_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connSS_7_data_availableTask_valid(_stealNet_io_connSS_7_data_availableTask_valid),
		.io_connSS_7_data_availableTask_bits(_stealNet_io_connSS_7_data_availableTask_bits),
		.io_connSS_7_data_qOutTask_ready(_stealNet_io_connSS_7_data_qOutTask_ready),
		.io_connSS_7_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connSS_7_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connSS_8_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_8_ctrl_serveStealReq_ready(_stealNet_io_connSS_8_ctrl_serveStealReq_ready),
		.io_connSS_8_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_8_ctrl_stealReq_ready(_stealNet_io_connSS_8_ctrl_stealReq_ready),
		.io_connSS_8_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connSS_8_data_availableTask_valid(_stealNet_io_connSS_8_data_availableTask_valid),
		.io_connSS_8_data_availableTask_bits(_stealNet_io_connSS_8_data_availableTask_bits),
		.io_connSS_8_data_qOutTask_ready(_stealNet_io_connSS_8_data_qOutTask_ready),
		.io_connSS_8_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connSS_8_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connSS_9_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_9_ctrl_serveStealReq_ready(_stealNet_io_connSS_9_ctrl_serveStealReq_ready),
		.io_connSS_9_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_9_ctrl_stealReq_ready(_stealNet_io_connSS_9_ctrl_stealReq_ready),
		.io_connSS_9_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connSS_9_data_availableTask_valid(_stealNet_io_connSS_9_data_availableTask_valid),
		.io_connSS_9_data_availableTask_bits(_stealNet_io_connSS_9_data_availableTask_bits),
		.io_connSS_9_data_qOutTask_ready(_stealNet_io_connSS_9_data_qOutTask_ready),
		.io_connSS_9_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connSS_9_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connSS_10_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_10_ctrl_serveStealReq_ready(_stealNet_io_connSS_10_ctrl_serveStealReq_ready),
		.io_connSS_10_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_10_ctrl_stealReq_ready(_stealNet_io_connSS_10_ctrl_stealReq_ready),
		.io_connSS_10_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connSS_10_data_availableTask_valid(_stealNet_io_connSS_10_data_availableTask_valid),
		.io_connSS_10_data_availableTask_bits(_stealNet_io_connSS_10_data_availableTask_bits),
		.io_connSS_10_data_qOutTask_ready(_stealNet_io_connSS_10_data_qOutTask_ready),
		.io_connSS_10_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connSS_10_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connSS_11_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_11_ctrl_serveStealReq_ready(_stealNet_io_connSS_11_ctrl_serveStealReq_ready),
		.io_connSS_11_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_11_ctrl_stealReq_ready(_stealNet_io_connSS_11_ctrl_stealReq_ready),
		.io_connSS_11_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connSS_11_data_availableTask_valid(_stealNet_io_connSS_11_data_availableTask_valid),
		.io_connSS_11_data_availableTask_bits(_stealNet_io_connSS_11_data_availableTask_bits),
		.io_connSS_11_data_qOutTask_ready(_stealNet_io_connSS_11_data_qOutTask_ready),
		.io_connSS_11_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connSS_11_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connSS_12_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_12_ctrl_serveStealReq_ready(_stealNet_io_connSS_12_ctrl_serveStealReq_ready),
		.io_connSS_12_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_12_ctrl_stealReq_ready(_stealNet_io_connSS_12_ctrl_stealReq_ready),
		.io_connSS_12_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connSS_12_data_availableTask_valid(_stealNet_io_connSS_12_data_availableTask_valid),
		.io_connSS_12_data_availableTask_bits(_stealNet_io_connSS_12_data_availableTask_bits),
		.io_connSS_12_data_qOutTask_ready(_stealNet_io_connSS_12_data_qOutTask_ready),
		.io_connSS_12_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connSS_12_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connSS_13_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_13_ctrl_serveStealReq_ready(_stealNet_io_connSS_13_ctrl_serveStealReq_ready),
		.io_connSS_13_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_13_ctrl_stealReq_ready(_stealNet_io_connSS_13_ctrl_stealReq_ready),
		.io_connSS_13_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connSS_13_data_availableTask_valid(_stealNet_io_connSS_13_data_availableTask_valid),
		.io_connSS_13_data_availableTask_bits(_stealNet_io_connSS_13_data_availableTask_bits),
		.io_connSS_13_data_qOutTask_ready(_stealNet_io_connSS_13_data_qOutTask_ready),
		.io_connSS_13_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connSS_13_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connSS_14_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_14_ctrl_serveStealReq_ready(_stealNet_io_connSS_14_ctrl_serveStealReq_ready),
		.io_connSS_14_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_14_ctrl_stealReq_ready(_stealNet_io_connSS_14_ctrl_stealReq_ready),
		.io_connSS_14_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connSS_14_data_availableTask_valid(_stealNet_io_connSS_14_data_availableTask_valid),
		.io_connSS_14_data_availableTask_bits(_stealNet_io_connSS_14_data_availableTask_bits),
		.io_connSS_14_data_qOutTask_ready(_stealNet_io_connSS_14_data_qOutTask_ready),
		.io_connSS_14_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connSS_14_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connSS_15_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_15_ctrl_serveStealReq_ready(_stealNet_io_connSS_15_ctrl_serveStealReq_ready),
		.io_connSS_15_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_15_ctrl_stealReq_ready(_stealNet_io_connSS_15_ctrl_stealReq_ready),
		.io_connSS_15_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connSS_15_data_availableTask_valid(_stealNet_io_connSS_15_data_availableTask_valid),
		.io_connSS_15_data_availableTask_bits(_stealNet_io_connSS_15_data_availableTask_bits),
		.io_connSS_15_data_qOutTask_ready(_stealNet_io_connSS_15_data_qOutTask_ready),
		.io_connSS_15_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connSS_15_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connSS_16_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_16_ctrl_serveStealReq_ready(_stealNet_io_connSS_16_ctrl_serveStealReq_ready),
		.io_connSS_16_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_16_ctrl_stealReq_ready(_stealNet_io_connSS_16_ctrl_stealReq_ready),
		.io_connSS_16_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connSS_16_data_availableTask_valid(_stealNet_io_connSS_16_data_availableTask_valid),
		.io_connSS_16_data_availableTask_bits(_stealNet_io_connSS_16_data_availableTask_bits),
		.io_connSS_16_data_qOutTask_ready(_stealNet_io_connSS_16_data_qOutTask_ready),
		.io_connSS_16_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connSS_16_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connSS_17_ctrl_serveStealReq_valid(_stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_17_ctrl_serveStealReq_ready(_stealNet_io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_17_ctrl_stealReq_valid(_stealServers_16_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_17_ctrl_stealReq_ready(_stealNet_io_connSS_17_ctrl_stealReq_ready),
		.io_connSS_17_data_availableTask_ready(_stealServers_16_io_connNetwork_data_availableTask_ready),
		.io_connSS_17_data_availableTask_valid(_stealNet_io_connSS_17_data_availableTask_valid),
		.io_connSS_17_data_availableTask_bits(_stealNet_io_connSS_17_data_availableTask_bits),
		.io_connSS_17_data_qOutTask_ready(_stealNet_io_connSS_17_data_qOutTask_ready),
		.io_connSS_17_data_qOutTask_valid(_stealServers_16_io_connNetwork_data_qOutTask_valid),
		.io_connSS_17_data_qOutTask_bits(_stealServers_16_io_connNetwork_data_qOutTask_bits),
		.io_connSS_18_ctrl_serveStealReq_valid(_stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_18_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_18_ctrl_stealReq_valid(_stealServers_17_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_18_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connSS_18_data_availableTask_ready(_stealServers_17_io_connNetwork_data_availableTask_ready),
		.io_connSS_18_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connSS_18_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connSS_18_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connSS_18_data_qOutTask_valid(_stealServers_17_io_connNetwork_data_qOutTask_valid),
		.io_connSS_18_data_qOutTask_bits(_stealServers_17_io_connNetwork_data_qOutTask_bits),
		.io_connSS_19_ctrl_serveStealReq_valid(_stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_19_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_19_ctrl_stealReq_valid(_stealServers_18_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_19_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connSS_19_data_availableTask_ready(_stealServers_18_io_connNetwork_data_availableTask_ready),
		.io_connSS_19_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connSS_19_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connSS_19_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connSS_19_data_qOutTask_valid(_stealServers_18_io_connNetwork_data_qOutTask_valid),
		.io_connSS_19_data_qOutTask_bits(_stealServers_18_io_connNetwork_data_qOutTask_bits),
		.io_connSS_20_ctrl_serveStealReq_valid(_stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_20_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_20_ctrl_stealReq_valid(_stealServers_19_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_20_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connSS_20_data_availableTask_ready(_stealServers_19_io_connNetwork_data_availableTask_ready),
		.io_connSS_20_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connSS_20_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connSS_20_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connSS_20_data_qOutTask_valid(_stealServers_19_io_connNetwork_data_qOutTask_valid),
		.io_connSS_20_data_qOutTask_bits(_stealServers_19_io_connNetwork_data_qOutTask_bits),
		.io_connSS_21_ctrl_serveStealReq_valid(_stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_21_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_21_ctrl_stealReq_valid(_stealServers_20_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_21_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connSS_21_data_availableTask_ready(_stealServers_20_io_connNetwork_data_availableTask_ready),
		.io_connSS_21_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connSS_21_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connSS_21_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connSS_21_data_qOutTask_valid(_stealServers_20_io_connNetwork_data_qOutTask_valid),
		.io_connSS_21_data_qOutTask_bits(_stealServers_20_io_connNetwork_data_qOutTask_bits),
		.io_connSS_22_ctrl_serveStealReq_valid(_stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_22_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_22_ctrl_stealReq_valid(_stealServers_21_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_22_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connSS_22_data_availableTask_ready(_stealServers_21_io_connNetwork_data_availableTask_ready),
		.io_connSS_22_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connSS_22_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connSS_22_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connSS_22_data_qOutTask_valid(_stealServers_21_io_connNetwork_data_qOutTask_valid),
		.io_connSS_22_data_qOutTask_bits(_stealServers_21_io_connNetwork_data_qOutTask_bits),
		.io_connSS_23_ctrl_serveStealReq_valid(_stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_23_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_23_ctrl_stealReq_valid(_stealServers_22_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_23_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connSS_23_data_availableTask_ready(_stealServers_22_io_connNetwork_data_availableTask_ready),
		.io_connSS_23_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connSS_23_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connSS_23_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connSS_23_data_qOutTask_valid(_stealServers_22_io_connNetwork_data_qOutTask_valid),
		.io_connSS_23_data_qOutTask_bits(_stealServers_22_io_connNetwork_data_qOutTask_bits),
		.io_connSS_24_ctrl_serveStealReq_valid(_stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_24_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_24_ctrl_stealReq_valid(_stealServers_23_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_24_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connSS_24_data_availableTask_ready(_stealServers_23_io_connNetwork_data_availableTask_ready),
		.io_connSS_24_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connSS_24_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connSS_24_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connSS_24_data_qOutTask_valid(_stealServers_23_io_connNetwork_data_qOutTask_valid),
		.io_connSS_24_data_qOutTask_bits(_stealServers_23_io_connNetwork_data_qOutTask_bits),
		.io_connSS_25_ctrl_serveStealReq_valid(_stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_25_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_25_ctrl_stealReq_valid(_stealServers_24_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_25_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connSS_25_data_availableTask_ready(_stealServers_24_io_connNetwork_data_availableTask_ready),
		.io_connSS_25_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connSS_25_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connSS_25_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connSS_25_data_qOutTask_valid(_stealServers_24_io_connNetwork_data_qOutTask_valid),
		.io_connSS_25_data_qOutTask_bits(_stealServers_24_io_connNetwork_data_qOutTask_bits),
		.io_connSS_26_ctrl_serveStealReq_valid(_stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_26_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_26_ctrl_stealReq_valid(_stealServers_25_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_26_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connSS_26_data_availableTask_ready(_stealServers_25_io_connNetwork_data_availableTask_ready),
		.io_connSS_26_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connSS_26_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connSS_26_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connSS_26_data_qOutTask_valid(_stealServers_25_io_connNetwork_data_qOutTask_valid),
		.io_connSS_26_data_qOutTask_bits(_stealServers_25_io_connNetwork_data_qOutTask_bits),
		.io_connSS_27_ctrl_serveStealReq_valid(_stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_27_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_27_ctrl_stealReq_valid(_stealServers_26_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_27_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connSS_27_data_availableTask_ready(_stealServers_26_io_connNetwork_data_availableTask_ready),
		.io_connSS_27_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connSS_27_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connSS_27_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connSS_27_data_qOutTask_valid(_stealServers_26_io_connNetwork_data_qOutTask_valid),
		.io_connSS_27_data_qOutTask_bits(_stealServers_26_io_connNetwork_data_qOutTask_bits),
		.io_connSS_28_ctrl_serveStealReq_valid(_stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_28_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_28_ctrl_stealReq_valid(_stealServers_27_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_28_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connSS_28_data_availableTask_ready(_stealServers_27_io_connNetwork_data_availableTask_ready),
		.io_connSS_28_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connSS_28_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connSS_28_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connSS_28_data_qOutTask_valid(_stealServers_27_io_connNetwork_data_qOutTask_valid),
		.io_connSS_28_data_qOutTask_bits(_stealServers_27_io_connNetwork_data_qOutTask_bits),
		.io_connSS_29_ctrl_serveStealReq_valid(_stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_29_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_29_ctrl_stealReq_valid(_stealServers_28_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_29_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connSS_29_data_availableTask_ready(_stealServers_28_io_connNetwork_data_availableTask_ready),
		.io_connSS_29_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connSS_29_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connSS_29_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connSS_29_data_qOutTask_valid(_stealServers_28_io_connNetwork_data_qOutTask_valid),
		.io_connSS_29_data_qOutTask_bits(_stealServers_28_io_connNetwork_data_qOutTask_bits),
		.io_connSS_30_ctrl_serveStealReq_valid(_stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_30_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_30_ctrl_stealReq_valid(_stealServers_29_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_30_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connSS_30_data_availableTask_ready(_stealServers_29_io_connNetwork_data_availableTask_ready),
		.io_connSS_30_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connSS_30_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connSS_30_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connSS_30_data_qOutTask_valid(_stealServers_29_io_connNetwork_data_qOutTask_valid),
		.io_connSS_30_data_qOutTask_bits(_stealServers_29_io_connNetwork_data_qOutTask_bits),
		.io_connSS_31_ctrl_serveStealReq_valid(_stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_31_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_31_ctrl_stealReq_valid(_stealServers_30_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_31_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connSS_31_data_availableTask_ready(_stealServers_30_io_connNetwork_data_availableTask_ready),
		.io_connSS_31_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connSS_31_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connSS_31_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connSS_31_data_qOutTask_valid(_stealServers_30_io_connNetwork_data_qOutTask_valid),
		.io_connSS_31_data_qOutTask_bits(_stealServers_30_io_connNetwork_data_qOutTask_bits),
		.io_connSS_32_ctrl_serveStealReq_valid(_stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_32_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_32_ctrl_stealReq_valid(_stealServers_31_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_32_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connSS_32_data_availableTask_ready(_stealServers_31_io_connNetwork_data_availableTask_ready),
		.io_connSS_32_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connSS_32_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connSS_32_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connSS_32_data_qOutTask_valid(_stealServers_31_io_connNetwork_data_qOutTask_valid),
		.io_connSS_32_data_qOutTask_bits(_stealServers_31_io_connNetwork_data_qOutTask_bits),
		.io_connSS_33_ctrl_serveStealReq_valid(_stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_33_ctrl_serveStealReq_ready(_stealNet_io_connSS_33_ctrl_serveStealReq_ready),
		.io_connSS_33_ctrl_stealReq_valid(_stealServers_32_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_33_ctrl_stealReq_ready(_stealNet_io_connSS_33_ctrl_stealReq_ready),
		.io_connSS_33_data_availableTask_ready(_stealServers_32_io_connNetwork_data_availableTask_ready),
		.io_connSS_33_data_availableTask_valid(_stealNet_io_connSS_33_data_availableTask_valid),
		.io_connSS_33_data_availableTask_bits(_stealNet_io_connSS_33_data_availableTask_bits),
		.io_connSS_33_data_qOutTask_ready(_stealNet_io_connSS_33_data_qOutTask_ready),
		.io_connSS_33_data_qOutTask_valid(_stealServers_32_io_connNetwork_data_qOutTask_valid),
		.io_connSS_33_data_qOutTask_bits(_stealServers_32_io_connNetwork_data_qOutTask_bits),
		.io_connSS_34_ctrl_serveStealReq_valid(_stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_34_ctrl_serveStealReq_ready(_stealNet_io_connSS_34_ctrl_serveStealReq_ready),
		.io_connSS_34_ctrl_stealReq_valid(_stealServers_33_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_34_ctrl_stealReq_ready(_stealNet_io_connSS_34_ctrl_stealReq_ready),
		.io_connSS_34_data_availableTask_ready(_stealServers_33_io_connNetwork_data_availableTask_ready),
		.io_connSS_34_data_availableTask_valid(_stealNet_io_connSS_34_data_availableTask_valid),
		.io_connSS_34_data_availableTask_bits(_stealNet_io_connSS_34_data_availableTask_bits),
		.io_connSS_34_data_qOutTask_ready(_stealNet_io_connSS_34_data_qOutTask_ready),
		.io_connSS_34_data_qOutTask_valid(_stealServers_33_io_connNetwork_data_qOutTask_valid),
		.io_connSS_34_data_qOutTask_bits(_stealServers_33_io_connNetwork_data_qOutTask_bits),
		.io_connSS_35_ctrl_serveStealReq_valid(_stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_35_ctrl_serveStealReq_ready(_stealNet_io_connSS_35_ctrl_serveStealReq_ready),
		.io_connSS_35_ctrl_stealReq_valid(_stealServers_34_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_35_ctrl_stealReq_ready(_stealNet_io_connSS_35_ctrl_stealReq_ready),
		.io_connSS_35_data_availableTask_ready(_stealServers_34_io_connNetwork_data_availableTask_ready),
		.io_connSS_35_data_availableTask_valid(_stealNet_io_connSS_35_data_availableTask_valid),
		.io_connSS_35_data_availableTask_bits(_stealNet_io_connSS_35_data_availableTask_bits),
		.io_connSS_35_data_qOutTask_ready(_stealNet_io_connSS_35_data_qOutTask_ready),
		.io_connSS_35_data_qOutTask_valid(_stealServers_34_io_connNetwork_data_qOutTask_valid),
		.io_connSS_35_data_qOutTask_bits(_stealServers_34_io_connNetwork_data_qOutTask_bits),
		.io_connSS_36_ctrl_serveStealReq_valid(_stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_36_ctrl_serveStealReq_ready(_stealNet_io_connSS_36_ctrl_serveStealReq_ready),
		.io_connSS_36_ctrl_stealReq_valid(_stealServers_35_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_36_ctrl_stealReq_ready(_stealNet_io_connSS_36_ctrl_stealReq_ready),
		.io_connSS_36_data_availableTask_ready(_stealServers_35_io_connNetwork_data_availableTask_ready),
		.io_connSS_36_data_availableTask_valid(_stealNet_io_connSS_36_data_availableTask_valid),
		.io_connSS_36_data_availableTask_bits(_stealNet_io_connSS_36_data_availableTask_bits),
		.io_connSS_36_data_qOutTask_ready(_stealNet_io_connSS_36_data_qOutTask_ready),
		.io_connSS_36_data_qOutTask_valid(_stealServers_35_io_connNetwork_data_qOutTask_valid),
		.io_connSS_36_data_qOutTask_bits(_stealServers_35_io_connNetwork_data_qOutTask_bits),
		.io_connSS_37_ctrl_serveStealReq_valid(_stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_37_ctrl_serveStealReq_ready(_stealNet_io_connSS_37_ctrl_serveStealReq_ready),
		.io_connSS_37_ctrl_stealReq_valid(_stealServers_36_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_37_ctrl_stealReq_ready(_stealNet_io_connSS_37_ctrl_stealReq_ready),
		.io_connSS_37_data_availableTask_ready(_stealServers_36_io_connNetwork_data_availableTask_ready),
		.io_connSS_37_data_availableTask_valid(_stealNet_io_connSS_37_data_availableTask_valid),
		.io_connSS_37_data_availableTask_bits(_stealNet_io_connSS_37_data_availableTask_bits),
		.io_connSS_37_data_qOutTask_ready(_stealNet_io_connSS_37_data_qOutTask_ready),
		.io_connSS_37_data_qOutTask_valid(_stealServers_36_io_connNetwork_data_qOutTask_valid),
		.io_connSS_37_data_qOutTask_bits(_stealServers_36_io_connNetwork_data_qOutTask_bits),
		.io_connSS_38_ctrl_serveStealReq_valid(_stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_38_ctrl_serveStealReq_ready(_stealNet_io_connSS_38_ctrl_serveStealReq_ready),
		.io_connSS_38_ctrl_stealReq_valid(_stealServers_37_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_38_ctrl_stealReq_ready(_stealNet_io_connSS_38_ctrl_stealReq_ready),
		.io_connSS_38_data_availableTask_ready(_stealServers_37_io_connNetwork_data_availableTask_ready),
		.io_connSS_38_data_availableTask_valid(_stealNet_io_connSS_38_data_availableTask_valid),
		.io_connSS_38_data_availableTask_bits(_stealNet_io_connSS_38_data_availableTask_bits),
		.io_connSS_38_data_qOutTask_ready(_stealNet_io_connSS_38_data_qOutTask_ready),
		.io_connSS_38_data_qOutTask_valid(_stealServers_37_io_connNetwork_data_qOutTask_valid),
		.io_connSS_38_data_qOutTask_bits(_stealServers_37_io_connNetwork_data_qOutTask_bits),
		.io_connSS_39_ctrl_serveStealReq_valid(_stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_39_ctrl_serveStealReq_ready(_stealNet_io_connSS_39_ctrl_serveStealReq_ready),
		.io_connSS_39_ctrl_stealReq_valid(_stealServers_38_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_39_ctrl_stealReq_ready(_stealNet_io_connSS_39_ctrl_stealReq_ready),
		.io_connSS_39_data_availableTask_ready(_stealServers_38_io_connNetwork_data_availableTask_ready),
		.io_connSS_39_data_availableTask_valid(_stealNet_io_connSS_39_data_availableTask_valid),
		.io_connSS_39_data_availableTask_bits(_stealNet_io_connSS_39_data_availableTask_bits),
		.io_connSS_39_data_qOutTask_ready(_stealNet_io_connSS_39_data_qOutTask_ready),
		.io_connSS_39_data_qOutTask_valid(_stealServers_38_io_connNetwork_data_qOutTask_valid),
		.io_connSS_39_data_qOutTask_bits(_stealServers_38_io_connNetwork_data_qOutTask_bits),
		.io_connSS_40_ctrl_serveStealReq_valid(_stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_40_ctrl_serveStealReq_ready(_stealNet_io_connSS_40_ctrl_serveStealReq_ready),
		.io_connSS_40_ctrl_stealReq_valid(_stealServers_39_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_40_ctrl_stealReq_ready(_stealNet_io_connSS_40_ctrl_stealReq_ready),
		.io_connSS_40_data_availableTask_ready(_stealServers_39_io_connNetwork_data_availableTask_ready),
		.io_connSS_40_data_availableTask_valid(_stealNet_io_connSS_40_data_availableTask_valid),
		.io_connSS_40_data_availableTask_bits(_stealNet_io_connSS_40_data_availableTask_bits),
		.io_connSS_40_data_qOutTask_ready(_stealNet_io_connSS_40_data_qOutTask_ready),
		.io_connSS_40_data_qOutTask_valid(_stealServers_39_io_connNetwork_data_qOutTask_valid),
		.io_connSS_40_data_qOutTask_bits(_stealServers_39_io_connNetwork_data_qOutTask_bits),
		.io_connSS_41_ctrl_serveStealReq_valid(_stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_41_ctrl_serveStealReq_ready(_stealNet_io_connSS_41_ctrl_serveStealReq_ready),
		.io_connSS_41_ctrl_stealReq_valid(_stealServers_40_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_41_ctrl_stealReq_ready(_stealNet_io_connSS_41_ctrl_stealReq_ready),
		.io_connSS_41_data_availableTask_ready(_stealServers_40_io_connNetwork_data_availableTask_ready),
		.io_connSS_41_data_availableTask_valid(_stealNet_io_connSS_41_data_availableTask_valid),
		.io_connSS_41_data_availableTask_bits(_stealNet_io_connSS_41_data_availableTask_bits),
		.io_connSS_41_data_qOutTask_ready(_stealNet_io_connSS_41_data_qOutTask_ready),
		.io_connSS_41_data_qOutTask_valid(_stealServers_40_io_connNetwork_data_qOutTask_valid),
		.io_connSS_41_data_qOutTask_bits(_stealServers_40_io_connNetwork_data_qOutTask_bits),
		.io_connSS_42_ctrl_serveStealReq_valid(_stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_42_ctrl_serveStealReq_ready(_stealNet_io_connSS_42_ctrl_serveStealReq_ready),
		.io_connSS_42_ctrl_stealReq_valid(_stealServers_41_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_42_ctrl_stealReq_ready(_stealNet_io_connSS_42_ctrl_stealReq_ready),
		.io_connSS_42_data_availableTask_ready(_stealServers_41_io_connNetwork_data_availableTask_ready),
		.io_connSS_42_data_availableTask_valid(_stealNet_io_connSS_42_data_availableTask_valid),
		.io_connSS_42_data_availableTask_bits(_stealNet_io_connSS_42_data_availableTask_bits),
		.io_connSS_42_data_qOutTask_ready(_stealNet_io_connSS_42_data_qOutTask_ready),
		.io_connSS_42_data_qOutTask_valid(_stealServers_41_io_connNetwork_data_qOutTask_valid),
		.io_connSS_42_data_qOutTask_bits(_stealServers_41_io_connNetwork_data_qOutTask_bits),
		.io_connSS_43_ctrl_serveStealReq_valid(_stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_43_ctrl_serveStealReq_ready(_stealNet_io_connSS_43_ctrl_serveStealReq_ready),
		.io_connSS_43_ctrl_stealReq_valid(_stealServers_42_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_43_ctrl_stealReq_ready(_stealNet_io_connSS_43_ctrl_stealReq_ready),
		.io_connSS_43_data_availableTask_ready(_stealServers_42_io_connNetwork_data_availableTask_ready),
		.io_connSS_43_data_availableTask_valid(_stealNet_io_connSS_43_data_availableTask_valid),
		.io_connSS_43_data_availableTask_bits(_stealNet_io_connSS_43_data_availableTask_bits),
		.io_connSS_43_data_qOutTask_ready(_stealNet_io_connSS_43_data_qOutTask_ready),
		.io_connSS_43_data_qOutTask_valid(_stealServers_42_io_connNetwork_data_qOutTask_valid),
		.io_connSS_43_data_qOutTask_bits(_stealServers_42_io_connNetwork_data_qOutTask_bits),
		.io_connSS_44_ctrl_serveStealReq_valid(_stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_44_ctrl_serveStealReq_ready(_stealNet_io_connSS_44_ctrl_serveStealReq_ready),
		.io_connSS_44_ctrl_stealReq_valid(_stealServers_43_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_44_ctrl_stealReq_ready(_stealNet_io_connSS_44_ctrl_stealReq_ready),
		.io_connSS_44_data_availableTask_ready(_stealServers_43_io_connNetwork_data_availableTask_ready),
		.io_connSS_44_data_availableTask_valid(_stealNet_io_connSS_44_data_availableTask_valid),
		.io_connSS_44_data_availableTask_bits(_stealNet_io_connSS_44_data_availableTask_bits),
		.io_connSS_44_data_qOutTask_ready(_stealNet_io_connSS_44_data_qOutTask_ready),
		.io_connSS_44_data_qOutTask_valid(_stealServers_43_io_connNetwork_data_qOutTask_valid),
		.io_connSS_44_data_qOutTask_bits(_stealServers_43_io_connNetwork_data_qOutTask_bits),
		.io_connSS_45_ctrl_serveStealReq_valid(_stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_45_ctrl_serveStealReq_ready(_stealNet_io_connSS_45_ctrl_serveStealReq_ready),
		.io_connSS_45_ctrl_stealReq_valid(_stealServers_44_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_45_ctrl_stealReq_ready(_stealNet_io_connSS_45_ctrl_stealReq_ready),
		.io_connSS_45_data_availableTask_ready(_stealServers_44_io_connNetwork_data_availableTask_ready),
		.io_connSS_45_data_availableTask_valid(_stealNet_io_connSS_45_data_availableTask_valid),
		.io_connSS_45_data_availableTask_bits(_stealNet_io_connSS_45_data_availableTask_bits),
		.io_connSS_45_data_qOutTask_ready(_stealNet_io_connSS_45_data_qOutTask_ready),
		.io_connSS_45_data_qOutTask_valid(_stealServers_44_io_connNetwork_data_qOutTask_valid),
		.io_connSS_45_data_qOutTask_bits(_stealServers_44_io_connNetwork_data_qOutTask_bits),
		.io_connSS_46_ctrl_serveStealReq_valid(_stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_46_ctrl_serveStealReq_ready(_stealNet_io_connSS_46_ctrl_serveStealReq_ready),
		.io_connSS_46_ctrl_stealReq_valid(_stealServers_45_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_46_ctrl_stealReq_ready(_stealNet_io_connSS_46_ctrl_stealReq_ready),
		.io_connSS_46_data_availableTask_ready(_stealServers_45_io_connNetwork_data_availableTask_ready),
		.io_connSS_46_data_availableTask_valid(_stealNet_io_connSS_46_data_availableTask_valid),
		.io_connSS_46_data_availableTask_bits(_stealNet_io_connSS_46_data_availableTask_bits),
		.io_connSS_46_data_qOutTask_ready(_stealNet_io_connSS_46_data_qOutTask_ready),
		.io_connSS_46_data_qOutTask_valid(_stealServers_45_io_connNetwork_data_qOutTask_valid),
		.io_connSS_46_data_qOutTask_bits(_stealServers_45_io_connNetwork_data_qOutTask_bits),
		.io_connSS_47_ctrl_serveStealReq_valid(_stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_47_ctrl_serveStealReq_ready(_stealNet_io_connSS_47_ctrl_serveStealReq_ready),
		.io_connSS_47_ctrl_stealReq_valid(_stealServers_46_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_47_ctrl_stealReq_ready(_stealNet_io_connSS_47_ctrl_stealReq_ready),
		.io_connSS_47_data_availableTask_ready(_stealServers_46_io_connNetwork_data_availableTask_ready),
		.io_connSS_47_data_availableTask_valid(_stealNet_io_connSS_47_data_availableTask_valid),
		.io_connSS_47_data_availableTask_bits(_stealNet_io_connSS_47_data_availableTask_bits),
		.io_connSS_47_data_qOutTask_ready(_stealNet_io_connSS_47_data_qOutTask_ready),
		.io_connSS_47_data_qOutTask_valid(_stealServers_46_io_connNetwork_data_qOutTask_valid),
		.io_connSS_47_data_qOutTask_bits(_stealServers_46_io_connNetwork_data_qOutTask_bits),
		.io_connSS_48_ctrl_serveStealReq_valid(_stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_48_ctrl_serveStealReq_ready(_stealNet_io_connSS_48_ctrl_serveStealReq_ready),
		.io_connSS_48_ctrl_stealReq_valid(_stealServers_47_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_48_ctrl_stealReq_ready(_stealNet_io_connSS_48_ctrl_stealReq_ready),
		.io_connSS_48_data_availableTask_ready(_stealServers_47_io_connNetwork_data_availableTask_ready),
		.io_connSS_48_data_availableTask_valid(_stealNet_io_connSS_48_data_availableTask_valid),
		.io_connSS_48_data_availableTask_bits(_stealNet_io_connSS_48_data_availableTask_bits),
		.io_connSS_48_data_qOutTask_ready(_stealNet_io_connSS_48_data_qOutTask_ready),
		.io_connSS_48_data_qOutTask_valid(_stealServers_47_io_connNetwork_data_qOutTask_valid),
		.io_connSS_48_data_qOutTask_bits(_stealServers_47_io_connNetwork_data_qOutTask_bits),
		.io_connSS_49_ctrl_serveStealReq_valid(_stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_49_ctrl_serveStealReq_ready(_stealNet_io_connSS_49_ctrl_serveStealReq_ready),
		.io_connSS_49_ctrl_stealReq_valid(_stealServers_48_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_49_ctrl_stealReq_ready(_stealNet_io_connSS_49_ctrl_stealReq_ready),
		.io_connSS_49_data_availableTask_ready(_stealServers_48_io_connNetwork_data_availableTask_ready),
		.io_connSS_49_data_availableTask_valid(_stealNet_io_connSS_49_data_availableTask_valid),
		.io_connSS_49_data_availableTask_bits(_stealNet_io_connSS_49_data_availableTask_bits),
		.io_connSS_49_data_qOutTask_ready(_stealNet_io_connSS_49_data_qOutTask_ready),
		.io_connSS_49_data_qOutTask_valid(_stealServers_48_io_connNetwork_data_qOutTask_valid),
		.io_connSS_49_data_qOutTask_bits(_stealServers_48_io_connNetwork_data_qOutTask_bits),
		.io_connSS_50_ctrl_serveStealReq_valid(_stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_50_ctrl_serveStealReq_ready(_stealNet_io_connSS_50_ctrl_serveStealReq_ready),
		.io_connSS_50_ctrl_stealReq_valid(_stealServers_49_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_50_ctrl_stealReq_ready(_stealNet_io_connSS_50_ctrl_stealReq_ready),
		.io_connSS_50_data_availableTask_ready(_stealServers_49_io_connNetwork_data_availableTask_ready),
		.io_connSS_50_data_availableTask_valid(_stealNet_io_connSS_50_data_availableTask_valid),
		.io_connSS_50_data_availableTask_bits(_stealNet_io_connSS_50_data_availableTask_bits),
		.io_connSS_50_data_qOutTask_ready(_stealNet_io_connSS_50_data_qOutTask_ready),
		.io_connSS_50_data_qOutTask_valid(_stealServers_49_io_connNetwork_data_qOutTask_valid),
		.io_connSS_50_data_qOutTask_bits(_stealServers_49_io_connNetwork_data_qOutTask_bits),
		.io_connSS_51_ctrl_serveStealReq_valid(_stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_51_ctrl_serveStealReq_ready(_stealNet_io_connSS_51_ctrl_serveStealReq_ready),
		.io_connSS_51_ctrl_stealReq_valid(_stealServers_50_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_51_ctrl_stealReq_ready(_stealNet_io_connSS_51_ctrl_stealReq_ready),
		.io_connSS_51_data_availableTask_ready(_stealServers_50_io_connNetwork_data_availableTask_ready),
		.io_connSS_51_data_availableTask_valid(_stealNet_io_connSS_51_data_availableTask_valid),
		.io_connSS_51_data_availableTask_bits(_stealNet_io_connSS_51_data_availableTask_bits),
		.io_connSS_51_data_qOutTask_ready(_stealNet_io_connSS_51_data_qOutTask_ready),
		.io_connSS_51_data_qOutTask_valid(_stealServers_50_io_connNetwork_data_qOutTask_valid),
		.io_connSS_51_data_qOutTask_bits(_stealServers_50_io_connNetwork_data_qOutTask_bits),
		.io_connSS_52_ctrl_serveStealReq_valid(_stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_52_ctrl_serveStealReq_ready(_stealNet_io_connSS_52_ctrl_serveStealReq_ready),
		.io_connSS_52_ctrl_stealReq_valid(_stealServers_51_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_52_ctrl_stealReq_ready(_stealNet_io_connSS_52_ctrl_stealReq_ready),
		.io_connSS_52_data_availableTask_ready(_stealServers_51_io_connNetwork_data_availableTask_ready),
		.io_connSS_52_data_availableTask_valid(_stealNet_io_connSS_52_data_availableTask_valid),
		.io_connSS_52_data_availableTask_bits(_stealNet_io_connSS_52_data_availableTask_bits),
		.io_connSS_52_data_qOutTask_ready(_stealNet_io_connSS_52_data_qOutTask_ready),
		.io_connSS_52_data_qOutTask_valid(_stealServers_51_io_connNetwork_data_qOutTask_valid),
		.io_connSS_52_data_qOutTask_bits(_stealServers_51_io_connNetwork_data_qOutTask_bits),
		.io_connSS_53_ctrl_serveStealReq_valid(_stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_53_ctrl_serveStealReq_ready(_stealNet_io_connSS_53_ctrl_serveStealReq_ready),
		.io_connSS_53_ctrl_stealReq_valid(_stealServers_52_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_53_ctrl_stealReq_ready(_stealNet_io_connSS_53_ctrl_stealReq_ready),
		.io_connSS_53_data_availableTask_ready(_stealServers_52_io_connNetwork_data_availableTask_ready),
		.io_connSS_53_data_availableTask_valid(_stealNet_io_connSS_53_data_availableTask_valid),
		.io_connSS_53_data_availableTask_bits(_stealNet_io_connSS_53_data_availableTask_bits),
		.io_connSS_53_data_qOutTask_ready(_stealNet_io_connSS_53_data_qOutTask_ready),
		.io_connSS_53_data_qOutTask_valid(_stealServers_52_io_connNetwork_data_qOutTask_valid),
		.io_connSS_53_data_qOutTask_bits(_stealServers_52_io_connNetwork_data_qOutTask_bits),
		.io_connSS_54_ctrl_serveStealReq_valid(_stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_54_ctrl_serveStealReq_ready(_stealNet_io_connSS_54_ctrl_serveStealReq_ready),
		.io_connSS_54_ctrl_stealReq_valid(_stealServers_53_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_54_ctrl_stealReq_ready(_stealNet_io_connSS_54_ctrl_stealReq_ready),
		.io_connSS_54_data_availableTask_ready(_stealServers_53_io_connNetwork_data_availableTask_ready),
		.io_connSS_54_data_availableTask_valid(_stealNet_io_connSS_54_data_availableTask_valid),
		.io_connSS_54_data_availableTask_bits(_stealNet_io_connSS_54_data_availableTask_bits),
		.io_connSS_54_data_qOutTask_ready(_stealNet_io_connSS_54_data_qOutTask_ready),
		.io_connSS_54_data_qOutTask_valid(_stealServers_53_io_connNetwork_data_qOutTask_valid),
		.io_connSS_54_data_qOutTask_bits(_stealServers_53_io_connNetwork_data_qOutTask_bits),
		.io_connSS_55_ctrl_serveStealReq_valid(_stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_55_ctrl_serveStealReq_ready(_stealNet_io_connSS_55_ctrl_serveStealReq_ready),
		.io_connSS_55_ctrl_stealReq_valid(_stealServers_54_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_55_ctrl_stealReq_ready(_stealNet_io_connSS_55_ctrl_stealReq_ready),
		.io_connSS_55_data_availableTask_ready(_stealServers_54_io_connNetwork_data_availableTask_ready),
		.io_connSS_55_data_availableTask_valid(_stealNet_io_connSS_55_data_availableTask_valid),
		.io_connSS_55_data_availableTask_bits(_stealNet_io_connSS_55_data_availableTask_bits),
		.io_connSS_55_data_qOutTask_ready(_stealNet_io_connSS_55_data_qOutTask_ready),
		.io_connSS_55_data_qOutTask_valid(_stealServers_54_io_connNetwork_data_qOutTask_valid),
		.io_connSS_55_data_qOutTask_bits(_stealServers_54_io_connNetwork_data_qOutTask_bits),
		.io_connSS_56_ctrl_serveStealReq_valid(_stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_56_ctrl_serveStealReq_ready(_stealNet_io_connSS_56_ctrl_serveStealReq_ready),
		.io_connSS_56_ctrl_stealReq_valid(_stealServers_55_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_56_ctrl_stealReq_ready(_stealNet_io_connSS_56_ctrl_stealReq_ready),
		.io_connSS_56_data_availableTask_ready(_stealServers_55_io_connNetwork_data_availableTask_ready),
		.io_connSS_56_data_availableTask_valid(_stealNet_io_connSS_56_data_availableTask_valid),
		.io_connSS_56_data_availableTask_bits(_stealNet_io_connSS_56_data_availableTask_bits),
		.io_connSS_56_data_qOutTask_ready(_stealNet_io_connSS_56_data_qOutTask_ready),
		.io_connSS_56_data_qOutTask_valid(_stealServers_55_io_connNetwork_data_qOutTask_valid),
		.io_connSS_56_data_qOutTask_bits(_stealServers_55_io_connNetwork_data_qOutTask_bits),
		.io_connSS_57_ctrl_serveStealReq_valid(_stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_57_ctrl_serveStealReq_ready(_stealNet_io_connSS_57_ctrl_serveStealReq_ready),
		.io_connSS_57_ctrl_stealReq_valid(_stealServers_56_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_57_ctrl_stealReq_ready(_stealNet_io_connSS_57_ctrl_stealReq_ready),
		.io_connSS_57_data_availableTask_ready(_stealServers_56_io_connNetwork_data_availableTask_ready),
		.io_connSS_57_data_availableTask_valid(_stealNet_io_connSS_57_data_availableTask_valid),
		.io_connSS_57_data_availableTask_bits(_stealNet_io_connSS_57_data_availableTask_bits),
		.io_connSS_57_data_qOutTask_ready(_stealNet_io_connSS_57_data_qOutTask_ready),
		.io_connSS_57_data_qOutTask_valid(_stealServers_56_io_connNetwork_data_qOutTask_valid),
		.io_connSS_57_data_qOutTask_bits(_stealServers_56_io_connNetwork_data_qOutTask_bits),
		.io_connSS_58_ctrl_serveStealReq_valid(_stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_58_ctrl_serveStealReq_ready(_stealNet_io_connSS_58_ctrl_serveStealReq_ready),
		.io_connSS_58_ctrl_stealReq_valid(_stealServers_57_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_58_ctrl_stealReq_ready(_stealNet_io_connSS_58_ctrl_stealReq_ready),
		.io_connSS_58_data_availableTask_ready(_stealServers_57_io_connNetwork_data_availableTask_ready),
		.io_connSS_58_data_availableTask_valid(_stealNet_io_connSS_58_data_availableTask_valid),
		.io_connSS_58_data_availableTask_bits(_stealNet_io_connSS_58_data_availableTask_bits),
		.io_connSS_58_data_qOutTask_ready(_stealNet_io_connSS_58_data_qOutTask_ready),
		.io_connSS_58_data_qOutTask_valid(_stealServers_57_io_connNetwork_data_qOutTask_valid),
		.io_connSS_58_data_qOutTask_bits(_stealServers_57_io_connNetwork_data_qOutTask_bits),
		.io_connSS_59_ctrl_serveStealReq_valid(_stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_59_ctrl_serveStealReq_ready(_stealNet_io_connSS_59_ctrl_serveStealReq_ready),
		.io_connSS_59_ctrl_stealReq_valid(_stealServers_58_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_59_ctrl_stealReq_ready(_stealNet_io_connSS_59_ctrl_stealReq_ready),
		.io_connSS_59_data_availableTask_ready(_stealServers_58_io_connNetwork_data_availableTask_ready),
		.io_connSS_59_data_availableTask_valid(_stealNet_io_connSS_59_data_availableTask_valid),
		.io_connSS_59_data_availableTask_bits(_stealNet_io_connSS_59_data_availableTask_bits),
		.io_connSS_59_data_qOutTask_ready(_stealNet_io_connSS_59_data_qOutTask_ready),
		.io_connSS_59_data_qOutTask_valid(_stealServers_58_io_connNetwork_data_qOutTask_valid),
		.io_connSS_59_data_qOutTask_bits(_stealServers_58_io_connNetwork_data_qOutTask_bits),
		.io_connSS_60_ctrl_serveStealReq_valid(_stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_60_ctrl_serveStealReq_ready(_stealNet_io_connSS_60_ctrl_serveStealReq_ready),
		.io_connSS_60_ctrl_stealReq_valid(_stealServers_59_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_60_ctrl_stealReq_ready(_stealNet_io_connSS_60_ctrl_stealReq_ready),
		.io_connSS_60_data_availableTask_ready(_stealServers_59_io_connNetwork_data_availableTask_ready),
		.io_connSS_60_data_availableTask_valid(_stealNet_io_connSS_60_data_availableTask_valid),
		.io_connSS_60_data_availableTask_bits(_stealNet_io_connSS_60_data_availableTask_bits),
		.io_connSS_60_data_qOutTask_ready(_stealNet_io_connSS_60_data_qOutTask_ready),
		.io_connSS_60_data_qOutTask_valid(_stealServers_59_io_connNetwork_data_qOutTask_valid),
		.io_connSS_60_data_qOutTask_bits(_stealServers_59_io_connNetwork_data_qOutTask_bits),
		.io_connSS_61_ctrl_serveStealReq_valid(_stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_61_ctrl_serveStealReq_ready(_stealNet_io_connSS_61_ctrl_serveStealReq_ready),
		.io_connSS_61_ctrl_stealReq_valid(_stealServers_60_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_61_ctrl_stealReq_ready(_stealNet_io_connSS_61_ctrl_stealReq_ready),
		.io_connSS_61_data_availableTask_ready(_stealServers_60_io_connNetwork_data_availableTask_ready),
		.io_connSS_61_data_availableTask_valid(_stealNet_io_connSS_61_data_availableTask_valid),
		.io_connSS_61_data_availableTask_bits(_stealNet_io_connSS_61_data_availableTask_bits),
		.io_connSS_61_data_qOutTask_ready(_stealNet_io_connSS_61_data_qOutTask_ready),
		.io_connSS_61_data_qOutTask_valid(_stealServers_60_io_connNetwork_data_qOutTask_valid),
		.io_connSS_61_data_qOutTask_bits(_stealServers_60_io_connNetwork_data_qOutTask_bits),
		.io_connSS_62_ctrl_serveStealReq_valid(_stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_62_ctrl_serveStealReq_ready(_stealNet_io_connSS_62_ctrl_serveStealReq_ready),
		.io_connSS_62_ctrl_stealReq_valid(_stealServers_61_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_62_ctrl_stealReq_ready(_stealNet_io_connSS_62_ctrl_stealReq_ready),
		.io_connSS_62_data_availableTask_ready(_stealServers_61_io_connNetwork_data_availableTask_ready),
		.io_connSS_62_data_availableTask_valid(_stealNet_io_connSS_62_data_availableTask_valid),
		.io_connSS_62_data_availableTask_bits(_stealNet_io_connSS_62_data_availableTask_bits),
		.io_connSS_62_data_qOutTask_ready(_stealNet_io_connSS_62_data_qOutTask_ready),
		.io_connSS_62_data_qOutTask_valid(_stealServers_61_io_connNetwork_data_qOutTask_valid),
		.io_connSS_62_data_qOutTask_bits(_stealServers_61_io_connNetwork_data_qOutTask_bits),
		.io_connSS_63_ctrl_serveStealReq_valid(_stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_63_ctrl_serveStealReq_ready(_stealNet_io_connSS_63_ctrl_serveStealReq_ready),
		.io_connSS_63_ctrl_stealReq_valid(_stealServers_62_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_63_ctrl_stealReq_ready(_stealNet_io_connSS_63_ctrl_stealReq_ready),
		.io_connSS_63_data_availableTask_ready(_stealServers_62_io_connNetwork_data_availableTask_ready),
		.io_connSS_63_data_availableTask_valid(_stealNet_io_connSS_63_data_availableTask_valid),
		.io_connSS_63_data_availableTask_bits(_stealNet_io_connSS_63_data_availableTask_bits),
		.io_connSS_63_data_qOutTask_ready(_stealNet_io_connSS_63_data_qOutTask_ready),
		.io_connSS_63_data_qOutTask_valid(_stealServers_62_io_connNetwork_data_qOutTask_valid),
		.io_connSS_63_data_qOutTask_bits(_stealServers_62_io_connNetwork_data_qOutTask_bits),
		.io_connSS_64_ctrl_serveStealReq_valid(_stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_64_ctrl_serveStealReq_ready(_stealNet_io_connSS_64_ctrl_serveStealReq_ready),
		.io_connSS_64_ctrl_stealReq_valid(_stealServers_63_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_64_ctrl_stealReq_ready(_stealNet_io_connSS_64_ctrl_stealReq_ready),
		.io_connSS_64_data_availableTask_ready(_stealServers_63_io_connNetwork_data_availableTask_ready),
		.io_connSS_64_data_availableTask_valid(_stealNet_io_connSS_64_data_availableTask_valid),
		.io_connSS_64_data_availableTask_bits(_stealNet_io_connSS_64_data_availableTask_bits),
		.io_connSS_64_data_qOutTask_ready(_stealNet_io_connSS_64_data_qOutTask_ready),
		.io_connSS_64_data_qOutTask_valid(_stealServers_63_io_connNetwork_data_qOutTask_valid),
		.io_connSS_64_data_qOutTask_bits(_stealServers_63_io_connNetwork_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerClient stealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_1_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_1_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_1_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_1_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_1_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_0_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_2_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_2_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_2_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_2_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_2_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_1_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_2(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_3_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_3_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_3_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_3_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_3_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_2_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_3(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_4_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_4_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_4_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_4_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_4_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_3_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_4(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_5_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_5_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_5_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_5_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_5_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_4_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_5(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_6_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_6_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_6_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_6_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_6_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_5_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_6(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_7_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_7_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_7_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_7_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_7_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_6_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_7(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_8_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_8_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_8_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_8_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_8_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_7_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_8(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_9_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_9_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_9_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_9_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_9_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_8_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_9(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_10_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_10_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_10_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_10_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_10_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_9_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_10(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_11_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_11_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_11_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_11_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_11_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_10_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_11(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_12_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_12_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_12_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_12_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_12_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_11_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_12(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_13_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_13_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_13_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_13_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_13_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_12_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_13(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_14_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_14_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_14_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_14_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_14_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_13_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_14(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_15_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_15_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_15_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_15_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_15_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_14_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_15(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_16_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_16_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_16_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_16_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_16_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_15_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_16(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_16_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_17_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_16_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_17_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_16_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_17_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_17_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_17_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_16_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_16_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_16_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_16_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_16_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_16_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_16_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_16_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_16_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_17(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_17_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_17_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_17_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_17_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_17_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_17_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_17_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_17_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_17_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_17_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_17_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_17_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_18(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_18_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_18_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_18_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_18_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_18_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_18_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_18_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_18_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_18_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_18_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_18_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_18_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_19(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_19_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_19_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_19_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_19_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_19_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_19_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_19_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_19_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_19_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_19_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_19_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_19_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_20(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_20_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_20_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_20_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_20_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_20_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_20_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_20_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_20_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_20_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_20_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_20_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_20_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_21(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_21_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_21_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_21_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_21_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_21_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_21_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_21_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_21_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_21_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_21_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_21_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_21_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_22(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_22_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_22_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_22_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_22_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_22_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_22_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_22_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_22_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_22_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_22_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_22_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_22_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_23(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_23_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_23_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_23_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_23_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_23_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_23_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_23_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_23_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_23_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_23_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_23_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_23_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_24(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_24_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_24_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_24_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_24_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_24_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_24_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_24_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_24_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_24_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_24_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_24_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_24_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_25(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_25_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_25_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_25_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_25_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_25_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_25_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_25_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_25_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_25_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_25_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_25_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_25_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_26(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_26_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_26_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_26_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_26_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_26_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_26_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_26_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_26_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_26_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_26_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_26_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_26_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_27(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_27_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_27_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_27_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_27_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_27_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_27_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_27_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_27_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_27_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_27_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_27_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_27_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_28(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_28_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_28_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_28_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_28_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_28_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_28_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_28_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_28_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_28_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_28_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_28_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_28_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_29(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_29_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_29_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_29_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_29_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_29_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_29_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_29_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_29_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_29_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_29_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_29_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_29_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_30(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_30_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_30_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_30_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_30_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_30_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_30_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_30_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_30_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_30_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_30_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_30_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_30_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_31(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_31_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_31_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_31_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_31_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_31_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_31_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_31_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_31_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_31_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_31_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_31_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_31_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_32(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_32_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_33_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_32_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_33_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_32_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_33_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_33_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_33_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_32_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_32_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_32_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_32_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_32_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_32_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_32_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_32_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_32_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_33(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_33_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_34_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_33_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_34_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_33_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_34_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_34_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_34_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_33_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_33_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_33_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_33_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_33_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_33_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_33_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_33_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_33_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_34(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_34_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_35_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_34_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_35_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_34_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_35_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_35_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_35_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_34_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_34_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_34_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_34_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_34_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_34_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_34_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_34_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_34_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_35(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_35_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_36_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_35_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_36_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_35_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_36_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_36_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_36_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_35_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_35_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_35_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_35_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_35_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_35_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_35_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_35_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_35_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_36(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_36_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_37_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_36_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_37_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_36_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_37_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_37_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_37_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_36_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_36_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_36_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_36_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_36_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_36_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_36_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_36_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_36_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_37(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_37_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_38_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_37_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_38_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_37_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_38_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_38_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_38_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_37_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_37_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_37_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_37_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_37_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_37_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_37_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_37_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_37_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_38(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_38_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_39_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_38_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_39_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_38_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_39_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_39_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_39_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_38_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_38_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_38_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_38_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_38_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_38_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_38_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_38_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_38_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_39(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_39_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_40_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_39_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_40_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_39_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_40_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_40_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_40_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_39_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_39_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_39_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_39_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_39_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_39_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_39_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_39_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_39_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_40(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_40_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_41_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_40_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_41_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_40_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_41_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_41_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_41_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_40_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_40_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_40_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_40_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_40_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_40_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_40_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_40_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_40_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_41(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_41_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_42_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_41_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_42_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_41_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_42_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_42_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_42_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_41_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_41_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_41_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_41_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_41_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_41_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_41_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_41_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_41_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_42(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_42_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_43_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_42_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_43_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_42_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_43_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_43_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_43_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_42_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_42_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_42_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_42_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_42_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_42_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_42_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_42_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_42_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_43(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_43_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_44_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_43_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_44_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_43_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_44_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_44_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_44_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_43_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_43_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_43_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_43_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_43_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_43_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_43_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_43_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_43_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_44(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_44_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_45_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_44_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_45_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_44_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_45_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_45_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_45_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_44_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_44_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_44_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_44_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_44_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_44_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_44_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_44_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_44_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_45(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_45_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_46_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_45_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_46_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_45_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_46_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_46_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_46_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_45_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_45_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_45_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_45_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_45_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_45_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_45_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_45_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_45_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_46(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_46_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_47_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_46_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_47_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_46_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_47_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_47_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_47_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_46_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_46_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_46_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_46_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_46_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_46_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_46_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_46_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_46_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_47(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_47_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_48_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_47_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_48_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_47_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_48_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_48_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_48_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_47_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_47_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_47_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_47_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_47_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_47_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_47_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_47_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_47_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_48(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_48_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_49_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_48_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_49_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_48_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_49_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_49_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_49_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_48_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_48_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_48_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_48_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_48_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_48_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_48_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_48_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_48_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_49(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_49_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_50_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_49_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_50_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_49_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_50_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_50_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_50_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_49_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_49_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_49_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_49_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_49_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_49_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_49_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_49_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_49_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_50(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_50_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_51_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_50_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_51_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_50_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_51_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_51_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_51_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_50_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_50_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_50_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_50_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_50_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_50_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_50_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_50_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_50_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_51(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_51_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_52_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_51_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_52_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_51_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_52_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_52_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_52_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_51_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_51_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_51_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_51_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_51_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_51_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_51_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_51_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_51_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_52(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_52_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_53_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_52_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_53_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_52_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_53_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_53_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_53_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_52_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_52_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_52_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_52_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_52_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_52_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_52_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_52_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_52_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_53(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_53_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_54_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_53_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_54_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_53_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_54_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_54_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_54_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_53_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_53_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_53_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_53_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_53_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_53_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_53_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_53_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_53_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_54(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_54_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_55_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_54_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_55_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_54_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_55_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_55_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_55_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_54_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_54_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_54_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_54_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_54_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_54_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_54_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_54_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_54_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_55(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_55_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_56_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_55_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_56_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_55_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_56_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_56_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_56_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_55_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_55_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_55_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_55_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_55_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_55_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_55_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_55_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_55_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_56(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_56_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_57_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_56_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_57_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_56_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_57_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_57_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_57_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_56_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_56_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_56_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_56_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_56_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_56_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_56_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_56_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_56_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_57(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_57_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_58_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_57_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_58_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_57_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_58_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_58_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_58_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_57_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_57_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_57_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_57_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_57_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_57_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_57_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_57_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_57_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_58(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_58_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_59_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_58_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_59_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_58_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_59_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_59_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_59_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_58_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_58_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_58_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_58_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_58_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_58_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_58_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_58_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_58_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_59(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_59_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_60_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_59_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_60_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_59_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_60_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_60_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_60_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_59_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_59_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_59_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_59_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_59_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_59_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_59_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_59_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_59_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_60(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_60_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_61_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_60_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_61_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_60_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_61_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_61_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_61_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_60_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_60_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_60_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_60_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_60_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_60_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_60_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_60_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_60_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_61(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_61_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_62_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_61_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_62_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_61_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_62_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_62_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_62_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_61_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_61_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_61_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_61_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_61_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_61_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_61_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_61_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_61_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_62(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_62_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_63_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_62_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_63_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_62_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_63_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_63_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_63_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_62_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_62_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_62_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_62_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_62_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_62_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_62_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_62_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_62_io_connVec_1_pop_bits)
	);
	SchedulerClient stealServers_63(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_63_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_64_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_63_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_64_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_63_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_64_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_64_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_64_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_63_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_63_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_63_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_63_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_63_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_63_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_63_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_63_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_63_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_0(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_0_push_ready),
		.io_connVec_0_push_valid(io_connPE_0_push_valid),
		.io_connVec_0_push_bits(io_connPE_0_push_bits),
		.io_connVec_0_pop_ready(io_connPE_0_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_0_pop_valid),
		.io_connVec_1_currLength(_taskQueues_0_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_1(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_1_push_ready),
		.io_connVec_0_push_valid(io_connPE_1_push_valid),
		.io_connVec_0_push_bits(io_connPE_1_push_bits),
		.io_connVec_0_pop_ready(io_connPE_1_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_1_pop_valid),
		.io_connVec_1_currLength(_taskQueues_1_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_2(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_2_push_ready),
		.io_connVec_0_push_valid(io_connPE_2_push_valid),
		.io_connVec_0_push_bits(io_connPE_2_push_bits),
		.io_connVec_0_pop_ready(io_connPE_2_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_2_pop_valid),
		.io_connVec_1_currLength(_taskQueues_2_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_3(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_3_push_ready),
		.io_connVec_0_push_valid(io_connPE_3_push_valid),
		.io_connVec_0_push_bits(io_connPE_3_push_bits),
		.io_connVec_0_pop_ready(io_connPE_3_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_3_pop_valid),
		.io_connVec_1_currLength(_taskQueues_3_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_4(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_4_push_ready),
		.io_connVec_0_push_valid(io_connPE_4_push_valid),
		.io_connVec_0_push_bits(io_connPE_4_push_bits),
		.io_connVec_0_pop_ready(io_connPE_4_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_4_pop_valid),
		.io_connVec_1_currLength(_taskQueues_4_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_5(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_5_push_ready),
		.io_connVec_0_push_valid(io_connPE_5_push_valid),
		.io_connVec_0_push_bits(io_connPE_5_push_bits),
		.io_connVec_0_pop_ready(io_connPE_5_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_5_pop_valid),
		.io_connVec_1_currLength(_taskQueues_5_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_6(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_6_push_ready),
		.io_connVec_0_push_valid(io_connPE_6_push_valid),
		.io_connVec_0_push_bits(io_connPE_6_push_bits),
		.io_connVec_0_pop_ready(io_connPE_6_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_6_pop_valid),
		.io_connVec_1_currLength(_taskQueues_6_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_7(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_7_push_ready),
		.io_connVec_0_push_valid(io_connPE_7_push_valid),
		.io_connVec_0_push_bits(io_connPE_7_push_bits),
		.io_connVec_0_pop_ready(io_connPE_7_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_7_pop_valid),
		.io_connVec_1_currLength(_taskQueues_7_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_8(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_8_push_ready),
		.io_connVec_0_push_valid(io_connPE_8_push_valid),
		.io_connVec_0_push_bits(io_connPE_8_push_bits),
		.io_connVec_0_pop_ready(io_connPE_8_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_8_pop_valid),
		.io_connVec_1_currLength(_taskQueues_8_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_9(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_9_push_ready),
		.io_connVec_0_push_valid(io_connPE_9_push_valid),
		.io_connVec_0_push_bits(io_connPE_9_push_bits),
		.io_connVec_0_pop_ready(io_connPE_9_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_9_pop_valid),
		.io_connVec_1_currLength(_taskQueues_9_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_10(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_10_push_ready),
		.io_connVec_0_push_valid(io_connPE_10_push_valid),
		.io_connVec_0_push_bits(io_connPE_10_push_bits),
		.io_connVec_0_pop_ready(io_connPE_10_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_10_pop_valid),
		.io_connVec_1_currLength(_taskQueues_10_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_11(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_11_push_ready),
		.io_connVec_0_push_valid(io_connPE_11_push_valid),
		.io_connVec_0_push_bits(io_connPE_11_push_bits),
		.io_connVec_0_pop_ready(io_connPE_11_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_11_pop_valid),
		.io_connVec_1_currLength(_taskQueues_11_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_12(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_12_push_ready),
		.io_connVec_0_push_valid(io_connPE_12_push_valid),
		.io_connVec_0_push_bits(io_connPE_12_push_bits),
		.io_connVec_0_pop_ready(io_connPE_12_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_12_pop_valid),
		.io_connVec_1_currLength(_taskQueues_12_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_13(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_13_push_ready),
		.io_connVec_0_push_valid(io_connPE_13_push_valid),
		.io_connVec_0_push_bits(io_connPE_13_push_bits),
		.io_connVec_0_pop_ready(io_connPE_13_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_13_pop_valid),
		.io_connVec_1_currLength(_taskQueues_13_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_14(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_14_push_ready),
		.io_connVec_0_push_valid(io_connPE_14_push_valid),
		.io_connVec_0_push_bits(io_connPE_14_push_bits),
		.io_connVec_0_pop_ready(io_connPE_14_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_14_pop_valid),
		.io_connVec_1_currLength(_taskQueues_14_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_15(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_15_push_ready),
		.io_connVec_0_push_valid(io_connPE_15_push_valid),
		.io_connVec_0_push_bits(io_connPE_15_push_bits),
		.io_connVec_0_pop_ready(io_connPE_15_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_15_pop_valid),
		.io_connVec_1_currLength(_taskQueues_15_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_16(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_16_push_ready),
		.io_connVec_0_push_valid(io_connPE_16_push_valid),
		.io_connVec_0_push_bits(io_connPE_16_push_bits),
		.io_connVec_0_pop_ready(io_connPE_16_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_16_pop_valid),
		.io_connVec_1_currLength(_taskQueues_16_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_16_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_16_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_16_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_16_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_16_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_16_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_17(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_17_push_ready),
		.io_connVec_0_push_valid(io_connPE_17_push_valid),
		.io_connVec_0_push_bits(io_connPE_17_push_bits),
		.io_connVec_0_pop_ready(io_connPE_17_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_17_pop_valid),
		.io_connVec_1_currLength(_taskQueues_17_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_17_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_17_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_17_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_17_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_17_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_17_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_18(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_18_push_ready),
		.io_connVec_0_push_valid(io_connPE_18_push_valid),
		.io_connVec_0_push_bits(io_connPE_18_push_bits),
		.io_connVec_0_pop_ready(io_connPE_18_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_18_pop_valid),
		.io_connVec_1_currLength(_taskQueues_18_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_18_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_18_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_18_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_18_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_18_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_18_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_19(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_19_push_ready),
		.io_connVec_0_push_valid(io_connPE_19_push_valid),
		.io_connVec_0_push_bits(io_connPE_19_push_bits),
		.io_connVec_0_pop_ready(io_connPE_19_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_19_pop_valid),
		.io_connVec_1_currLength(_taskQueues_19_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_19_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_19_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_19_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_19_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_19_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_19_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_20(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_20_push_ready),
		.io_connVec_0_push_valid(io_connPE_20_push_valid),
		.io_connVec_0_push_bits(io_connPE_20_push_bits),
		.io_connVec_0_pop_ready(io_connPE_20_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_20_pop_valid),
		.io_connVec_1_currLength(_taskQueues_20_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_20_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_20_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_20_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_20_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_20_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_20_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_21(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_21_push_ready),
		.io_connVec_0_push_valid(io_connPE_21_push_valid),
		.io_connVec_0_push_bits(io_connPE_21_push_bits),
		.io_connVec_0_pop_ready(io_connPE_21_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_21_pop_valid),
		.io_connVec_1_currLength(_taskQueues_21_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_21_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_21_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_21_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_21_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_21_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_21_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_22(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_22_push_ready),
		.io_connVec_0_push_valid(io_connPE_22_push_valid),
		.io_connVec_0_push_bits(io_connPE_22_push_bits),
		.io_connVec_0_pop_ready(io_connPE_22_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_22_pop_valid),
		.io_connVec_1_currLength(_taskQueues_22_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_22_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_22_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_22_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_22_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_22_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_22_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_23(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_23_push_ready),
		.io_connVec_0_push_valid(io_connPE_23_push_valid),
		.io_connVec_0_push_bits(io_connPE_23_push_bits),
		.io_connVec_0_pop_ready(io_connPE_23_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_23_pop_valid),
		.io_connVec_1_currLength(_taskQueues_23_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_23_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_23_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_23_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_23_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_23_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_23_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_24(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_24_push_ready),
		.io_connVec_0_push_valid(io_connPE_24_push_valid),
		.io_connVec_0_push_bits(io_connPE_24_push_bits),
		.io_connVec_0_pop_ready(io_connPE_24_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_24_pop_valid),
		.io_connVec_1_currLength(_taskQueues_24_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_24_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_24_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_24_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_24_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_24_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_24_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_25(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_25_push_ready),
		.io_connVec_0_push_valid(io_connPE_25_push_valid),
		.io_connVec_0_push_bits(io_connPE_25_push_bits),
		.io_connVec_0_pop_ready(io_connPE_25_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_25_pop_valid),
		.io_connVec_1_currLength(_taskQueues_25_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_25_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_25_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_25_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_25_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_25_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_25_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_26(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_26_push_ready),
		.io_connVec_0_push_valid(io_connPE_26_push_valid),
		.io_connVec_0_push_bits(io_connPE_26_push_bits),
		.io_connVec_0_pop_ready(io_connPE_26_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_26_pop_valid),
		.io_connVec_1_currLength(_taskQueues_26_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_26_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_26_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_26_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_26_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_26_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_26_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_27(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_27_push_ready),
		.io_connVec_0_push_valid(io_connPE_27_push_valid),
		.io_connVec_0_push_bits(io_connPE_27_push_bits),
		.io_connVec_0_pop_ready(io_connPE_27_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_27_pop_valid),
		.io_connVec_1_currLength(_taskQueues_27_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_27_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_27_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_27_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_27_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_27_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_27_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_28(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_28_push_ready),
		.io_connVec_0_push_valid(io_connPE_28_push_valid),
		.io_connVec_0_push_bits(io_connPE_28_push_bits),
		.io_connVec_0_pop_ready(io_connPE_28_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_28_pop_valid),
		.io_connVec_1_currLength(_taskQueues_28_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_28_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_28_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_28_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_28_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_28_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_28_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_29(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_29_push_ready),
		.io_connVec_0_push_valid(io_connPE_29_push_valid),
		.io_connVec_0_push_bits(io_connPE_29_push_bits),
		.io_connVec_0_pop_ready(io_connPE_29_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_29_pop_valid),
		.io_connVec_1_currLength(_taskQueues_29_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_29_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_29_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_29_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_29_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_29_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_29_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_30(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_30_push_ready),
		.io_connVec_0_push_valid(io_connPE_30_push_valid),
		.io_connVec_0_push_bits(io_connPE_30_push_bits),
		.io_connVec_0_pop_ready(io_connPE_30_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_30_pop_valid),
		.io_connVec_1_currLength(_taskQueues_30_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_30_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_30_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_30_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_30_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_30_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_30_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_31(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_31_push_ready),
		.io_connVec_0_push_valid(io_connPE_31_push_valid),
		.io_connVec_0_push_bits(io_connPE_31_push_bits),
		.io_connVec_0_pop_ready(io_connPE_31_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_31_pop_valid),
		.io_connVec_1_currLength(_taskQueues_31_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_31_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_31_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_31_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_31_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_31_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_31_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_32(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_32_push_ready),
		.io_connVec_0_push_valid(io_connPE_32_push_valid),
		.io_connVec_0_push_bits(io_connPE_32_push_bits),
		.io_connVec_0_pop_ready(io_connPE_32_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_32_pop_valid),
		.io_connVec_1_currLength(_taskQueues_32_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_32_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_32_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_32_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_32_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_32_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_32_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_33(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_33_push_ready),
		.io_connVec_0_push_valid(io_connPE_33_push_valid),
		.io_connVec_0_push_bits(io_connPE_33_push_bits),
		.io_connVec_0_pop_ready(io_connPE_33_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_33_pop_valid),
		.io_connVec_1_currLength(_taskQueues_33_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_33_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_33_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_33_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_33_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_33_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_33_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_34(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_34_push_ready),
		.io_connVec_0_push_valid(io_connPE_34_push_valid),
		.io_connVec_0_push_bits(io_connPE_34_push_bits),
		.io_connVec_0_pop_ready(io_connPE_34_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_34_pop_valid),
		.io_connVec_1_currLength(_taskQueues_34_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_34_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_34_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_34_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_34_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_34_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_34_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_35(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_35_push_ready),
		.io_connVec_0_push_valid(io_connPE_35_push_valid),
		.io_connVec_0_push_bits(io_connPE_35_push_bits),
		.io_connVec_0_pop_ready(io_connPE_35_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_35_pop_valid),
		.io_connVec_1_currLength(_taskQueues_35_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_35_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_35_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_35_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_35_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_35_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_35_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_36(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_36_push_ready),
		.io_connVec_0_push_valid(io_connPE_36_push_valid),
		.io_connVec_0_push_bits(io_connPE_36_push_bits),
		.io_connVec_0_pop_ready(io_connPE_36_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_36_pop_valid),
		.io_connVec_1_currLength(_taskQueues_36_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_36_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_36_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_36_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_36_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_36_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_36_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_37(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_37_push_ready),
		.io_connVec_0_push_valid(io_connPE_37_push_valid),
		.io_connVec_0_push_bits(io_connPE_37_push_bits),
		.io_connVec_0_pop_ready(io_connPE_37_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_37_pop_valid),
		.io_connVec_1_currLength(_taskQueues_37_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_37_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_37_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_37_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_37_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_37_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_37_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_38(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_38_push_ready),
		.io_connVec_0_push_valid(io_connPE_38_push_valid),
		.io_connVec_0_push_bits(io_connPE_38_push_bits),
		.io_connVec_0_pop_ready(io_connPE_38_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_38_pop_valid),
		.io_connVec_1_currLength(_taskQueues_38_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_38_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_38_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_38_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_38_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_38_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_38_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_39(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_39_push_ready),
		.io_connVec_0_push_valid(io_connPE_39_push_valid),
		.io_connVec_0_push_bits(io_connPE_39_push_bits),
		.io_connVec_0_pop_ready(io_connPE_39_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_39_pop_valid),
		.io_connVec_1_currLength(_taskQueues_39_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_39_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_39_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_39_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_39_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_39_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_39_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_40(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_40_push_ready),
		.io_connVec_0_push_valid(io_connPE_40_push_valid),
		.io_connVec_0_push_bits(io_connPE_40_push_bits),
		.io_connVec_0_pop_ready(io_connPE_40_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_40_pop_valid),
		.io_connVec_1_currLength(_taskQueues_40_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_40_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_40_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_40_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_40_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_40_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_40_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_41(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_41_push_ready),
		.io_connVec_0_push_valid(io_connPE_41_push_valid),
		.io_connVec_0_push_bits(io_connPE_41_push_bits),
		.io_connVec_0_pop_ready(io_connPE_41_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_41_pop_valid),
		.io_connVec_1_currLength(_taskQueues_41_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_41_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_41_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_41_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_41_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_41_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_41_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_42(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_42_push_ready),
		.io_connVec_0_push_valid(io_connPE_42_push_valid),
		.io_connVec_0_push_bits(io_connPE_42_push_bits),
		.io_connVec_0_pop_ready(io_connPE_42_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_42_pop_valid),
		.io_connVec_1_currLength(_taskQueues_42_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_42_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_42_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_42_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_42_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_42_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_42_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_43(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_43_push_ready),
		.io_connVec_0_push_valid(io_connPE_43_push_valid),
		.io_connVec_0_push_bits(io_connPE_43_push_bits),
		.io_connVec_0_pop_ready(io_connPE_43_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_43_pop_valid),
		.io_connVec_1_currLength(_taskQueues_43_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_43_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_43_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_43_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_43_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_43_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_43_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_44(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_44_push_ready),
		.io_connVec_0_push_valid(io_connPE_44_push_valid),
		.io_connVec_0_push_bits(io_connPE_44_push_bits),
		.io_connVec_0_pop_ready(io_connPE_44_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_44_pop_valid),
		.io_connVec_1_currLength(_taskQueues_44_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_44_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_44_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_44_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_44_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_44_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_44_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_45(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_45_push_ready),
		.io_connVec_0_push_valid(io_connPE_45_push_valid),
		.io_connVec_0_push_bits(io_connPE_45_push_bits),
		.io_connVec_0_pop_ready(io_connPE_45_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_45_pop_valid),
		.io_connVec_1_currLength(_taskQueues_45_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_45_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_45_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_45_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_45_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_45_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_45_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_46(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_46_push_ready),
		.io_connVec_0_push_valid(io_connPE_46_push_valid),
		.io_connVec_0_push_bits(io_connPE_46_push_bits),
		.io_connVec_0_pop_ready(io_connPE_46_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_46_pop_valid),
		.io_connVec_1_currLength(_taskQueues_46_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_46_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_46_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_46_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_46_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_46_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_46_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_47(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_47_push_ready),
		.io_connVec_0_push_valid(io_connPE_47_push_valid),
		.io_connVec_0_push_bits(io_connPE_47_push_bits),
		.io_connVec_0_pop_ready(io_connPE_47_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_47_pop_valid),
		.io_connVec_1_currLength(_taskQueues_47_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_47_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_47_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_47_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_47_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_47_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_47_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_48(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_48_push_ready),
		.io_connVec_0_push_valid(io_connPE_48_push_valid),
		.io_connVec_0_push_bits(io_connPE_48_push_bits),
		.io_connVec_0_pop_ready(io_connPE_48_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_48_pop_valid),
		.io_connVec_1_currLength(_taskQueues_48_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_48_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_48_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_48_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_48_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_48_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_48_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_49(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_49_push_ready),
		.io_connVec_0_push_valid(io_connPE_49_push_valid),
		.io_connVec_0_push_bits(io_connPE_49_push_bits),
		.io_connVec_0_pop_ready(io_connPE_49_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_49_pop_valid),
		.io_connVec_1_currLength(_taskQueues_49_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_49_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_49_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_49_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_49_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_49_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_49_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_50(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_50_push_ready),
		.io_connVec_0_push_valid(io_connPE_50_push_valid),
		.io_connVec_0_push_bits(io_connPE_50_push_bits),
		.io_connVec_0_pop_ready(io_connPE_50_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_50_pop_valid),
		.io_connVec_1_currLength(_taskQueues_50_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_50_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_50_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_50_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_50_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_50_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_50_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_51(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_51_push_ready),
		.io_connVec_0_push_valid(io_connPE_51_push_valid),
		.io_connVec_0_push_bits(io_connPE_51_push_bits),
		.io_connVec_0_pop_ready(io_connPE_51_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_51_pop_valid),
		.io_connVec_1_currLength(_taskQueues_51_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_51_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_51_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_51_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_51_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_51_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_51_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_52(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_52_push_ready),
		.io_connVec_0_push_valid(io_connPE_52_push_valid),
		.io_connVec_0_push_bits(io_connPE_52_push_bits),
		.io_connVec_0_pop_ready(io_connPE_52_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_52_pop_valid),
		.io_connVec_1_currLength(_taskQueues_52_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_52_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_52_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_52_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_52_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_52_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_52_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_53(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_53_push_ready),
		.io_connVec_0_push_valid(io_connPE_53_push_valid),
		.io_connVec_0_push_bits(io_connPE_53_push_bits),
		.io_connVec_0_pop_ready(io_connPE_53_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_53_pop_valid),
		.io_connVec_1_currLength(_taskQueues_53_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_53_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_53_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_53_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_53_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_53_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_53_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_54(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_54_push_ready),
		.io_connVec_0_push_valid(io_connPE_54_push_valid),
		.io_connVec_0_push_bits(io_connPE_54_push_bits),
		.io_connVec_0_pop_ready(io_connPE_54_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_54_pop_valid),
		.io_connVec_1_currLength(_taskQueues_54_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_54_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_54_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_54_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_54_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_54_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_54_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_55(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_55_push_ready),
		.io_connVec_0_push_valid(io_connPE_55_push_valid),
		.io_connVec_0_push_bits(io_connPE_55_push_bits),
		.io_connVec_0_pop_ready(io_connPE_55_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_55_pop_valid),
		.io_connVec_1_currLength(_taskQueues_55_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_55_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_55_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_55_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_55_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_55_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_55_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_56(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_56_push_ready),
		.io_connVec_0_push_valid(io_connPE_56_push_valid),
		.io_connVec_0_push_bits(io_connPE_56_push_bits),
		.io_connVec_0_pop_ready(io_connPE_56_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_56_pop_valid),
		.io_connVec_1_currLength(_taskQueues_56_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_56_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_56_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_56_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_56_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_56_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_56_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_57(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_57_push_ready),
		.io_connVec_0_push_valid(io_connPE_57_push_valid),
		.io_connVec_0_push_bits(io_connPE_57_push_bits),
		.io_connVec_0_pop_ready(io_connPE_57_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_57_pop_valid),
		.io_connVec_1_currLength(_taskQueues_57_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_57_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_57_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_57_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_57_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_57_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_57_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_58(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_58_push_ready),
		.io_connVec_0_push_valid(io_connPE_58_push_valid),
		.io_connVec_0_push_bits(io_connPE_58_push_bits),
		.io_connVec_0_pop_ready(io_connPE_58_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_58_pop_valid),
		.io_connVec_1_currLength(_taskQueues_58_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_58_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_58_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_58_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_58_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_58_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_58_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_59(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_59_push_ready),
		.io_connVec_0_push_valid(io_connPE_59_push_valid),
		.io_connVec_0_push_bits(io_connPE_59_push_bits),
		.io_connVec_0_pop_ready(io_connPE_59_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_59_pop_valid),
		.io_connVec_1_currLength(_taskQueues_59_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_59_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_59_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_59_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_59_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_59_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_59_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_60(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_60_push_ready),
		.io_connVec_0_push_valid(io_connPE_60_push_valid),
		.io_connVec_0_push_bits(io_connPE_60_push_bits),
		.io_connVec_0_pop_ready(io_connPE_60_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_60_pop_valid),
		.io_connVec_1_currLength(_taskQueues_60_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_60_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_60_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_60_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_60_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_60_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_60_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_61(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_61_push_ready),
		.io_connVec_0_push_valid(io_connPE_61_push_valid),
		.io_connVec_0_push_bits(io_connPE_61_push_bits),
		.io_connVec_0_pop_ready(io_connPE_61_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_61_pop_valid),
		.io_connVec_1_currLength(_taskQueues_61_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_61_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_61_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_61_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_61_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_61_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_61_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_62(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_62_push_ready),
		.io_connVec_0_push_valid(io_connPE_62_push_valid),
		.io_connVec_0_push_bits(io_connPE_62_push_bits),
		.io_connVec_0_pop_ready(io_connPE_62_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_62_pop_valid),
		.io_connVec_1_currLength(_taskQueues_62_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_62_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_62_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_62_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_62_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_62_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_62_io_connVec_1_pop_bits)
	);
	hw_deque taskQueues_63(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_push_ready(io_connPE_63_push_ready),
		.io_connVec_0_push_valid(io_connPE_63_push_valid),
		.io_connVec_0_push_bits(io_connPE_63_push_bits),
		.io_connVec_0_pop_ready(io_connPE_63_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_63_pop_valid),
		.io_connVec_1_currLength(_taskQueues_63_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_63_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_63_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_63_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_63_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_63_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_63_io_connVec_1_pop_bits)
	);
endmodule
module ram_2x9 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [8:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [8:0] W0_data;
	reg [8:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 9'bxxxxxxxxx);
endmodule
module Queue2_AddressChannel_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_prot,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_prot
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [5:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_prot;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [5:0] io_deq_bits_addr;
	output wire [2:0] io_deq_bits_prot;
	wire [8:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x9 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({io_enq_bits_prot, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[5:0];
	assign io_deq_bits_prot = _ram_ext_R0_data[8:6];
endmodule
module Queue1_AddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_prot,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [5:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_prot;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [5:0] io_deq_bits_addr;
	reg [8:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_prot, io_enq_bits_addr};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_addr = ram[5:0];
endmodule
module Queue1_ReadDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	reg [65:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {2'h0, io_enq_bits_data};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[63:0];
	assign io_deq_bits_resp = ram[65:64];
endmodule
module Queue1_WriteDataChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [7:0] io_enq_bits_strb;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [7:0] io_deq_bits_strb;
	reg [71:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= {io_enq_bits_strb, io_enq_bits_data};
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
	assign io_deq_bits_data = ram[63:0];
	assign io_deq_bits_strb = ram[71:64];
endmodule
module Queue1_WriteResponseChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_deq_ready,
	io_deq_valid
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_deq_ready;
	output wire io_deq_valid;
	reg full;
	always @(posedge clock)
		if (reset)
			full <= 1'h0;
		else begin : sv2v_autoblock_1
			reg do_enq;
			do_enq = ~full & io_enq_valid;
			if (~(do_enq == (io_deq_ready & full)))
				full <= do_enq;
		end
	assign io_enq_ready = ~full;
	assign io_deq_valid = full;
endmodule
module Queue1_UInt (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_bits,
	io_count
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [255:0] io_enq_bits;
	input io_deq_ready;
	output wire [255:0] io_deq_bits;
	output wire io_count;
	reg [255:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= io_enq_bits;
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_bits = ram;
	assign io_count = full;
endmodule
module SchedulerServer (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_axi_mgmt_ar_ready,
	io_axi_mgmt_ar_valid,
	io_axi_mgmt_ar_bits_addr,
	io_axi_mgmt_ar_bits_prot,
	io_axi_mgmt_r_ready,
	io_axi_mgmt_r_valid,
	io_axi_mgmt_r_bits_data,
	io_axi_mgmt_r_bits_resp,
	io_axi_mgmt_aw_ready,
	io_axi_mgmt_aw_valid,
	io_axi_mgmt_aw_bits_addr,
	io_axi_mgmt_aw_bits_prot,
	io_axi_mgmt_w_ready,
	io_axi_mgmt_w_valid,
	io_axi_mgmt_w_bits_data,
	io_axi_mgmt_w_bits_strb,
	io_axi_mgmt_b_ready,
	io_axi_mgmt_b_valid,
	io_axi_mgmt_b_bits_resp,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_read_burst_len,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_write_last,
	io_ntwDataUnitOccupancy
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [255:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [255:0] io_connNetwork_data_qOutTask_bits;
	output wire io_axi_mgmt_ar_ready;
	input io_axi_mgmt_ar_valid;
	input [5:0] io_axi_mgmt_ar_bits_addr;
	input [2:0] io_axi_mgmt_ar_bits_prot;
	input io_axi_mgmt_r_ready;
	output wire io_axi_mgmt_r_valid;
	output wire [63:0] io_axi_mgmt_r_bits_data;
	output wire [1:0] io_axi_mgmt_r_bits_resp;
	output wire io_axi_mgmt_aw_ready;
	input io_axi_mgmt_aw_valid;
	input [5:0] io_axi_mgmt_aw_bits_addr;
	input [2:0] io_axi_mgmt_aw_bits_prot;
	output wire io_axi_mgmt_w_ready;
	input io_axi_mgmt_w_valid;
	input [63:0] io_axi_mgmt_w_bits_data;
	input [7:0] io_axi_mgmt_w_bits_strb;
	input io_axi_mgmt_b_ready;
	output wire io_axi_mgmt_b_valid;
	output wire [1:0] io_axi_mgmt_b_bits_resp;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [255:0] io_read_data_bits;
	output wire [3:0] io_read_burst_len;
	input io_write_address_ready;
	output wire io_write_address_valid;
	output wire [63:0] io_write_address_bits;
	input io_write_data_ready;
	output wire io_write_data_valid;
	output wire [255:0] io_write_data_bits;
	output wire io_write_last;
	input io_ntwDataUnitOccupancy;
	wire [63:0] currLen;
	wire _taskQueueBuffer_io_enq_ready;
	wire [255:0] _taskQueueBuffer_io_deq_bits;
	wire _taskQueueBuffer_io_count;
	wire _wrRespQueue__io_enq_ready;
	wire _wrRespQueue__io_deq_valid;
	wire _wrReqData__deq_q_io_enq_ready;
	wire _wrReqData__deq_q_io_deq_valid;
	wire [63:0] _wrReqData__deq_q_io_deq_bits_data;
	wire [7:0] _wrReqData__deq_q_io_deq_bits_strb;
	wire _wrReq__deq_q_io_enq_ready;
	wire _wrReq__deq_q_io_deq_valid;
	wire [5:0] _wrReq__deq_q_io_deq_bits_addr;
	wire _rdRespQueue__io_enq_ready;
	wire _rdRespQueue__io_deq_valid;
	wire [63:0] _rdRespQueue__io_deq_bits_data;
	wire [1:0] _rdRespQueue__io_deq_bits_resp;
	wire _rdReq__deq_q_io_enq_ready;
	wire _rdReq__deq_q_io_deq_valid;
	wire [5:0] _rdReq__deq_q_io_deq_bits_addr;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	wire rdReq = _rdReq__deq_q_io_deq_valid & _rdRespQueue__io_enq_ready;
	wire wrReq = (_wrReq__deq_q_io_deq_valid & _wrReqData__deq_q_io_deq_valid) & _wrRespQueue__io_enq_ready;
	reg [63:0] rAddr;
	reg [63:0] rPause;
	reg [63:0] procInterrupt;
	reg [63:0] maxLength;
	reg [3:0] stateReg;
	reg [63:0] contentionCounter;
	reg networkCongested;
	reg [63:0] fifoTailReg;
	reg [63:0] fifoHeadReg;
	reg popOrPush;
	reg [4:0] memDataCounter;
	wire _GEN = stateReg == 4'h2;
	wire _GEN_0 = stateReg == 4'h4;
	wire _GEN_1 = stateReg == 4'h3;
	wire _GEN_2 = memDataCounter == 5'h01;
	wire _GEN_3 = _GEN | _GEN_0;
	wire _GEN_4 = stateReg == 4'h6;
	wire _GEN_5 = stateReg == 4'h5;
	wire _GEN_6 = (_GEN_0 | _GEN_1) | _GEN_4;
	wire _GEN_7 = _GEN | _GEN_6;
	wire _GEN_8 = stateReg == 4'h7;
	wire _GEN_9 = (_GEN | _GEN_0) | _GEN_1;
	wire _GEN_10 = _GEN_4 | _GEN_5;
	reg [63:0] lengthHistroy;
	wire _GEN_11 = fifoTailReg > fifoHeadReg;
	wire [63:0] _currLen_T = fifoTailReg - fifoHeadReg;
	wire _GEN_12 = fifoTailReg < fifoHeadReg;
	wire [63:0] _currLen_T_4 = (maxLength - fifoHeadReg) + fifoTailReg;
	wire [63:0] _currLen_T_6 = lengthHistroy + 64'h0000000000000001;
	assign currLen = (_GEN_11 ? _currLen_T : (_GEN_12 ? _currLen_T_4 : (popOrPush ? 64'h0000000000000000 : _currLen_T_6)));
	wire [511:0] _GEN_13 = {128'hffffffffffffffffffffffffffffffff, procInterrupt, fifoHeadReg, fifoTailReg, maxLength, rAddr, rPause};
	always @(posedge clock)
		if (reset) begin
			rAddr <= 64'h0000000000000000;
			rPause <= 64'h0000000000000000;
			procInterrupt <= 64'h0000000000000000;
			maxLength <= 64'h0000000000000000;
			stateReg <= 4'h0;
			contentionCounter <= 64'h0000000000000000;
			networkCongested <= 1'h0;
			fifoTailReg <= 64'h0000000000000000;
			fifoHeadReg <= 64'h0000000000000000;
			popOrPush <= 1'h1;
			memDataCounter <= 5'h00;
			lengthHistroy <= 64'h0000000000000000;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_14;
			reg _GEN_15;
			reg _GEN_16;
			reg [63:0] _GEN_17;
			reg _GEN_18;
			reg _GEN_19;
			reg _GEN_20;
			reg [63:0] _GEN_21;
			_GEN_20 = rPause == 64'h0000000000000000;
			_GEN_14 = stateReg == 4'h0;
			_GEN_15 = ((currLen == maxLength) & networkCongested) | (maxLength < (currLen + 64'h0000000000000001));
			_GEN_16 = io_write_data_ready & _GEN_2;
			_GEN_17 = maxLength - 64'h0000000000000001;
			_GEN_18 = _GEN_14 | _GEN_3;
			_GEN_19 = io_read_data_valid & _GEN_2;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h1))
				rAddr <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rAddr[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rAddr[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rAddr[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rAddr[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rAddr[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rAddr[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rAddr[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rAddr[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h0))
				rPause <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rPause[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rPause[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rPause[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rPause[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rPause[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rPause[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rPause[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rPause[7:0])};
			else if (_GEN_14 & (|procInterrupt | _GEN_15))
				rPause <= 64'hffffffffffffffff;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h5))
				procInterrupt <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : procInterrupt[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : procInterrupt[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : procInterrupt[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : procInterrupt[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : procInterrupt[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : procInterrupt[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : procInterrupt[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : procInterrupt[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h2))
				maxLength <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : maxLength[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : maxLength[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : maxLength[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : maxLength[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : maxLength[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : maxLength[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : maxLength[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : maxLength[7:0])};
			_GEN_21 = {stateReg, stateReg, stateReg, stateReg, stateReg, (_GEN_20 ? 4'h0 : 4'ha), (_GEN_20 ? 4'h0 : 4'h9), (io_connNetwork_ctrl_serveStealReq_ready ? 4'h7 : (networkCongested | (|procInterrupt) ? 4'h0 : stateReg)), (io_connNetwork_data_qOutTask_ready | networkCongested ? 4'h0 : 4'h7), (io_read_address_ready ? 4'h5 : stateReg), (_GEN_19 ? 4'h8 : stateReg), (io_write_address_ready ? 4'h3 : stateReg), (_GEN_16 ? 4'h0 : stateReg), (~_taskQueueBuffer_io_count & io_connNetwork_data_availableTask_valid ? 4'h4 : (io_connNetwork_data_availableTask_valid & networkCongested ? 4'h2 : (networkCongested ? stateReg : 4'h0))), stateReg, (|procInterrupt ? 4'ha : (_GEN_15 ? 4'h9 : (networkCongested & _taskQueueBuffer_io_count ? 4'h4 : (networkCongested ? 4'h2 : ((~networkCongested & |currLen) & ~_taskQueueBuffer_io_count ? 4'h6 : (~networkCongested & _taskQueueBuffer_io_count ? 4'h7 : stateReg))))))};
			stateReg <= _GEN_21[stateReg * 4+:4];
			if ((~io_connNetwork_ctrl_serveStealReq_ready & io_ntwDataUnitOccupancy) & (contentionCounter != 64'h0000000000000040))
				contentionCounter <= contentionCounter + 64'h0000000000000001;
			else if ((io_connNetwork_ctrl_serveStealReq_ready & |contentionCounter) & ~io_ntwDataUnitOccupancy)
				contentionCounter <= contentionCounter - 64'h0000000000000001;
			networkCongested <= (contentionCounter > 64'h0000000000000035) | ((contentionCounter > 64'h0000000000000033) & networkCongested);
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h3))
				fifoTailReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoTailReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoTailReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoTailReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoTailReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoTailReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoTailReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoTailReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoTailReg[7:0])};
			else if (_GEN_18 | ~_GEN_1)
				;
			else begin : sv2v_autoblock_2
				reg _GEN_22;
				_GEN_22 = fifoTailReg < _GEN_17;
				if (_GEN_16) begin
					if (_GEN_22)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
				else if (io_write_data_ready) begin
					if (_GEN_22)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
			end
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h4))
				fifoHeadReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoHeadReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoHeadReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoHeadReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoHeadReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoHeadReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoHeadReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoHeadReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoHeadReg[7:0])};
			else if ((_GEN_14 | _GEN_7) | ~_GEN_5)
				;
			else begin : sv2v_autoblock_3
				reg _GEN_23;
				_GEN_23 = fifoHeadReg < _GEN_17;
				if (_GEN_19) begin
					if (_GEN_23)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
				else if (io_read_data_valid) begin
					if (_GEN_23)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
			end
			if (~_GEN_18) begin
				if (_GEN_1)
					popOrPush <= ~_GEN_16 & popOrPush;
				else
					popOrPush <= ((~_GEN_4 & _GEN_5) & _GEN_19) | popOrPush;
			end
			if (~(_GEN_14 | _GEN)) begin
				if (_GEN_0) begin
					if (io_write_address_ready)
						memDataCounter <= 5'h01;
				end
				else if (_GEN_1) begin
					if (_GEN_16 | ~io_write_data_ready)
						;
					else
						memDataCounter <= memDataCounter - 5'h01;
				end
				else if (_GEN_4) begin
					if (io_read_address_ready)
						memDataCounter <= (currLen == 64'h0000000000000000 ? currLen[4:0] : 5'h01);
				end
				else if ((~_GEN_5 | _GEN_19) | ~io_read_data_valid)
					;
				else
					memDataCounter <= memDataCounter - 5'h01;
			end
			if (_GEN_11 | _GEN_12) begin
				if (_GEN_11)
					lengthHistroy <= _currLen_T;
				else if (_GEN_12)
					lengthHistroy <= _currLen_T_4;
				else if (popOrPush)
					lengthHistroy <= 64'h0000000000000000;
				else
					lengthHistroy <= _currLen_T_6;
			end
		end
	Queue2_AddressChannel_2 s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_ar_ready),
		.io_enq_valid(io_axi_mgmt_ar_valid),
		.io_enq_bits_addr(io_axi_mgmt_ar_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_ar_bits_prot),
		.io_deq_ready(_rdReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_rdRespQueue__io_deq_valid),
		.io_enq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_enq_bits_resp(_rdRespQueue__io_deq_bits_resp),
		.io_deq_ready(io_axi_mgmt_r_ready),
		.io_deq_valid(io_axi_mgmt_r_valid),
		.io_deq_bits_data(io_axi_mgmt_r_bits_data),
		.io_deq_bits_resp(io_axi_mgmt_r_bits_resp)
	);
	Queue2_AddressChannel_2 s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_aw_ready),
		.io_enq_valid(io_axi_mgmt_aw_valid),
		.io_enq_bits_addr(io_axi_mgmt_aw_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_aw_bits_prot),
		.io_deq_ready(_wrReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_w_ready),
		.io_enq_valid(io_axi_mgmt_w_valid),
		.io_enq_bits_data(io_axi_mgmt_w_bits_data),
		.io_enq_bits_strb(io_axi_mgmt_w_bits_strb),
		.io_deq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_wrRespQueue__io_deq_valid),
		.io_enq_bits_resp(2'h0),
		.io_deq_ready(io_axi_mgmt_b_ready),
		.io_deq_valid(io_axi_mgmt_b_valid),
		.io_deq_bits_resp(io_axi_mgmt_b_bits_resp)
	);
	Queue1_AddressChannel rdReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_deq_ready(rdReq),
		.io_deq_valid(_rdReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_rdReq__deq_q_io_deq_bits_addr)
	);
	Queue1_ReadDataChannel rdRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdRespQueue__io_enq_ready),
		.io_enq_valid(rdReq),
		.io_enq_bits_data(_GEN_13[_rdReq__deq_q_io_deq_bits_addr[5:3] * 64+:64]),
		.io_deq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_deq_valid(_rdRespQueue__io_deq_valid),
		.io_deq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_deq_bits_resp(_rdRespQueue__io_deq_bits_resp)
	);
	Queue1_AddressChannel wrReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_wrReq__deq_q_io_deq_bits_addr)
	);
	Queue1_WriteDataChannel wrReqData__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_enq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_enq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReqData__deq_q_io_deq_valid),
		.io_deq_bits_data(_wrReqData__deq_q_io_deq_bits_data),
		.io_deq_bits_strb(_wrReqData__deq_q_io_deq_bits_strb)
	);
	Queue1_WriteResponseChannel wrRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrRespQueue__io_enq_ready),
		.io_enq_valid(wrReq),
		.io_deq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_deq_valid(_wrRespQueue__io_deq_valid)
	);
	Queue1_UInt taskQueueBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_taskQueueBuffer_io_enq_ready),
		.io_enq_valid((_GEN ? io_connNetwork_data_availableTask_valid : (~_GEN_6 & _GEN_5) & io_read_data_valid)),
		.io_enq_bits((_GEN ? io_connNetwork_data_availableTask_bits : (_GEN_6 | ~_GEN_5 ? 256'h0000000000000000000000000000000000000000000000000000000000000000 : io_read_data_bits))),
		.io_deq_ready(~_GEN_3 & (_GEN_1 ? io_write_data_ready : (~_GEN_10 & _GEN_8) & io_connNetwork_data_qOutTask_ready)),
		.io_deq_bits(_taskQueueBuffer_io_deq_bits),
		.io_count(_taskQueueBuffer_io_count)
	);
	assign io_connNetwork_ctrl_serveStealReq_valid = ~(((((_GEN | _GEN_0) | _GEN_1) | _GEN_4) | _GEN_5) | _GEN_8) & (stateReg == 4'h8);
	assign io_connNetwork_data_availableTask_ready = _GEN & _taskQueueBuffer_io_enq_ready;
	assign io_connNetwork_data_qOutTask_valid = ~(((_GEN | _GEN_0) | _GEN_1) | _GEN_10) & _GEN_8;
	assign io_connNetwork_data_qOutTask_bits = _taskQueueBuffer_io_deq_bits;
	assign io_read_address_valid = ~_GEN_9 & _GEN_4;
	assign io_read_address_bits = (_GEN_9 | ~_GEN_4 ? 64'h0000000000000000 : {fifoHeadReg[58:0], 5'h00} + rAddr);
	assign io_read_data_ready = ~_GEN_7 & _GEN_5;
	assign io_read_burst_len = (_GEN_9 | ~(_GEN_4 & (currLen == 64'h0000000000000000)) ? 4'h0 : currLen[3:0] - 4'h1);
	assign io_write_address_valid = ~_GEN & _GEN_0;
	assign io_write_address_bits = (_GEN | ~_GEN_0 ? 64'h0000000000000000 : {fifoTailReg[58:0], 5'h00} + rAddr);
	assign io_write_data_valid = ~_GEN_3 & _GEN_1;
	assign io_write_data_bits = _taskQueueBuffer_io_deq_bits;
	assign io_write_last = (~_GEN_3 & _GEN_1) & _GEN_2;
endmodule
module RVtoAXIBridge (
	clock,
	reset,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_writeBurst_last,
	io_readBurst_len,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_ar_bits_len,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data,
	axi_aw_ready,
	axi_aw_valid,
	axi_aw_bits_addr,
	axi_w_ready,
	axi_w_valid,
	axi_w_bits_data,
	axi_w_bits_last,
	axi_b_valid
);
	input clock;
	input reset;
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [255:0] io_read_data_bits;
	output wire io_write_address_ready;
	input io_write_address_valid;
	input [63:0] io_write_address_bits;
	output wire io_write_data_ready;
	input io_write_data_valid;
	input [255:0] io_write_data_bits;
	input io_writeBurst_last;
	input [3:0] io_readBurst_len;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire [7:0] axi_ar_bits_len;
	output wire axi_r_ready;
	input axi_r_valid;
	input [255:0] axi_r_bits_data;
	input axi_aw_ready;
	output wire axi_aw_valid;
	output wire [63:0] axi_aw_bits_addr;
	input axi_w_ready;
	output wire axi_w_valid;
	output wire [255:0] axi_w_bits_data;
	output wire axi_w_bits_last;
	input axi_b_valid;
	reg writeHandshakeDetector;
	wire axi_w_valid_0 = (io_write_data_valid & axi_w_ready) & ~writeHandshakeDetector;
	always @(posedge clock)
		if (reset)
			writeHandshakeDetector <= 1'h0;
		else if (axi_w_valid_0)
			writeHandshakeDetector <= io_writeBurst_last | writeHandshakeDetector;
		else
			writeHandshakeDetector <= ~axi_b_valid & writeHandshakeDetector;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign io_write_address_ready = axi_aw_ready;
	assign io_write_data_ready = axi_w_ready & ~writeHandshakeDetector;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_ar_bits_len = {4'h0, io_readBurst_len};
	assign axi_r_ready = io_read_data_ready;
	assign axi_aw_valid = io_write_address_valid;
	assign axi_aw_bits_addr = io_write_address_bits;
	assign axi_w_valid = axi_w_valid_0;
	assign axi_w_bits_data = io_write_data_bits;
	assign axi_w_bits_last = io_writeBurst_last;
endmodule
module Counter (
	clock,
	reset,
	io_incEn,
	io_decEn,
	io_empty,
	io_full
);
	input clock;
	input reset;
	input io_incEn;
	input io_decEn;
	output wire io_empty;
	output wire io_full;
	reg [1:0] rCounter;
	always @(posedge clock)
		if (reset)
			rCounter <= 2'h0;
		else if (~(io_incEn & io_decEn)) begin
			if (io_incEn)
				rCounter <= rCounter + 2'h1;
			else if (io_decEn)
				rCounter <= rCounter - 2'h1;
		end
	assign io_empty = rCounter == 2'h0;
	assign io_full = &rCounter;
endmodule
module ram_2x93 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [92:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [92:0] W0_data;
	reg [92:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 93'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue2_WriteAddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_size,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input [2:0] io_enq_bits_size;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [92:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x93 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({18'h00001, io_enq_bits_size, 8'h00, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[63:0];
	assign io_deq_bits_len = _ram_ext_R0_data[71:64];
	assign io_deq_bits_size = _ram_ext_R0_data[74:72];
	assign io_deq_bits_burst = _ram_ext_R0_data[76:75];
	assign io_deq_bits_lock = _ram_ext_R0_data[77];
	assign io_deq_bits_cache = _ram_ext_R0_data[81:78];
	assign io_deq_bits_prot = _ram_ext_R0_data[84:82];
	assign io_deq_bits_qos = _ram_ext_R0_data[88:85];
	assign io_deq_bits_region = _ram_ext_R0_data[92:89];
endmodule
module Queue2_ReadAddressChannel (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst,
	io_deq_bits_lock,
	io_deq_bits_cache,
	io_deq_bits_prot,
	io_deq_bits_qos,
	io_deq_bits_region
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	output wire io_deq_bits_lock;
	output wire [3:0] io_deq_bits_cache;
	output wire [2:0] io_deq_bits_prot;
	output wire [3:0] io_deq_bits_qos;
	output wire [3:0] io_deq_bits_region;
	wire [92:0] _ram_ext_R0_data;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_2x93 ram_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(_ram_ext_R0_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data({18'h00001, io_enq_bits_size, io_enq_bits_len, io_enq_bits_addr})
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
	assign io_deq_bits_addr = _ram_ext_R0_data[63:0];
	assign io_deq_bits_len = _ram_ext_R0_data[71:64];
	assign io_deq_bits_size = _ram_ext_R0_data[74:72];
	assign io_deq_bits_burst = _ram_ext_R0_data[76:75];
	assign io_deq_bits_lock = _ram_ext_R0_data[77];
	assign io_deq_bits_cache = _ram_ext_R0_data[81:78];
	assign io_deq_bits_prot = _ram_ext_R0_data[84:82];
	assign io_deq_bits_qos = _ram_ext_R0_data[88:85];
	assign io_deq_bits_region = _ram_ext_R0_data[92:89];
endmodule
module AxiWriteBuffer (
	clock,
	reset,
	s_axi_ar_ready,
	s_axi_ar_valid,
	s_axi_ar_bits_addr,
	s_axi_ar_bits_len,
	s_axi_r_ready,
	s_axi_r_valid,
	s_axi_r_bits_data,
	s_axi_aw_ready,
	s_axi_aw_valid,
	s_axi_aw_bits_addr,
	s_axi_w_ready,
	s_axi_w_valid,
	s_axi_w_bits_data,
	s_axi_w_bits_last,
	s_axi_b_valid,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_data,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_last,
	m_axi_b_valid
);
	input clock;
	input reset;
	output wire s_axi_ar_ready;
	input s_axi_ar_valid;
	input [63:0] s_axi_ar_bits_addr;
	input [7:0] s_axi_ar_bits_len;
	input s_axi_r_ready;
	output wire s_axi_r_valid;
	output wire [255:0] s_axi_r_bits_data;
	output wire s_axi_aw_ready;
	input s_axi_aw_valid;
	input [63:0] s_axi_aw_bits_addr;
	output wire s_axi_w_ready;
	input s_axi_w_valid;
	input [255:0] s_axi_w_bits_data;
	input s_axi_w_bits_last;
	output wire s_axi_b_valid;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [255:0] m_axi_r_bits_data;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [255:0] m_axi_w_bits_data;
	output wire m_axi_w_bits_last;
	input m_axi_b_valid;
	wire s_axi_aw_ready_0;
	wire _sinkBuffered__sinkBuffer_1_io_enq_ready;
	wire _sinkBuffered__sinkBuffer_io_enq_ready;
	wire _counter_io_empty;
	wire _counter_io_full;
	wire _counter_io_incEn_T = s_axi_aw_ready_0 & s_axi_aw_valid;
	assign s_axi_aw_ready_0 = (_sinkBuffered__sinkBuffer_io_enq_ready & s_axi_aw_valid) & ~_counter_io_full;
	wire s_axi_ar_ready_0 = ((_sinkBuffered__sinkBuffer_1_io_enq_ready & s_axi_ar_valid) & _counter_io_empty) & ~_counter_io_incEn_T;
	Counter counter(
		.clock(clock),
		.reset(reset),
		.io_incEn(_counter_io_incEn_T),
		.io_decEn(m_axi_b_valid),
		.io_empty(_counter_io_empty),
		.io_full(_counter_io_full)
	);
	Queue2_WriteAddressChannel sinkBuffered__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_io_enq_ready),
		.io_enq_valid(s_axi_aw_ready_0),
		.io_enq_bits_addr(s_axi_aw_bits_addr),
		.io_enq_bits_size(3'h5),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_ReadAddressChannel sinkBuffered__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(s_axi_ar_ready_0),
		.io_enq_bits_addr(s_axi_ar_bits_addr),
		.io_enq_bits_len(s_axi_ar_bits_len),
		.io_enq_bits_size(3'h5),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	assign s_axi_ar_ready = s_axi_ar_ready_0;
	assign s_axi_r_valid = m_axi_r_valid;
	assign s_axi_r_bits_data = m_axi_r_bits_data;
	assign s_axi_aw_ready = s_axi_aw_ready_0;
	assign s_axi_w_ready = m_axi_w_ready;
	assign s_axi_b_valid = m_axi_b_valid;
	assign m_axi_r_ready = s_axi_r_ready;
	assign m_axi_w_valid = s_axi_w_valid;
	assign m_axi_w_bits_data = s_axi_w_bits_data;
	assign m_axi_w_bits_last = s_axi_w_bits_last;
endmodule
module AxisDownscaler (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataOut_TREADY,
	io_dataOut_TVALID
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	reg writeCounter;
	always @(posedge clock)
		if (reset)
			writeCounter <= 1'h0;
		else
			writeCounter <= ~io_dataIn_TVALID & writeCounter;
	assign io_dataIn_TREADY = 1'h1;
	assign io_dataOut_TVALID = 1'h0;
endmodule
module AxisDataWidthConverter (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataOut_TREADY,
	io_dataOut_TVALID
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	AxisDownscaler downScaler(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_dataIn_TREADY),
		.io_dataIn_TVALID(io_dataIn_TVALID),
		.io_dataOut_TREADY(io_dataOut_TREADY),
		.io_dataOut_TVALID(io_dataOut_TVALID)
	);
endmodule
module AxisUpscaler (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [31:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [255:0] io_dataOut_TDATA;
	reg [255:0] buffer;
	reg readCounter;
	reg stateReg;
	always @(posedge clock)
		if (reset) begin
			buffer <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			readCounter <= 1'h0;
			stateReg <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg _GEN;
			_GEN = stateReg & io_dataOut_TREADY;
			if (stateReg | ~io_dataIn_TVALID)
				;
			else
				buffer <= {buffer[255:159], buffer[158:0] | ({127'h00000000000000000000000000000000, io_dataIn_TDATA} << {153'h000000000000000000000000000000000000000, readCounter, 5'h00})};
			if (stateReg)
				readCounter <= ~_GEN & readCounter;
			else if (io_dataIn_TVALID)
				readCounter <= readCounter - 1'h1;
			stateReg <= (~stateReg | ~_GEN) & stateReg;
		end
	assign io_dataIn_TREADY = ~stateReg;
	assign io_dataOut_TVALID = stateReg;
	assign io_dataOut_TDATA = buffer;
endmodule
module AxisDataWidthConverter_64 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [31:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [255:0] io_dataOut_TDATA;
	AxisUpscaler upScaler(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_dataIn_TREADY),
		.io_dataIn_TVALID(io_dataIn_TVALID),
		.io_dataIn_TDATA(io_dataIn_TDATA),
		.io_dataOut_TREADY(io_dataOut_TREADY),
		.io_dataOut_TVALID(io_dataOut_TVALID),
		.io_dataOut_TDATA(io_dataOut_TDATA)
	);
endmodule
module Scheduler (
	clock,
	reset,
	io_export_taskOut_0_TREADY,
	io_export_taskOut_0_TVALID,
	io_export_taskOut_1_TREADY,
	io_export_taskOut_1_TVALID,
	io_export_taskOut_2_TREADY,
	io_export_taskOut_2_TVALID,
	io_export_taskOut_3_TREADY,
	io_export_taskOut_3_TVALID,
	io_export_taskOut_4_TREADY,
	io_export_taskOut_4_TVALID,
	io_export_taskOut_5_TREADY,
	io_export_taskOut_5_TVALID,
	io_export_taskOut_6_TREADY,
	io_export_taskOut_6_TVALID,
	io_export_taskOut_7_TREADY,
	io_export_taskOut_7_TVALID,
	io_export_taskOut_8_TREADY,
	io_export_taskOut_8_TVALID,
	io_export_taskOut_9_TREADY,
	io_export_taskOut_9_TVALID,
	io_export_taskOut_10_TREADY,
	io_export_taskOut_10_TVALID,
	io_export_taskOut_11_TREADY,
	io_export_taskOut_11_TVALID,
	io_export_taskOut_12_TREADY,
	io_export_taskOut_12_TVALID,
	io_export_taskOut_13_TREADY,
	io_export_taskOut_13_TVALID,
	io_export_taskOut_14_TREADY,
	io_export_taskOut_14_TVALID,
	io_export_taskOut_15_TREADY,
	io_export_taskOut_15_TVALID,
	io_export_taskOut_16_TREADY,
	io_export_taskOut_16_TVALID,
	io_export_taskOut_17_TREADY,
	io_export_taskOut_17_TVALID,
	io_export_taskOut_18_TREADY,
	io_export_taskOut_18_TVALID,
	io_export_taskOut_19_TREADY,
	io_export_taskOut_19_TVALID,
	io_export_taskOut_20_TREADY,
	io_export_taskOut_20_TVALID,
	io_export_taskOut_21_TREADY,
	io_export_taskOut_21_TVALID,
	io_export_taskOut_22_TREADY,
	io_export_taskOut_22_TVALID,
	io_export_taskOut_23_TREADY,
	io_export_taskOut_23_TVALID,
	io_export_taskOut_24_TREADY,
	io_export_taskOut_24_TVALID,
	io_export_taskOut_25_TREADY,
	io_export_taskOut_25_TVALID,
	io_export_taskOut_26_TREADY,
	io_export_taskOut_26_TVALID,
	io_export_taskOut_27_TREADY,
	io_export_taskOut_27_TVALID,
	io_export_taskOut_28_TREADY,
	io_export_taskOut_28_TVALID,
	io_export_taskOut_29_TREADY,
	io_export_taskOut_29_TVALID,
	io_export_taskOut_30_TREADY,
	io_export_taskOut_30_TVALID,
	io_export_taskOut_31_TREADY,
	io_export_taskOut_31_TVALID,
	io_export_taskOut_32_TREADY,
	io_export_taskOut_32_TVALID,
	io_export_taskOut_33_TREADY,
	io_export_taskOut_33_TVALID,
	io_export_taskOut_34_TREADY,
	io_export_taskOut_34_TVALID,
	io_export_taskOut_35_TREADY,
	io_export_taskOut_35_TVALID,
	io_export_taskOut_36_TREADY,
	io_export_taskOut_36_TVALID,
	io_export_taskOut_37_TREADY,
	io_export_taskOut_37_TVALID,
	io_export_taskOut_38_TREADY,
	io_export_taskOut_38_TVALID,
	io_export_taskOut_39_TREADY,
	io_export_taskOut_39_TVALID,
	io_export_taskOut_40_TREADY,
	io_export_taskOut_40_TVALID,
	io_export_taskOut_41_TREADY,
	io_export_taskOut_41_TVALID,
	io_export_taskOut_42_TREADY,
	io_export_taskOut_42_TVALID,
	io_export_taskOut_43_TREADY,
	io_export_taskOut_43_TVALID,
	io_export_taskOut_44_TREADY,
	io_export_taskOut_44_TVALID,
	io_export_taskOut_45_TREADY,
	io_export_taskOut_45_TVALID,
	io_export_taskOut_46_TREADY,
	io_export_taskOut_46_TVALID,
	io_export_taskOut_47_TREADY,
	io_export_taskOut_47_TVALID,
	io_export_taskOut_48_TREADY,
	io_export_taskOut_48_TVALID,
	io_export_taskOut_49_TREADY,
	io_export_taskOut_49_TVALID,
	io_export_taskOut_50_TREADY,
	io_export_taskOut_50_TVALID,
	io_export_taskOut_51_TREADY,
	io_export_taskOut_51_TVALID,
	io_export_taskOut_52_TREADY,
	io_export_taskOut_52_TVALID,
	io_export_taskOut_53_TREADY,
	io_export_taskOut_53_TVALID,
	io_export_taskOut_54_TREADY,
	io_export_taskOut_54_TVALID,
	io_export_taskOut_55_TREADY,
	io_export_taskOut_55_TVALID,
	io_export_taskOut_56_TREADY,
	io_export_taskOut_56_TVALID,
	io_export_taskOut_57_TREADY,
	io_export_taskOut_57_TVALID,
	io_export_taskOut_58_TREADY,
	io_export_taskOut_58_TVALID,
	io_export_taskOut_59_TREADY,
	io_export_taskOut_59_TVALID,
	io_export_taskOut_60_TREADY,
	io_export_taskOut_60_TVALID,
	io_export_taskOut_61_TREADY,
	io_export_taskOut_61_TVALID,
	io_export_taskOut_62_TREADY,
	io_export_taskOut_62_TVALID,
	io_export_taskOut_63_TREADY,
	io_export_taskOut_63_TVALID,
	io_export_taskIn_0_TREADY,
	io_export_taskIn_0_TVALID,
	io_export_taskIn_0_TDATA,
	io_export_taskIn_1_TREADY,
	io_export_taskIn_1_TVALID,
	io_export_taskIn_1_TDATA,
	io_export_taskIn_2_TREADY,
	io_export_taskIn_2_TVALID,
	io_export_taskIn_2_TDATA,
	io_export_taskIn_3_TREADY,
	io_export_taskIn_3_TVALID,
	io_export_taskIn_3_TDATA,
	io_export_taskIn_4_TREADY,
	io_export_taskIn_4_TVALID,
	io_export_taskIn_4_TDATA,
	io_export_taskIn_5_TREADY,
	io_export_taskIn_5_TVALID,
	io_export_taskIn_5_TDATA,
	io_export_taskIn_6_TREADY,
	io_export_taskIn_6_TVALID,
	io_export_taskIn_6_TDATA,
	io_export_taskIn_7_TREADY,
	io_export_taskIn_7_TVALID,
	io_export_taskIn_7_TDATA,
	io_export_taskIn_8_TREADY,
	io_export_taskIn_8_TVALID,
	io_export_taskIn_8_TDATA,
	io_export_taskIn_9_TREADY,
	io_export_taskIn_9_TVALID,
	io_export_taskIn_9_TDATA,
	io_export_taskIn_10_TREADY,
	io_export_taskIn_10_TVALID,
	io_export_taskIn_10_TDATA,
	io_export_taskIn_11_TREADY,
	io_export_taskIn_11_TVALID,
	io_export_taskIn_11_TDATA,
	io_export_taskIn_12_TREADY,
	io_export_taskIn_12_TVALID,
	io_export_taskIn_12_TDATA,
	io_export_taskIn_13_TREADY,
	io_export_taskIn_13_TVALID,
	io_export_taskIn_13_TDATA,
	io_export_taskIn_14_TREADY,
	io_export_taskIn_14_TVALID,
	io_export_taskIn_14_TDATA,
	io_export_taskIn_15_TREADY,
	io_export_taskIn_15_TVALID,
	io_export_taskIn_15_TDATA,
	io_export_taskIn_16_TREADY,
	io_export_taskIn_16_TVALID,
	io_export_taskIn_16_TDATA,
	io_export_taskIn_17_TREADY,
	io_export_taskIn_17_TVALID,
	io_export_taskIn_17_TDATA,
	io_export_taskIn_18_TREADY,
	io_export_taskIn_18_TVALID,
	io_export_taskIn_18_TDATA,
	io_export_taskIn_19_TREADY,
	io_export_taskIn_19_TVALID,
	io_export_taskIn_19_TDATA,
	io_export_taskIn_20_TREADY,
	io_export_taskIn_20_TVALID,
	io_export_taskIn_20_TDATA,
	io_export_taskIn_21_TREADY,
	io_export_taskIn_21_TVALID,
	io_export_taskIn_21_TDATA,
	io_export_taskIn_22_TREADY,
	io_export_taskIn_22_TVALID,
	io_export_taskIn_22_TDATA,
	io_export_taskIn_23_TREADY,
	io_export_taskIn_23_TVALID,
	io_export_taskIn_23_TDATA,
	io_export_taskIn_24_TREADY,
	io_export_taskIn_24_TVALID,
	io_export_taskIn_24_TDATA,
	io_export_taskIn_25_TREADY,
	io_export_taskIn_25_TVALID,
	io_export_taskIn_25_TDATA,
	io_export_taskIn_26_TREADY,
	io_export_taskIn_26_TVALID,
	io_export_taskIn_26_TDATA,
	io_export_taskIn_27_TREADY,
	io_export_taskIn_27_TVALID,
	io_export_taskIn_27_TDATA,
	io_export_taskIn_28_TREADY,
	io_export_taskIn_28_TVALID,
	io_export_taskIn_28_TDATA,
	io_export_taskIn_29_TREADY,
	io_export_taskIn_29_TVALID,
	io_export_taskIn_29_TDATA,
	io_export_taskIn_30_TREADY,
	io_export_taskIn_30_TVALID,
	io_export_taskIn_30_TDATA,
	io_export_taskIn_31_TREADY,
	io_export_taskIn_31_TVALID,
	io_export_taskIn_31_TDATA,
	io_export_taskIn_32_TREADY,
	io_export_taskIn_32_TVALID,
	io_export_taskIn_32_TDATA,
	io_export_taskIn_33_TREADY,
	io_export_taskIn_33_TVALID,
	io_export_taskIn_33_TDATA,
	io_export_taskIn_34_TREADY,
	io_export_taskIn_34_TVALID,
	io_export_taskIn_34_TDATA,
	io_export_taskIn_35_TREADY,
	io_export_taskIn_35_TVALID,
	io_export_taskIn_35_TDATA,
	io_export_taskIn_36_TREADY,
	io_export_taskIn_36_TVALID,
	io_export_taskIn_36_TDATA,
	io_export_taskIn_37_TREADY,
	io_export_taskIn_37_TVALID,
	io_export_taskIn_37_TDATA,
	io_export_taskIn_38_TREADY,
	io_export_taskIn_38_TVALID,
	io_export_taskIn_38_TDATA,
	io_export_taskIn_39_TREADY,
	io_export_taskIn_39_TVALID,
	io_export_taskIn_39_TDATA,
	io_export_taskIn_40_TREADY,
	io_export_taskIn_40_TVALID,
	io_export_taskIn_40_TDATA,
	io_export_taskIn_41_TREADY,
	io_export_taskIn_41_TVALID,
	io_export_taskIn_41_TDATA,
	io_export_taskIn_42_TREADY,
	io_export_taskIn_42_TVALID,
	io_export_taskIn_42_TDATA,
	io_export_taskIn_43_TREADY,
	io_export_taskIn_43_TVALID,
	io_export_taskIn_43_TDATA,
	io_export_taskIn_44_TREADY,
	io_export_taskIn_44_TVALID,
	io_export_taskIn_44_TDATA,
	io_export_taskIn_45_TREADY,
	io_export_taskIn_45_TVALID,
	io_export_taskIn_45_TDATA,
	io_export_taskIn_46_TREADY,
	io_export_taskIn_46_TVALID,
	io_export_taskIn_46_TDATA,
	io_export_taskIn_47_TREADY,
	io_export_taskIn_47_TVALID,
	io_export_taskIn_47_TDATA,
	io_export_taskIn_48_TREADY,
	io_export_taskIn_48_TVALID,
	io_export_taskIn_48_TDATA,
	io_export_taskIn_49_TREADY,
	io_export_taskIn_49_TVALID,
	io_export_taskIn_49_TDATA,
	io_export_taskIn_50_TREADY,
	io_export_taskIn_50_TVALID,
	io_export_taskIn_50_TDATA,
	io_export_taskIn_51_TREADY,
	io_export_taskIn_51_TVALID,
	io_export_taskIn_51_TDATA,
	io_export_taskIn_52_TREADY,
	io_export_taskIn_52_TVALID,
	io_export_taskIn_52_TDATA,
	io_export_taskIn_53_TREADY,
	io_export_taskIn_53_TVALID,
	io_export_taskIn_53_TDATA,
	io_export_taskIn_54_TREADY,
	io_export_taskIn_54_TVALID,
	io_export_taskIn_54_TDATA,
	io_export_taskIn_55_TREADY,
	io_export_taskIn_55_TVALID,
	io_export_taskIn_55_TDATA,
	io_export_taskIn_56_TREADY,
	io_export_taskIn_56_TVALID,
	io_export_taskIn_56_TDATA,
	io_export_taskIn_57_TREADY,
	io_export_taskIn_57_TVALID,
	io_export_taskIn_57_TDATA,
	io_export_taskIn_58_TREADY,
	io_export_taskIn_58_TVALID,
	io_export_taskIn_58_TDATA,
	io_export_taskIn_59_TREADY,
	io_export_taskIn_59_TVALID,
	io_export_taskIn_59_TDATA,
	io_export_taskIn_60_TREADY,
	io_export_taskIn_60_TVALID,
	io_export_taskIn_60_TDATA,
	io_export_taskIn_61_TREADY,
	io_export_taskIn_61_TVALID,
	io_export_taskIn_61_TDATA,
	io_export_taskIn_62_TREADY,
	io_export_taskIn_62_TVALID,
	io_export_taskIn_62_TDATA,
	io_export_taskIn_63_TREADY,
	io_export_taskIn_63_TVALID,
	io_export_taskIn_63_TDATA,
	io_internal_vss_axi_full_0_ar_ready,
	io_internal_vss_axi_full_0_ar_valid,
	io_internal_vss_axi_full_0_ar_bits_addr,
	io_internal_vss_axi_full_0_ar_bits_len,
	io_internal_vss_axi_full_0_ar_bits_size,
	io_internal_vss_axi_full_0_ar_bits_burst,
	io_internal_vss_axi_full_0_ar_bits_lock,
	io_internal_vss_axi_full_0_ar_bits_cache,
	io_internal_vss_axi_full_0_ar_bits_prot,
	io_internal_vss_axi_full_0_ar_bits_qos,
	io_internal_vss_axi_full_0_ar_bits_region,
	io_internal_vss_axi_full_0_r_ready,
	io_internal_vss_axi_full_0_r_valid,
	io_internal_vss_axi_full_0_r_bits_data,
	io_internal_vss_axi_full_0_aw_ready,
	io_internal_vss_axi_full_0_aw_valid,
	io_internal_vss_axi_full_0_aw_bits_addr,
	io_internal_vss_axi_full_0_aw_bits_len,
	io_internal_vss_axi_full_0_aw_bits_size,
	io_internal_vss_axi_full_0_aw_bits_burst,
	io_internal_vss_axi_full_0_aw_bits_lock,
	io_internal_vss_axi_full_0_aw_bits_cache,
	io_internal_vss_axi_full_0_aw_bits_prot,
	io_internal_vss_axi_full_0_aw_bits_qos,
	io_internal_vss_axi_full_0_aw_bits_region,
	io_internal_vss_axi_full_0_w_ready,
	io_internal_vss_axi_full_0_w_valid,
	io_internal_vss_axi_full_0_w_bits_data,
	io_internal_vss_axi_full_0_w_bits_last,
	io_internal_vss_axi_full_0_b_valid,
	io_internal_axi_mgmt_vss_0_ar_ready,
	io_internal_axi_mgmt_vss_0_ar_valid,
	io_internal_axi_mgmt_vss_0_ar_bits_addr,
	io_internal_axi_mgmt_vss_0_ar_bits_prot,
	io_internal_axi_mgmt_vss_0_r_ready,
	io_internal_axi_mgmt_vss_0_r_valid,
	io_internal_axi_mgmt_vss_0_r_bits_data,
	io_internal_axi_mgmt_vss_0_r_bits_resp,
	io_internal_axi_mgmt_vss_0_aw_ready,
	io_internal_axi_mgmt_vss_0_aw_valid,
	io_internal_axi_mgmt_vss_0_aw_bits_addr,
	io_internal_axi_mgmt_vss_0_aw_bits_prot,
	io_internal_axi_mgmt_vss_0_w_ready,
	io_internal_axi_mgmt_vss_0_w_valid,
	io_internal_axi_mgmt_vss_0_w_bits_data,
	io_internal_axi_mgmt_vss_0_w_bits_strb,
	io_internal_axi_mgmt_vss_0_b_ready,
	io_internal_axi_mgmt_vss_0_b_valid,
	io_internal_axi_mgmt_vss_0_b_bits_resp
);
	input clock;
	input reset;
	input io_export_taskOut_0_TREADY;
	output wire io_export_taskOut_0_TVALID;
	input io_export_taskOut_1_TREADY;
	output wire io_export_taskOut_1_TVALID;
	input io_export_taskOut_2_TREADY;
	output wire io_export_taskOut_2_TVALID;
	input io_export_taskOut_3_TREADY;
	output wire io_export_taskOut_3_TVALID;
	input io_export_taskOut_4_TREADY;
	output wire io_export_taskOut_4_TVALID;
	input io_export_taskOut_5_TREADY;
	output wire io_export_taskOut_5_TVALID;
	input io_export_taskOut_6_TREADY;
	output wire io_export_taskOut_6_TVALID;
	input io_export_taskOut_7_TREADY;
	output wire io_export_taskOut_7_TVALID;
	input io_export_taskOut_8_TREADY;
	output wire io_export_taskOut_8_TVALID;
	input io_export_taskOut_9_TREADY;
	output wire io_export_taskOut_9_TVALID;
	input io_export_taskOut_10_TREADY;
	output wire io_export_taskOut_10_TVALID;
	input io_export_taskOut_11_TREADY;
	output wire io_export_taskOut_11_TVALID;
	input io_export_taskOut_12_TREADY;
	output wire io_export_taskOut_12_TVALID;
	input io_export_taskOut_13_TREADY;
	output wire io_export_taskOut_13_TVALID;
	input io_export_taskOut_14_TREADY;
	output wire io_export_taskOut_14_TVALID;
	input io_export_taskOut_15_TREADY;
	output wire io_export_taskOut_15_TVALID;
	input io_export_taskOut_16_TREADY;
	output wire io_export_taskOut_16_TVALID;
	input io_export_taskOut_17_TREADY;
	output wire io_export_taskOut_17_TVALID;
	input io_export_taskOut_18_TREADY;
	output wire io_export_taskOut_18_TVALID;
	input io_export_taskOut_19_TREADY;
	output wire io_export_taskOut_19_TVALID;
	input io_export_taskOut_20_TREADY;
	output wire io_export_taskOut_20_TVALID;
	input io_export_taskOut_21_TREADY;
	output wire io_export_taskOut_21_TVALID;
	input io_export_taskOut_22_TREADY;
	output wire io_export_taskOut_22_TVALID;
	input io_export_taskOut_23_TREADY;
	output wire io_export_taskOut_23_TVALID;
	input io_export_taskOut_24_TREADY;
	output wire io_export_taskOut_24_TVALID;
	input io_export_taskOut_25_TREADY;
	output wire io_export_taskOut_25_TVALID;
	input io_export_taskOut_26_TREADY;
	output wire io_export_taskOut_26_TVALID;
	input io_export_taskOut_27_TREADY;
	output wire io_export_taskOut_27_TVALID;
	input io_export_taskOut_28_TREADY;
	output wire io_export_taskOut_28_TVALID;
	input io_export_taskOut_29_TREADY;
	output wire io_export_taskOut_29_TVALID;
	input io_export_taskOut_30_TREADY;
	output wire io_export_taskOut_30_TVALID;
	input io_export_taskOut_31_TREADY;
	output wire io_export_taskOut_31_TVALID;
	input io_export_taskOut_32_TREADY;
	output wire io_export_taskOut_32_TVALID;
	input io_export_taskOut_33_TREADY;
	output wire io_export_taskOut_33_TVALID;
	input io_export_taskOut_34_TREADY;
	output wire io_export_taskOut_34_TVALID;
	input io_export_taskOut_35_TREADY;
	output wire io_export_taskOut_35_TVALID;
	input io_export_taskOut_36_TREADY;
	output wire io_export_taskOut_36_TVALID;
	input io_export_taskOut_37_TREADY;
	output wire io_export_taskOut_37_TVALID;
	input io_export_taskOut_38_TREADY;
	output wire io_export_taskOut_38_TVALID;
	input io_export_taskOut_39_TREADY;
	output wire io_export_taskOut_39_TVALID;
	input io_export_taskOut_40_TREADY;
	output wire io_export_taskOut_40_TVALID;
	input io_export_taskOut_41_TREADY;
	output wire io_export_taskOut_41_TVALID;
	input io_export_taskOut_42_TREADY;
	output wire io_export_taskOut_42_TVALID;
	input io_export_taskOut_43_TREADY;
	output wire io_export_taskOut_43_TVALID;
	input io_export_taskOut_44_TREADY;
	output wire io_export_taskOut_44_TVALID;
	input io_export_taskOut_45_TREADY;
	output wire io_export_taskOut_45_TVALID;
	input io_export_taskOut_46_TREADY;
	output wire io_export_taskOut_46_TVALID;
	input io_export_taskOut_47_TREADY;
	output wire io_export_taskOut_47_TVALID;
	input io_export_taskOut_48_TREADY;
	output wire io_export_taskOut_48_TVALID;
	input io_export_taskOut_49_TREADY;
	output wire io_export_taskOut_49_TVALID;
	input io_export_taskOut_50_TREADY;
	output wire io_export_taskOut_50_TVALID;
	input io_export_taskOut_51_TREADY;
	output wire io_export_taskOut_51_TVALID;
	input io_export_taskOut_52_TREADY;
	output wire io_export_taskOut_52_TVALID;
	input io_export_taskOut_53_TREADY;
	output wire io_export_taskOut_53_TVALID;
	input io_export_taskOut_54_TREADY;
	output wire io_export_taskOut_54_TVALID;
	input io_export_taskOut_55_TREADY;
	output wire io_export_taskOut_55_TVALID;
	input io_export_taskOut_56_TREADY;
	output wire io_export_taskOut_56_TVALID;
	input io_export_taskOut_57_TREADY;
	output wire io_export_taskOut_57_TVALID;
	input io_export_taskOut_58_TREADY;
	output wire io_export_taskOut_58_TVALID;
	input io_export_taskOut_59_TREADY;
	output wire io_export_taskOut_59_TVALID;
	input io_export_taskOut_60_TREADY;
	output wire io_export_taskOut_60_TVALID;
	input io_export_taskOut_61_TREADY;
	output wire io_export_taskOut_61_TVALID;
	input io_export_taskOut_62_TREADY;
	output wire io_export_taskOut_62_TVALID;
	input io_export_taskOut_63_TREADY;
	output wire io_export_taskOut_63_TVALID;
	output wire io_export_taskIn_0_TREADY;
	input io_export_taskIn_0_TVALID;
	input [31:0] io_export_taskIn_0_TDATA;
	output wire io_export_taskIn_1_TREADY;
	input io_export_taskIn_1_TVALID;
	input [31:0] io_export_taskIn_1_TDATA;
	output wire io_export_taskIn_2_TREADY;
	input io_export_taskIn_2_TVALID;
	input [31:0] io_export_taskIn_2_TDATA;
	output wire io_export_taskIn_3_TREADY;
	input io_export_taskIn_3_TVALID;
	input [31:0] io_export_taskIn_3_TDATA;
	output wire io_export_taskIn_4_TREADY;
	input io_export_taskIn_4_TVALID;
	input [31:0] io_export_taskIn_4_TDATA;
	output wire io_export_taskIn_5_TREADY;
	input io_export_taskIn_5_TVALID;
	input [31:0] io_export_taskIn_5_TDATA;
	output wire io_export_taskIn_6_TREADY;
	input io_export_taskIn_6_TVALID;
	input [31:0] io_export_taskIn_6_TDATA;
	output wire io_export_taskIn_7_TREADY;
	input io_export_taskIn_7_TVALID;
	input [31:0] io_export_taskIn_7_TDATA;
	output wire io_export_taskIn_8_TREADY;
	input io_export_taskIn_8_TVALID;
	input [31:0] io_export_taskIn_8_TDATA;
	output wire io_export_taskIn_9_TREADY;
	input io_export_taskIn_9_TVALID;
	input [31:0] io_export_taskIn_9_TDATA;
	output wire io_export_taskIn_10_TREADY;
	input io_export_taskIn_10_TVALID;
	input [31:0] io_export_taskIn_10_TDATA;
	output wire io_export_taskIn_11_TREADY;
	input io_export_taskIn_11_TVALID;
	input [31:0] io_export_taskIn_11_TDATA;
	output wire io_export_taskIn_12_TREADY;
	input io_export_taskIn_12_TVALID;
	input [31:0] io_export_taskIn_12_TDATA;
	output wire io_export_taskIn_13_TREADY;
	input io_export_taskIn_13_TVALID;
	input [31:0] io_export_taskIn_13_TDATA;
	output wire io_export_taskIn_14_TREADY;
	input io_export_taskIn_14_TVALID;
	input [31:0] io_export_taskIn_14_TDATA;
	output wire io_export_taskIn_15_TREADY;
	input io_export_taskIn_15_TVALID;
	input [31:0] io_export_taskIn_15_TDATA;
	output wire io_export_taskIn_16_TREADY;
	input io_export_taskIn_16_TVALID;
	input [31:0] io_export_taskIn_16_TDATA;
	output wire io_export_taskIn_17_TREADY;
	input io_export_taskIn_17_TVALID;
	input [31:0] io_export_taskIn_17_TDATA;
	output wire io_export_taskIn_18_TREADY;
	input io_export_taskIn_18_TVALID;
	input [31:0] io_export_taskIn_18_TDATA;
	output wire io_export_taskIn_19_TREADY;
	input io_export_taskIn_19_TVALID;
	input [31:0] io_export_taskIn_19_TDATA;
	output wire io_export_taskIn_20_TREADY;
	input io_export_taskIn_20_TVALID;
	input [31:0] io_export_taskIn_20_TDATA;
	output wire io_export_taskIn_21_TREADY;
	input io_export_taskIn_21_TVALID;
	input [31:0] io_export_taskIn_21_TDATA;
	output wire io_export_taskIn_22_TREADY;
	input io_export_taskIn_22_TVALID;
	input [31:0] io_export_taskIn_22_TDATA;
	output wire io_export_taskIn_23_TREADY;
	input io_export_taskIn_23_TVALID;
	input [31:0] io_export_taskIn_23_TDATA;
	output wire io_export_taskIn_24_TREADY;
	input io_export_taskIn_24_TVALID;
	input [31:0] io_export_taskIn_24_TDATA;
	output wire io_export_taskIn_25_TREADY;
	input io_export_taskIn_25_TVALID;
	input [31:0] io_export_taskIn_25_TDATA;
	output wire io_export_taskIn_26_TREADY;
	input io_export_taskIn_26_TVALID;
	input [31:0] io_export_taskIn_26_TDATA;
	output wire io_export_taskIn_27_TREADY;
	input io_export_taskIn_27_TVALID;
	input [31:0] io_export_taskIn_27_TDATA;
	output wire io_export_taskIn_28_TREADY;
	input io_export_taskIn_28_TVALID;
	input [31:0] io_export_taskIn_28_TDATA;
	output wire io_export_taskIn_29_TREADY;
	input io_export_taskIn_29_TVALID;
	input [31:0] io_export_taskIn_29_TDATA;
	output wire io_export_taskIn_30_TREADY;
	input io_export_taskIn_30_TVALID;
	input [31:0] io_export_taskIn_30_TDATA;
	output wire io_export_taskIn_31_TREADY;
	input io_export_taskIn_31_TVALID;
	input [31:0] io_export_taskIn_31_TDATA;
	output wire io_export_taskIn_32_TREADY;
	input io_export_taskIn_32_TVALID;
	input [31:0] io_export_taskIn_32_TDATA;
	output wire io_export_taskIn_33_TREADY;
	input io_export_taskIn_33_TVALID;
	input [31:0] io_export_taskIn_33_TDATA;
	output wire io_export_taskIn_34_TREADY;
	input io_export_taskIn_34_TVALID;
	input [31:0] io_export_taskIn_34_TDATA;
	output wire io_export_taskIn_35_TREADY;
	input io_export_taskIn_35_TVALID;
	input [31:0] io_export_taskIn_35_TDATA;
	output wire io_export_taskIn_36_TREADY;
	input io_export_taskIn_36_TVALID;
	input [31:0] io_export_taskIn_36_TDATA;
	output wire io_export_taskIn_37_TREADY;
	input io_export_taskIn_37_TVALID;
	input [31:0] io_export_taskIn_37_TDATA;
	output wire io_export_taskIn_38_TREADY;
	input io_export_taskIn_38_TVALID;
	input [31:0] io_export_taskIn_38_TDATA;
	output wire io_export_taskIn_39_TREADY;
	input io_export_taskIn_39_TVALID;
	input [31:0] io_export_taskIn_39_TDATA;
	output wire io_export_taskIn_40_TREADY;
	input io_export_taskIn_40_TVALID;
	input [31:0] io_export_taskIn_40_TDATA;
	output wire io_export_taskIn_41_TREADY;
	input io_export_taskIn_41_TVALID;
	input [31:0] io_export_taskIn_41_TDATA;
	output wire io_export_taskIn_42_TREADY;
	input io_export_taskIn_42_TVALID;
	input [31:0] io_export_taskIn_42_TDATA;
	output wire io_export_taskIn_43_TREADY;
	input io_export_taskIn_43_TVALID;
	input [31:0] io_export_taskIn_43_TDATA;
	output wire io_export_taskIn_44_TREADY;
	input io_export_taskIn_44_TVALID;
	input [31:0] io_export_taskIn_44_TDATA;
	output wire io_export_taskIn_45_TREADY;
	input io_export_taskIn_45_TVALID;
	input [31:0] io_export_taskIn_45_TDATA;
	output wire io_export_taskIn_46_TREADY;
	input io_export_taskIn_46_TVALID;
	input [31:0] io_export_taskIn_46_TDATA;
	output wire io_export_taskIn_47_TREADY;
	input io_export_taskIn_47_TVALID;
	input [31:0] io_export_taskIn_47_TDATA;
	output wire io_export_taskIn_48_TREADY;
	input io_export_taskIn_48_TVALID;
	input [31:0] io_export_taskIn_48_TDATA;
	output wire io_export_taskIn_49_TREADY;
	input io_export_taskIn_49_TVALID;
	input [31:0] io_export_taskIn_49_TDATA;
	output wire io_export_taskIn_50_TREADY;
	input io_export_taskIn_50_TVALID;
	input [31:0] io_export_taskIn_50_TDATA;
	output wire io_export_taskIn_51_TREADY;
	input io_export_taskIn_51_TVALID;
	input [31:0] io_export_taskIn_51_TDATA;
	output wire io_export_taskIn_52_TREADY;
	input io_export_taskIn_52_TVALID;
	input [31:0] io_export_taskIn_52_TDATA;
	output wire io_export_taskIn_53_TREADY;
	input io_export_taskIn_53_TVALID;
	input [31:0] io_export_taskIn_53_TDATA;
	output wire io_export_taskIn_54_TREADY;
	input io_export_taskIn_54_TVALID;
	input [31:0] io_export_taskIn_54_TDATA;
	output wire io_export_taskIn_55_TREADY;
	input io_export_taskIn_55_TVALID;
	input [31:0] io_export_taskIn_55_TDATA;
	output wire io_export_taskIn_56_TREADY;
	input io_export_taskIn_56_TVALID;
	input [31:0] io_export_taskIn_56_TDATA;
	output wire io_export_taskIn_57_TREADY;
	input io_export_taskIn_57_TVALID;
	input [31:0] io_export_taskIn_57_TDATA;
	output wire io_export_taskIn_58_TREADY;
	input io_export_taskIn_58_TVALID;
	input [31:0] io_export_taskIn_58_TDATA;
	output wire io_export_taskIn_59_TREADY;
	input io_export_taskIn_59_TVALID;
	input [31:0] io_export_taskIn_59_TDATA;
	output wire io_export_taskIn_60_TREADY;
	input io_export_taskIn_60_TVALID;
	input [31:0] io_export_taskIn_60_TDATA;
	output wire io_export_taskIn_61_TREADY;
	input io_export_taskIn_61_TVALID;
	input [31:0] io_export_taskIn_61_TDATA;
	output wire io_export_taskIn_62_TREADY;
	input io_export_taskIn_62_TVALID;
	input [31:0] io_export_taskIn_62_TDATA;
	output wire io_export_taskIn_63_TREADY;
	input io_export_taskIn_63_TVALID;
	input [31:0] io_export_taskIn_63_TDATA;
	input io_internal_vss_axi_full_0_ar_ready;
	output wire io_internal_vss_axi_full_0_ar_valid;
	output wire [63:0] io_internal_vss_axi_full_0_ar_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_ar_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_ar_bits_burst;
	output wire io_internal_vss_axi_full_0_ar_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_region;
	output wire io_internal_vss_axi_full_0_r_ready;
	input io_internal_vss_axi_full_0_r_valid;
	input [255:0] io_internal_vss_axi_full_0_r_bits_data;
	input io_internal_vss_axi_full_0_aw_ready;
	output wire io_internal_vss_axi_full_0_aw_valid;
	output wire [63:0] io_internal_vss_axi_full_0_aw_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_aw_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_aw_bits_burst;
	output wire io_internal_vss_axi_full_0_aw_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_region;
	input io_internal_vss_axi_full_0_w_ready;
	output wire io_internal_vss_axi_full_0_w_valid;
	output wire [255:0] io_internal_vss_axi_full_0_w_bits_data;
	output wire io_internal_vss_axi_full_0_w_bits_last;
	input io_internal_vss_axi_full_0_b_valid;
	output wire io_internal_axi_mgmt_vss_0_ar_ready;
	input io_internal_axi_mgmt_vss_0_ar_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_ar_bits_prot;
	input io_internal_axi_mgmt_vss_0_r_ready;
	output wire io_internal_axi_mgmt_vss_0_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vss_0_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vss_0_r_bits_resp;
	output wire io_internal_axi_mgmt_vss_0_aw_ready;
	input io_internal_axi_mgmt_vss_0_aw_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_aw_bits_prot;
	output wire io_internal_axi_mgmt_vss_0_w_ready;
	input io_internal_axi_mgmt_vss_0_w_valid;
	input [63:0] io_internal_axi_mgmt_vss_0_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vss_0_w_bits_strb;
	input io_internal_axi_mgmt_vss_0_b_ready;
	output wire io_internal_axi_mgmt_vss_0_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vss_0_b_bits_resp;
	wire _axis_stream_converters_in_63_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_63_io_dataOut_TDATA;
	wire _axis_stream_converters_in_62_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_62_io_dataOut_TDATA;
	wire _axis_stream_converters_in_61_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_61_io_dataOut_TDATA;
	wire _axis_stream_converters_in_60_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_60_io_dataOut_TDATA;
	wire _axis_stream_converters_in_59_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_59_io_dataOut_TDATA;
	wire _axis_stream_converters_in_58_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_58_io_dataOut_TDATA;
	wire _axis_stream_converters_in_57_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_57_io_dataOut_TDATA;
	wire _axis_stream_converters_in_56_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_56_io_dataOut_TDATA;
	wire _axis_stream_converters_in_55_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_55_io_dataOut_TDATA;
	wire _axis_stream_converters_in_54_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_54_io_dataOut_TDATA;
	wire _axis_stream_converters_in_53_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_53_io_dataOut_TDATA;
	wire _axis_stream_converters_in_52_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_52_io_dataOut_TDATA;
	wire _axis_stream_converters_in_51_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_51_io_dataOut_TDATA;
	wire _axis_stream_converters_in_50_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_50_io_dataOut_TDATA;
	wire _axis_stream_converters_in_49_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_49_io_dataOut_TDATA;
	wire _axis_stream_converters_in_48_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_48_io_dataOut_TDATA;
	wire _axis_stream_converters_in_47_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_47_io_dataOut_TDATA;
	wire _axis_stream_converters_in_46_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_46_io_dataOut_TDATA;
	wire _axis_stream_converters_in_45_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_45_io_dataOut_TDATA;
	wire _axis_stream_converters_in_44_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_44_io_dataOut_TDATA;
	wire _axis_stream_converters_in_43_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_43_io_dataOut_TDATA;
	wire _axis_stream_converters_in_42_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_42_io_dataOut_TDATA;
	wire _axis_stream_converters_in_41_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_41_io_dataOut_TDATA;
	wire _axis_stream_converters_in_40_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_40_io_dataOut_TDATA;
	wire _axis_stream_converters_in_39_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_39_io_dataOut_TDATA;
	wire _axis_stream_converters_in_38_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_38_io_dataOut_TDATA;
	wire _axis_stream_converters_in_37_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_37_io_dataOut_TDATA;
	wire _axis_stream_converters_in_36_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_36_io_dataOut_TDATA;
	wire _axis_stream_converters_in_35_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_35_io_dataOut_TDATA;
	wire _axis_stream_converters_in_34_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_34_io_dataOut_TDATA;
	wire _axis_stream_converters_in_33_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_33_io_dataOut_TDATA;
	wire _axis_stream_converters_in_32_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_32_io_dataOut_TDATA;
	wire _axis_stream_converters_in_31_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_31_io_dataOut_TDATA;
	wire _axis_stream_converters_in_30_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_30_io_dataOut_TDATA;
	wire _axis_stream_converters_in_29_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_29_io_dataOut_TDATA;
	wire _axis_stream_converters_in_28_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_28_io_dataOut_TDATA;
	wire _axis_stream_converters_in_27_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_27_io_dataOut_TDATA;
	wire _axis_stream_converters_in_26_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_26_io_dataOut_TDATA;
	wire _axis_stream_converters_in_25_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_25_io_dataOut_TDATA;
	wire _axis_stream_converters_in_24_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_24_io_dataOut_TDATA;
	wire _axis_stream_converters_in_23_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_23_io_dataOut_TDATA;
	wire _axis_stream_converters_in_22_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_22_io_dataOut_TDATA;
	wire _axis_stream_converters_in_21_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_21_io_dataOut_TDATA;
	wire _axis_stream_converters_in_20_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_20_io_dataOut_TDATA;
	wire _axis_stream_converters_in_19_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_19_io_dataOut_TDATA;
	wire _axis_stream_converters_in_18_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_18_io_dataOut_TDATA;
	wire _axis_stream_converters_in_17_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_17_io_dataOut_TDATA;
	wire _axis_stream_converters_in_16_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_16_io_dataOut_TDATA;
	wire _axis_stream_converters_in_15_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_15_io_dataOut_TDATA;
	wire _axis_stream_converters_in_14_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_14_io_dataOut_TDATA;
	wire _axis_stream_converters_in_13_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_13_io_dataOut_TDATA;
	wire _axis_stream_converters_in_12_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_12_io_dataOut_TDATA;
	wire _axis_stream_converters_in_11_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_11_io_dataOut_TDATA;
	wire _axis_stream_converters_in_10_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_10_io_dataOut_TDATA;
	wire _axis_stream_converters_in_9_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_9_io_dataOut_TDATA;
	wire _axis_stream_converters_in_8_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_8_io_dataOut_TDATA;
	wire _axis_stream_converters_in_7_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_7_io_dataOut_TDATA;
	wire _axis_stream_converters_in_6_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_6_io_dataOut_TDATA;
	wire _axis_stream_converters_in_5_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_5_io_dataOut_TDATA;
	wire _axis_stream_converters_in_4_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_4_io_dataOut_TDATA;
	wire _axis_stream_converters_in_3_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_3_io_dataOut_TDATA;
	wire _axis_stream_converters_in_2_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_2_io_dataOut_TDATA;
	wire _axis_stream_converters_in_1_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_1_io_dataOut_TDATA;
	wire _axis_stream_converters_in_0_io_dataOut_TVALID;
	wire [255:0] _axis_stream_converters_in_0_io_dataOut_TDATA;
	wire _axis_stream_converters_out_63_io_dataIn_TREADY;
	wire _axis_stream_converters_out_62_io_dataIn_TREADY;
	wire _axis_stream_converters_out_61_io_dataIn_TREADY;
	wire _axis_stream_converters_out_60_io_dataIn_TREADY;
	wire _axis_stream_converters_out_59_io_dataIn_TREADY;
	wire _axis_stream_converters_out_58_io_dataIn_TREADY;
	wire _axis_stream_converters_out_57_io_dataIn_TREADY;
	wire _axis_stream_converters_out_56_io_dataIn_TREADY;
	wire _axis_stream_converters_out_55_io_dataIn_TREADY;
	wire _axis_stream_converters_out_54_io_dataIn_TREADY;
	wire _axis_stream_converters_out_53_io_dataIn_TREADY;
	wire _axis_stream_converters_out_52_io_dataIn_TREADY;
	wire _axis_stream_converters_out_51_io_dataIn_TREADY;
	wire _axis_stream_converters_out_50_io_dataIn_TREADY;
	wire _axis_stream_converters_out_49_io_dataIn_TREADY;
	wire _axis_stream_converters_out_48_io_dataIn_TREADY;
	wire _axis_stream_converters_out_47_io_dataIn_TREADY;
	wire _axis_stream_converters_out_46_io_dataIn_TREADY;
	wire _axis_stream_converters_out_45_io_dataIn_TREADY;
	wire _axis_stream_converters_out_44_io_dataIn_TREADY;
	wire _axis_stream_converters_out_43_io_dataIn_TREADY;
	wire _axis_stream_converters_out_42_io_dataIn_TREADY;
	wire _axis_stream_converters_out_41_io_dataIn_TREADY;
	wire _axis_stream_converters_out_40_io_dataIn_TREADY;
	wire _axis_stream_converters_out_39_io_dataIn_TREADY;
	wire _axis_stream_converters_out_38_io_dataIn_TREADY;
	wire _axis_stream_converters_out_37_io_dataIn_TREADY;
	wire _axis_stream_converters_out_36_io_dataIn_TREADY;
	wire _axis_stream_converters_out_35_io_dataIn_TREADY;
	wire _axis_stream_converters_out_34_io_dataIn_TREADY;
	wire _axis_stream_converters_out_33_io_dataIn_TREADY;
	wire _axis_stream_converters_out_32_io_dataIn_TREADY;
	wire _axis_stream_converters_out_31_io_dataIn_TREADY;
	wire _axis_stream_converters_out_30_io_dataIn_TREADY;
	wire _axis_stream_converters_out_29_io_dataIn_TREADY;
	wire _axis_stream_converters_out_28_io_dataIn_TREADY;
	wire _axis_stream_converters_out_27_io_dataIn_TREADY;
	wire _axis_stream_converters_out_26_io_dataIn_TREADY;
	wire _axis_stream_converters_out_25_io_dataIn_TREADY;
	wire _axis_stream_converters_out_24_io_dataIn_TREADY;
	wire _axis_stream_converters_out_23_io_dataIn_TREADY;
	wire _axis_stream_converters_out_22_io_dataIn_TREADY;
	wire _axis_stream_converters_out_21_io_dataIn_TREADY;
	wire _axis_stream_converters_out_20_io_dataIn_TREADY;
	wire _axis_stream_converters_out_19_io_dataIn_TREADY;
	wire _axis_stream_converters_out_18_io_dataIn_TREADY;
	wire _axis_stream_converters_out_17_io_dataIn_TREADY;
	wire _axis_stream_converters_out_16_io_dataIn_TREADY;
	wire _axis_stream_converters_out_15_io_dataIn_TREADY;
	wire _axis_stream_converters_out_14_io_dataIn_TREADY;
	wire _axis_stream_converters_out_13_io_dataIn_TREADY;
	wire _axis_stream_converters_out_12_io_dataIn_TREADY;
	wire _axis_stream_converters_out_11_io_dataIn_TREADY;
	wire _axis_stream_converters_out_10_io_dataIn_TREADY;
	wire _axis_stream_converters_out_9_io_dataIn_TREADY;
	wire _axis_stream_converters_out_8_io_dataIn_TREADY;
	wire _axis_stream_converters_out_7_io_dataIn_TREADY;
	wire _axis_stream_converters_out_6_io_dataIn_TREADY;
	wire _axis_stream_converters_out_5_io_dataIn_TREADY;
	wire _axis_stream_converters_out_4_io_dataIn_TREADY;
	wire _axis_stream_converters_out_3_io_dataIn_TREADY;
	wire _axis_stream_converters_out_2_io_dataIn_TREADY;
	wire _axis_stream_converters_out_1_io_dataIn_TREADY;
	wire _axis_stream_converters_out_0_io_dataIn_TREADY;
	wire _module_s_axi_ar_ready;
	wire _module_s_axi_r_valid;
	wire [255:0] _module_s_axi_r_bits_data;
	wire _module_s_axi_aw_ready;
	wire _module_s_axi_w_ready;
	wire _module_s_axi_b_valid;
	wire _vssRvm_0_io_read_address_ready;
	wire _vssRvm_0_io_read_data_valid;
	wire [255:0] _vssRvm_0_io_read_data_bits;
	wire _vssRvm_0_io_write_address_ready;
	wire _vssRvm_0_io_write_data_ready;
	wire _vssRvm_0_axi_ar_valid;
	wire [63:0] _vssRvm_0_axi_ar_bits_addr;
	wire [7:0] _vssRvm_0_axi_ar_bits_len;
	wire _vssRvm_0_axi_r_ready;
	wire _vssRvm_0_axi_aw_valid;
	wire [63:0] _vssRvm_0_axi_aw_bits_addr;
	wire _vssRvm_0_axi_w_valid;
	wire [255:0] _vssRvm_0_axi_w_bits_data;
	wire _vssRvm_0_axi_w_bits_last;
	wire _virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _virtualStealServers_0_io_connNetwork_data_availableTask_ready;
	wire _virtualStealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [255:0] _virtualStealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _virtualStealServers_0_io_read_address_valid;
	wire [63:0] _virtualStealServers_0_io_read_address_bits;
	wire _virtualStealServers_0_io_read_data_ready;
	wire [3:0] _virtualStealServers_0_io_read_burst_len;
	wire _virtualStealServers_0_io_write_address_valid;
	wire [63:0] _virtualStealServers_0_io_write_address_bits;
	wire _virtualStealServers_0_io_write_data_valid;
	wire [255:0] _virtualStealServers_0_io_write_data_bits;
	wire _virtualStealServers_0_io_write_last;
	wire _stealNW_TQ_io_connPE_0_push_ready;
	wire _stealNW_TQ_io_connPE_0_pop_valid;
	wire _stealNW_TQ_io_connPE_1_push_ready;
	wire _stealNW_TQ_io_connPE_1_pop_valid;
	wire _stealNW_TQ_io_connPE_2_push_ready;
	wire _stealNW_TQ_io_connPE_2_pop_valid;
	wire _stealNW_TQ_io_connPE_3_push_ready;
	wire _stealNW_TQ_io_connPE_3_pop_valid;
	wire _stealNW_TQ_io_connPE_4_push_ready;
	wire _stealNW_TQ_io_connPE_4_pop_valid;
	wire _stealNW_TQ_io_connPE_5_push_ready;
	wire _stealNW_TQ_io_connPE_5_pop_valid;
	wire _stealNW_TQ_io_connPE_6_push_ready;
	wire _stealNW_TQ_io_connPE_6_pop_valid;
	wire _stealNW_TQ_io_connPE_7_push_ready;
	wire _stealNW_TQ_io_connPE_7_pop_valid;
	wire _stealNW_TQ_io_connPE_8_push_ready;
	wire _stealNW_TQ_io_connPE_8_pop_valid;
	wire _stealNW_TQ_io_connPE_9_push_ready;
	wire _stealNW_TQ_io_connPE_9_pop_valid;
	wire _stealNW_TQ_io_connPE_10_push_ready;
	wire _stealNW_TQ_io_connPE_10_pop_valid;
	wire _stealNW_TQ_io_connPE_11_push_ready;
	wire _stealNW_TQ_io_connPE_11_pop_valid;
	wire _stealNW_TQ_io_connPE_12_push_ready;
	wire _stealNW_TQ_io_connPE_12_pop_valid;
	wire _stealNW_TQ_io_connPE_13_push_ready;
	wire _stealNW_TQ_io_connPE_13_pop_valid;
	wire _stealNW_TQ_io_connPE_14_push_ready;
	wire _stealNW_TQ_io_connPE_14_pop_valid;
	wire _stealNW_TQ_io_connPE_15_push_ready;
	wire _stealNW_TQ_io_connPE_15_pop_valid;
	wire _stealNW_TQ_io_connPE_16_push_ready;
	wire _stealNW_TQ_io_connPE_16_pop_valid;
	wire _stealNW_TQ_io_connPE_17_push_ready;
	wire _stealNW_TQ_io_connPE_17_pop_valid;
	wire _stealNW_TQ_io_connPE_18_push_ready;
	wire _stealNW_TQ_io_connPE_18_pop_valid;
	wire _stealNW_TQ_io_connPE_19_push_ready;
	wire _stealNW_TQ_io_connPE_19_pop_valid;
	wire _stealNW_TQ_io_connPE_20_push_ready;
	wire _stealNW_TQ_io_connPE_20_pop_valid;
	wire _stealNW_TQ_io_connPE_21_push_ready;
	wire _stealNW_TQ_io_connPE_21_pop_valid;
	wire _stealNW_TQ_io_connPE_22_push_ready;
	wire _stealNW_TQ_io_connPE_22_pop_valid;
	wire _stealNW_TQ_io_connPE_23_push_ready;
	wire _stealNW_TQ_io_connPE_23_pop_valid;
	wire _stealNW_TQ_io_connPE_24_push_ready;
	wire _stealNW_TQ_io_connPE_24_pop_valid;
	wire _stealNW_TQ_io_connPE_25_push_ready;
	wire _stealNW_TQ_io_connPE_25_pop_valid;
	wire _stealNW_TQ_io_connPE_26_push_ready;
	wire _stealNW_TQ_io_connPE_26_pop_valid;
	wire _stealNW_TQ_io_connPE_27_push_ready;
	wire _stealNW_TQ_io_connPE_27_pop_valid;
	wire _stealNW_TQ_io_connPE_28_push_ready;
	wire _stealNW_TQ_io_connPE_28_pop_valid;
	wire _stealNW_TQ_io_connPE_29_push_ready;
	wire _stealNW_TQ_io_connPE_29_pop_valid;
	wire _stealNW_TQ_io_connPE_30_push_ready;
	wire _stealNW_TQ_io_connPE_30_pop_valid;
	wire _stealNW_TQ_io_connPE_31_push_ready;
	wire _stealNW_TQ_io_connPE_31_pop_valid;
	wire _stealNW_TQ_io_connPE_32_push_ready;
	wire _stealNW_TQ_io_connPE_32_pop_valid;
	wire _stealNW_TQ_io_connPE_33_push_ready;
	wire _stealNW_TQ_io_connPE_33_pop_valid;
	wire _stealNW_TQ_io_connPE_34_push_ready;
	wire _stealNW_TQ_io_connPE_34_pop_valid;
	wire _stealNW_TQ_io_connPE_35_push_ready;
	wire _stealNW_TQ_io_connPE_35_pop_valid;
	wire _stealNW_TQ_io_connPE_36_push_ready;
	wire _stealNW_TQ_io_connPE_36_pop_valid;
	wire _stealNW_TQ_io_connPE_37_push_ready;
	wire _stealNW_TQ_io_connPE_37_pop_valid;
	wire _stealNW_TQ_io_connPE_38_push_ready;
	wire _stealNW_TQ_io_connPE_38_pop_valid;
	wire _stealNW_TQ_io_connPE_39_push_ready;
	wire _stealNW_TQ_io_connPE_39_pop_valid;
	wire _stealNW_TQ_io_connPE_40_push_ready;
	wire _stealNW_TQ_io_connPE_40_pop_valid;
	wire _stealNW_TQ_io_connPE_41_push_ready;
	wire _stealNW_TQ_io_connPE_41_pop_valid;
	wire _stealNW_TQ_io_connPE_42_push_ready;
	wire _stealNW_TQ_io_connPE_42_pop_valid;
	wire _stealNW_TQ_io_connPE_43_push_ready;
	wire _stealNW_TQ_io_connPE_43_pop_valid;
	wire _stealNW_TQ_io_connPE_44_push_ready;
	wire _stealNW_TQ_io_connPE_44_pop_valid;
	wire _stealNW_TQ_io_connPE_45_push_ready;
	wire _stealNW_TQ_io_connPE_45_pop_valid;
	wire _stealNW_TQ_io_connPE_46_push_ready;
	wire _stealNW_TQ_io_connPE_46_pop_valid;
	wire _stealNW_TQ_io_connPE_47_push_ready;
	wire _stealNW_TQ_io_connPE_47_pop_valid;
	wire _stealNW_TQ_io_connPE_48_push_ready;
	wire _stealNW_TQ_io_connPE_48_pop_valid;
	wire _stealNW_TQ_io_connPE_49_push_ready;
	wire _stealNW_TQ_io_connPE_49_pop_valid;
	wire _stealNW_TQ_io_connPE_50_push_ready;
	wire _stealNW_TQ_io_connPE_50_pop_valid;
	wire _stealNW_TQ_io_connPE_51_push_ready;
	wire _stealNW_TQ_io_connPE_51_pop_valid;
	wire _stealNW_TQ_io_connPE_52_push_ready;
	wire _stealNW_TQ_io_connPE_52_pop_valid;
	wire _stealNW_TQ_io_connPE_53_push_ready;
	wire _stealNW_TQ_io_connPE_53_pop_valid;
	wire _stealNW_TQ_io_connPE_54_push_ready;
	wire _stealNW_TQ_io_connPE_54_pop_valid;
	wire _stealNW_TQ_io_connPE_55_push_ready;
	wire _stealNW_TQ_io_connPE_55_pop_valid;
	wire _stealNW_TQ_io_connPE_56_push_ready;
	wire _stealNW_TQ_io_connPE_56_pop_valid;
	wire _stealNW_TQ_io_connPE_57_push_ready;
	wire _stealNW_TQ_io_connPE_57_pop_valid;
	wire _stealNW_TQ_io_connPE_58_push_ready;
	wire _stealNW_TQ_io_connPE_58_pop_valid;
	wire _stealNW_TQ_io_connPE_59_push_ready;
	wire _stealNW_TQ_io_connPE_59_pop_valid;
	wire _stealNW_TQ_io_connPE_60_push_ready;
	wire _stealNW_TQ_io_connPE_60_pop_valid;
	wire _stealNW_TQ_io_connPE_61_push_ready;
	wire _stealNW_TQ_io_connPE_61_pop_valid;
	wire _stealNW_TQ_io_connPE_62_push_ready;
	wire _stealNW_TQ_io_connPE_62_pop_valid;
	wire _stealNW_TQ_io_connPE_63_push_ready;
	wire _stealNW_TQ_io_connPE_63_pop_valid;
	wire _stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready;
	wire _stealNW_TQ_io_connVSS_0_data_availableTask_valid;
	wire [255:0] _stealNW_TQ_io_connVSS_0_data_availableTask_bits;
	wire _stealNW_TQ_io_connVSS_0_data_qOutTask_ready;
	wire _stealNW_TQ_io_ntwDataUnitOccupancyVSS_0;
	SchedulerLocalNetwork stealNW_TQ(
		.clock(clock),
		.reset(reset),
		.io_connPE_0_push_ready(_stealNW_TQ_io_connPE_0_push_ready),
		.io_connPE_0_push_valid(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_connPE_0_push_bits(_axis_stream_converters_in_0_io_dataOut_TDATA),
		.io_connPE_0_pop_ready(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_connPE_0_pop_valid(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_connPE_1_push_ready(_stealNW_TQ_io_connPE_1_push_ready),
		.io_connPE_1_push_valid(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_connPE_1_push_bits(_axis_stream_converters_in_1_io_dataOut_TDATA),
		.io_connPE_1_pop_ready(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_connPE_1_pop_valid(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_connPE_2_push_ready(_stealNW_TQ_io_connPE_2_push_ready),
		.io_connPE_2_push_valid(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_connPE_2_push_bits(_axis_stream_converters_in_2_io_dataOut_TDATA),
		.io_connPE_2_pop_ready(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_connPE_2_pop_valid(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_connPE_3_push_ready(_stealNW_TQ_io_connPE_3_push_ready),
		.io_connPE_3_push_valid(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_connPE_3_push_bits(_axis_stream_converters_in_3_io_dataOut_TDATA),
		.io_connPE_3_pop_ready(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_connPE_3_pop_valid(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_connPE_4_push_ready(_stealNW_TQ_io_connPE_4_push_ready),
		.io_connPE_4_push_valid(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_connPE_4_push_bits(_axis_stream_converters_in_4_io_dataOut_TDATA),
		.io_connPE_4_pop_ready(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_connPE_4_pop_valid(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_connPE_5_push_ready(_stealNW_TQ_io_connPE_5_push_ready),
		.io_connPE_5_push_valid(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_connPE_5_push_bits(_axis_stream_converters_in_5_io_dataOut_TDATA),
		.io_connPE_5_pop_ready(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_connPE_5_pop_valid(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_connPE_6_push_ready(_stealNW_TQ_io_connPE_6_push_ready),
		.io_connPE_6_push_valid(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_connPE_6_push_bits(_axis_stream_converters_in_6_io_dataOut_TDATA),
		.io_connPE_6_pop_ready(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_connPE_6_pop_valid(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_connPE_7_push_ready(_stealNW_TQ_io_connPE_7_push_ready),
		.io_connPE_7_push_valid(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_connPE_7_push_bits(_axis_stream_converters_in_7_io_dataOut_TDATA),
		.io_connPE_7_pop_ready(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_connPE_7_pop_valid(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_connPE_8_push_ready(_stealNW_TQ_io_connPE_8_push_ready),
		.io_connPE_8_push_valid(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_connPE_8_push_bits(_axis_stream_converters_in_8_io_dataOut_TDATA),
		.io_connPE_8_pop_ready(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_connPE_8_pop_valid(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_connPE_9_push_ready(_stealNW_TQ_io_connPE_9_push_ready),
		.io_connPE_9_push_valid(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_connPE_9_push_bits(_axis_stream_converters_in_9_io_dataOut_TDATA),
		.io_connPE_9_pop_ready(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_connPE_9_pop_valid(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_connPE_10_push_ready(_stealNW_TQ_io_connPE_10_push_ready),
		.io_connPE_10_push_valid(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_connPE_10_push_bits(_axis_stream_converters_in_10_io_dataOut_TDATA),
		.io_connPE_10_pop_ready(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_connPE_10_pop_valid(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_connPE_11_push_ready(_stealNW_TQ_io_connPE_11_push_ready),
		.io_connPE_11_push_valid(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_connPE_11_push_bits(_axis_stream_converters_in_11_io_dataOut_TDATA),
		.io_connPE_11_pop_ready(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_connPE_11_pop_valid(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_connPE_12_push_ready(_stealNW_TQ_io_connPE_12_push_ready),
		.io_connPE_12_push_valid(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_connPE_12_push_bits(_axis_stream_converters_in_12_io_dataOut_TDATA),
		.io_connPE_12_pop_ready(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_connPE_12_pop_valid(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_connPE_13_push_ready(_stealNW_TQ_io_connPE_13_push_ready),
		.io_connPE_13_push_valid(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_connPE_13_push_bits(_axis_stream_converters_in_13_io_dataOut_TDATA),
		.io_connPE_13_pop_ready(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_connPE_13_pop_valid(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_connPE_14_push_ready(_stealNW_TQ_io_connPE_14_push_ready),
		.io_connPE_14_push_valid(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_connPE_14_push_bits(_axis_stream_converters_in_14_io_dataOut_TDATA),
		.io_connPE_14_pop_ready(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_connPE_14_pop_valid(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_connPE_15_push_ready(_stealNW_TQ_io_connPE_15_push_ready),
		.io_connPE_15_push_valid(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_connPE_15_push_bits(_axis_stream_converters_in_15_io_dataOut_TDATA),
		.io_connPE_15_pop_ready(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_connPE_15_pop_valid(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_connPE_16_push_ready(_stealNW_TQ_io_connPE_16_push_ready),
		.io_connPE_16_push_valid(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_connPE_16_push_bits(_axis_stream_converters_in_16_io_dataOut_TDATA),
		.io_connPE_16_pop_ready(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_connPE_16_pop_valid(_stealNW_TQ_io_connPE_16_pop_valid),
		.io_connPE_17_push_ready(_stealNW_TQ_io_connPE_17_push_ready),
		.io_connPE_17_push_valid(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_connPE_17_push_bits(_axis_stream_converters_in_17_io_dataOut_TDATA),
		.io_connPE_17_pop_ready(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_connPE_17_pop_valid(_stealNW_TQ_io_connPE_17_pop_valid),
		.io_connPE_18_push_ready(_stealNW_TQ_io_connPE_18_push_ready),
		.io_connPE_18_push_valid(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_connPE_18_push_bits(_axis_stream_converters_in_18_io_dataOut_TDATA),
		.io_connPE_18_pop_ready(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_connPE_18_pop_valid(_stealNW_TQ_io_connPE_18_pop_valid),
		.io_connPE_19_push_ready(_stealNW_TQ_io_connPE_19_push_ready),
		.io_connPE_19_push_valid(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_connPE_19_push_bits(_axis_stream_converters_in_19_io_dataOut_TDATA),
		.io_connPE_19_pop_ready(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_connPE_19_pop_valid(_stealNW_TQ_io_connPE_19_pop_valid),
		.io_connPE_20_push_ready(_stealNW_TQ_io_connPE_20_push_ready),
		.io_connPE_20_push_valid(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_connPE_20_push_bits(_axis_stream_converters_in_20_io_dataOut_TDATA),
		.io_connPE_20_pop_ready(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_connPE_20_pop_valid(_stealNW_TQ_io_connPE_20_pop_valid),
		.io_connPE_21_push_ready(_stealNW_TQ_io_connPE_21_push_ready),
		.io_connPE_21_push_valid(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_connPE_21_push_bits(_axis_stream_converters_in_21_io_dataOut_TDATA),
		.io_connPE_21_pop_ready(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_connPE_21_pop_valid(_stealNW_TQ_io_connPE_21_pop_valid),
		.io_connPE_22_push_ready(_stealNW_TQ_io_connPE_22_push_ready),
		.io_connPE_22_push_valid(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_connPE_22_push_bits(_axis_stream_converters_in_22_io_dataOut_TDATA),
		.io_connPE_22_pop_ready(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_connPE_22_pop_valid(_stealNW_TQ_io_connPE_22_pop_valid),
		.io_connPE_23_push_ready(_stealNW_TQ_io_connPE_23_push_ready),
		.io_connPE_23_push_valid(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_connPE_23_push_bits(_axis_stream_converters_in_23_io_dataOut_TDATA),
		.io_connPE_23_pop_ready(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_connPE_23_pop_valid(_stealNW_TQ_io_connPE_23_pop_valid),
		.io_connPE_24_push_ready(_stealNW_TQ_io_connPE_24_push_ready),
		.io_connPE_24_push_valid(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_connPE_24_push_bits(_axis_stream_converters_in_24_io_dataOut_TDATA),
		.io_connPE_24_pop_ready(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_connPE_24_pop_valid(_stealNW_TQ_io_connPE_24_pop_valid),
		.io_connPE_25_push_ready(_stealNW_TQ_io_connPE_25_push_ready),
		.io_connPE_25_push_valid(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_connPE_25_push_bits(_axis_stream_converters_in_25_io_dataOut_TDATA),
		.io_connPE_25_pop_ready(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_connPE_25_pop_valid(_stealNW_TQ_io_connPE_25_pop_valid),
		.io_connPE_26_push_ready(_stealNW_TQ_io_connPE_26_push_ready),
		.io_connPE_26_push_valid(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_connPE_26_push_bits(_axis_stream_converters_in_26_io_dataOut_TDATA),
		.io_connPE_26_pop_ready(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_connPE_26_pop_valid(_stealNW_TQ_io_connPE_26_pop_valid),
		.io_connPE_27_push_ready(_stealNW_TQ_io_connPE_27_push_ready),
		.io_connPE_27_push_valid(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_connPE_27_push_bits(_axis_stream_converters_in_27_io_dataOut_TDATA),
		.io_connPE_27_pop_ready(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_connPE_27_pop_valid(_stealNW_TQ_io_connPE_27_pop_valid),
		.io_connPE_28_push_ready(_stealNW_TQ_io_connPE_28_push_ready),
		.io_connPE_28_push_valid(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_connPE_28_push_bits(_axis_stream_converters_in_28_io_dataOut_TDATA),
		.io_connPE_28_pop_ready(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_connPE_28_pop_valid(_stealNW_TQ_io_connPE_28_pop_valid),
		.io_connPE_29_push_ready(_stealNW_TQ_io_connPE_29_push_ready),
		.io_connPE_29_push_valid(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_connPE_29_push_bits(_axis_stream_converters_in_29_io_dataOut_TDATA),
		.io_connPE_29_pop_ready(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_connPE_29_pop_valid(_stealNW_TQ_io_connPE_29_pop_valid),
		.io_connPE_30_push_ready(_stealNW_TQ_io_connPE_30_push_ready),
		.io_connPE_30_push_valid(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_connPE_30_push_bits(_axis_stream_converters_in_30_io_dataOut_TDATA),
		.io_connPE_30_pop_ready(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_connPE_30_pop_valid(_stealNW_TQ_io_connPE_30_pop_valid),
		.io_connPE_31_push_ready(_stealNW_TQ_io_connPE_31_push_ready),
		.io_connPE_31_push_valid(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_connPE_31_push_bits(_axis_stream_converters_in_31_io_dataOut_TDATA),
		.io_connPE_31_pop_ready(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_connPE_31_pop_valid(_stealNW_TQ_io_connPE_31_pop_valid),
		.io_connPE_32_push_ready(_stealNW_TQ_io_connPE_32_push_ready),
		.io_connPE_32_push_valid(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_connPE_32_push_bits(_axis_stream_converters_in_32_io_dataOut_TDATA),
		.io_connPE_32_pop_ready(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_connPE_32_pop_valid(_stealNW_TQ_io_connPE_32_pop_valid),
		.io_connPE_33_push_ready(_stealNW_TQ_io_connPE_33_push_ready),
		.io_connPE_33_push_valid(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_connPE_33_push_bits(_axis_stream_converters_in_33_io_dataOut_TDATA),
		.io_connPE_33_pop_ready(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_connPE_33_pop_valid(_stealNW_TQ_io_connPE_33_pop_valid),
		.io_connPE_34_push_ready(_stealNW_TQ_io_connPE_34_push_ready),
		.io_connPE_34_push_valid(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_connPE_34_push_bits(_axis_stream_converters_in_34_io_dataOut_TDATA),
		.io_connPE_34_pop_ready(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_connPE_34_pop_valid(_stealNW_TQ_io_connPE_34_pop_valid),
		.io_connPE_35_push_ready(_stealNW_TQ_io_connPE_35_push_ready),
		.io_connPE_35_push_valid(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_connPE_35_push_bits(_axis_stream_converters_in_35_io_dataOut_TDATA),
		.io_connPE_35_pop_ready(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_connPE_35_pop_valid(_stealNW_TQ_io_connPE_35_pop_valid),
		.io_connPE_36_push_ready(_stealNW_TQ_io_connPE_36_push_ready),
		.io_connPE_36_push_valid(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_connPE_36_push_bits(_axis_stream_converters_in_36_io_dataOut_TDATA),
		.io_connPE_36_pop_ready(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_connPE_36_pop_valid(_stealNW_TQ_io_connPE_36_pop_valid),
		.io_connPE_37_push_ready(_stealNW_TQ_io_connPE_37_push_ready),
		.io_connPE_37_push_valid(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_connPE_37_push_bits(_axis_stream_converters_in_37_io_dataOut_TDATA),
		.io_connPE_37_pop_ready(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_connPE_37_pop_valid(_stealNW_TQ_io_connPE_37_pop_valid),
		.io_connPE_38_push_ready(_stealNW_TQ_io_connPE_38_push_ready),
		.io_connPE_38_push_valid(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_connPE_38_push_bits(_axis_stream_converters_in_38_io_dataOut_TDATA),
		.io_connPE_38_pop_ready(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_connPE_38_pop_valid(_stealNW_TQ_io_connPE_38_pop_valid),
		.io_connPE_39_push_ready(_stealNW_TQ_io_connPE_39_push_ready),
		.io_connPE_39_push_valid(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_connPE_39_push_bits(_axis_stream_converters_in_39_io_dataOut_TDATA),
		.io_connPE_39_pop_ready(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_connPE_39_pop_valid(_stealNW_TQ_io_connPE_39_pop_valid),
		.io_connPE_40_push_ready(_stealNW_TQ_io_connPE_40_push_ready),
		.io_connPE_40_push_valid(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_connPE_40_push_bits(_axis_stream_converters_in_40_io_dataOut_TDATA),
		.io_connPE_40_pop_ready(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_connPE_40_pop_valid(_stealNW_TQ_io_connPE_40_pop_valid),
		.io_connPE_41_push_ready(_stealNW_TQ_io_connPE_41_push_ready),
		.io_connPE_41_push_valid(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_connPE_41_push_bits(_axis_stream_converters_in_41_io_dataOut_TDATA),
		.io_connPE_41_pop_ready(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_connPE_41_pop_valid(_stealNW_TQ_io_connPE_41_pop_valid),
		.io_connPE_42_push_ready(_stealNW_TQ_io_connPE_42_push_ready),
		.io_connPE_42_push_valid(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_connPE_42_push_bits(_axis_stream_converters_in_42_io_dataOut_TDATA),
		.io_connPE_42_pop_ready(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_connPE_42_pop_valid(_stealNW_TQ_io_connPE_42_pop_valid),
		.io_connPE_43_push_ready(_stealNW_TQ_io_connPE_43_push_ready),
		.io_connPE_43_push_valid(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_connPE_43_push_bits(_axis_stream_converters_in_43_io_dataOut_TDATA),
		.io_connPE_43_pop_ready(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_connPE_43_pop_valid(_stealNW_TQ_io_connPE_43_pop_valid),
		.io_connPE_44_push_ready(_stealNW_TQ_io_connPE_44_push_ready),
		.io_connPE_44_push_valid(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_connPE_44_push_bits(_axis_stream_converters_in_44_io_dataOut_TDATA),
		.io_connPE_44_pop_ready(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_connPE_44_pop_valid(_stealNW_TQ_io_connPE_44_pop_valid),
		.io_connPE_45_push_ready(_stealNW_TQ_io_connPE_45_push_ready),
		.io_connPE_45_push_valid(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_connPE_45_push_bits(_axis_stream_converters_in_45_io_dataOut_TDATA),
		.io_connPE_45_pop_ready(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_connPE_45_pop_valid(_stealNW_TQ_io_connPE_45_pop_valid),
		.io_connPE_46_push_ready(_stealNW_TQ_io_connPE_46_push_ready),
		.io_connPE_46_push_valid(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_connPE_46_push_bits(_axis_stream_converters_in_46_io_dataOut_TDATA),
		.io_connPE_46_pop_ready(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_connPE_46_pop_valid(_stealNW_TQ_io_connPE_46_pop_valid),
		.io_connPE_47_push_ready(_stealNW_TQ_io_connPE_47_push_ready),
		.io_connPE_47_push_valid(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_connPE_47_push_bits(_axis_stream_converters_in_47_io_dataOut_TDATA),
		.io_connPE_47_pop_ready(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_connPE_47_pop_valid(_stealNW_TQ_io_connPE_47_pop_valid),
		.io_connPE_48_push_ready(_stealNW_TQ_io_connPE_48_push_ready),
		.io_connPE_48_push_valid(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_connPE_48_push_bits(_axis_stream_converters_in_48_io_dataOut_TDATA),
		.io_connPE_48_pop_ready(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_connPE_48_pop_valid(_stealNW_TQ_io_connPE_48_pop_valid),
		.io_connPE_49_push_ready(_stealNW_TQ_io_connPE_49_push_ready),
		.io_connPE_49_push_valid(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_connPE_49_push_bits(_axis_stream_converters_in_49_io_dataOut_TDATA),
		.io_connPE_49_pop_ready(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_connPE_49_pop_valid(_stealNW_TQ_io_connPE_49_pop_valid),
		.io_connPE_50_push_ready(_stealNW_TQ_io_connPE_50_push_ready),
		.io_connPE_50_push_valid(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_connPE_50_push_bits(_axis_stream_converters_in_50_io_dataOut_TDATA),
		.io_connPE_50_pop_ready(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_connPE_50_pop_valid(_stealNW_TQ_io_connPE_50_pop_valid),
		.io_connPE_51_push_ready(_stealNW_TQ_io_connPE_51_push_ready),
		.io_connPE_51_push_valid(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_connPE_51_push_bits(_axis_stream_converters_in_51_io_dataOut_TDATA),
		.io_connPE_51_pop_ready(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_connPE_51_pop_valid(_stealNW_TQ_io_connPE_51_pop_valid),
		.io_connPE_52_push_ready(_stealNW_TQ_io_connPE_52_push_ready),
		.io_connPE_52_push_valid(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_connPE_52_push_bits(_axis_stream_converters_in_52_io_dataOut_TDATA),
		.io_connPE_52_pop_ready(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_connPE_52_pop_valid(_stealNW_TQ_io_connPE_52_pop_valid),
		.io_connPE_53_push_ready(_stealNW_TQ_io_connPE_53_push_ready),
		.io_connPE_53_push_valid(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_connPE_53_push_bits(_axis_stream_converters_in_53_io_dataOut_TDATA),
		.io_connPE_53_pop_ready(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_connPE_53_pop_valid(_stealNW_TQ_io_connPE_53_pop_valid),
		.io_connPE_54_push_ready(_stealNW_TQ_io_connPE_54_push_ready),
		.io_connPE_54_push_valid(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_connPE_54_push_bits(_axis_stream_converters_in_54_io_dataOut_TDATA),
		.io_connPE_54_pop_ready(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_connPE_54_pop_valid(_stealNW_TQ_io_connPE_54_pop_valid),
		.io_connPE_55_push_ready(_stealNW_TQ_io_connPE_55_push_ready),
		.io_connPE_55_push_valid(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_connPE_55_push_bits(_axis_stream_converters_in_55_io_dataOut_TDATA),
		.io_connPE_55_pop_ready(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_connPE_55_pop_valid(_stealNW_TQ_io_connPE_55_pop_valid),
		.io_connPE_56_push_ready(_stealNW_TQ_io_connPE_56_push_ready),
		.io_connPE_56_push_valid(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_connPE_56_push_bits(_axis_stream_converters_in_56_io_dataOut_TDATA),
		.io_connPE_56_pop_ready(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_connPE_56_pop_valid(_stealNW_TQ_io_connPE_56_pop_valid),
		.io_connPE_57_push_ready(_stealNW_TQ_io_connPE_57_push_ready),
		.io_connPE_57_push_valid(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_connPE_57_push_bits(_axis_stream_converters_in_57_io_dataOut_TDATA),
		.io_connPE_57_pop_ready(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_connPE_57_pop_valid(_stealNW_TQ_io_connPE_57_pop_valid),
		.io_connPE_58_push_ready(_stealNW_TQ_io_connPE_58_push_ready),
		.io_connPE_58_push_valid(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_connPE_58_push_bits(_axis_stream_converters_in_58_io_dataOut_TDATA),
		.io_connPE_58_pop_ready(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_connPE_58_pop_valid(_stealNW_TQ_io_connPE_58_pop_valid),
		.io_connPE_59_push_ready(_stealNW_TQ_io_connPE_59_push_ready),
		.io_connPE_59_push_valid(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_connPE_59_push_bits(_axis_stream_converters_in_59_io_dataOut_TDATA),
		.io_connPE_59_pop_ready(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_connPE_59_pop_valid(_stealNW_TQ_io_connPE_59_pop_valid),
		.io_connPE_60_push_ready(_stealNW_TQ_io_connPE_60_push_ready),
		.io_connPE_60_push_valid(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_connPE_60_push_bits(_axis_stream_converters_in_60_io_dataOut_TDATA),
		.io_connPE_60_pop_ready(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_connPE_60_pop_valid(_stealNW_TQ_io_connPE_60_pop_valid),
		.io_connPE_61_push_ready(_stealNW_TQ_io_connPE_61_push_ready),
		.io_connPE_61_push_valid(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_connPE_61_push_bits(_axis_stream_converters_in_61_io_dataOut_TDATA),
		.io_connPE_61_pop_ready(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_connPE_61_pop_valid(_stealNW_TQ_io_connPE_61_pop_valid),
		.io_connPE_62_push_ready(_stealNW_TQ_io_connPE_62_push_ready),
		.io_connPE_62_push_valid(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_connPE_62_push_bits(_axis_stream_converters_in_62_io_dataOut_TDATA),
		.io_connPE_62_pop_ready(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_connPE_62_pop_valid(_stealNW_TQ_io_connPE_62_pop_valid),
		.io_connPE_63_push_ready(_stealNW_TQ_io_connPE_63_push_ready),
		.io_connPE_63_push_valid(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_connPE_63_push_bits(_axis_stream_converters_in_63_io_dataOut_TDATA),
		.io_connPE_63_pop_ready(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_connPE_63_pop_valid(_stealNW_TQ_io_connPE_63_pop_valid),
		.io_connVSS_0_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connVSS_0_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connVSS_0_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connVSS_0_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connVSS_0_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connVSS_0_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connVSS_0_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connVSS_0_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerServer virtualStealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connNetwork_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vss_0_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vss_0_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vss_0_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vss_0_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vss_0_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vss_0_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vss_0_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vss_0_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vss_0_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vss_0_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vss_0_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vss_0_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vss_0_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vss_0_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vss_0_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vss_0_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vss_0_b_bits_resp),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_read_burst_len(_virtualStealServers_0_io_read_burst_len),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_write_last(_virtualStealServers_0_io_write_last),
		.io_ntwDataUnitOccupancy(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
	);
	RVtoAXIBridge vssRvm_0(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_writeBurst_last(_virtualStealServers_0_io_write_last),
		.io_readBurst_len(_virtualStealServers_0_io_read_burst_len),
		.axi_ar_ready(_module_s_axi_ar_ready),
		.axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.axi_r_ready(_vssRvm_0_axi_r_ready),
		.axi_r_valid(_module_s_axi_r_valid),
		.axi_r_bits_data(_module_s_axi_r_bits_data),
		.axi_aw_ready(_module_s_axi_aw_ready),
		.axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.axi_w_ready(_module_s_axi_w_ready),
		.axi_w_valid(_vssRvm_0_axi_w_valid),
		.axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.axi_b_valid(_module_s_axi_b_valid)
	);
	AxiWriteBuffer module_0(
		.clock(clock),
		.reset(reset),
		.s_axi_ar_ready(_module_s_axi_ar_ready),
		.s_axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.s_axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.s_axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.s_axi_r_ready(_vssRvm_0_axi_r_ready),
		.s_axi_r_valid(_module_s_axi_r_valid),
		.s_axi_r_bits_data(_module_s_axi_r_bits_data),
		.s_axi_aw_ready(_module_s_axi_aw_ready),
		.s_axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.s_axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.s_axi_w_ready(_module_s_axi_w_ready),
		.s_axi_w_valid(_vssRvm_0_axi_w_valid),
		.s_axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.s_axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.s_axi_b_valid(_module_s_axi_b_valid),
		.m_axi_ar_ready(io_internal_vss_axi_full_0_ar_ready),
		.m_axi_ar_valid(io_internal_vss_axi_full_0_ar_valid),
		.m_axi_ar_bits_addr(io_internal_vss_axi_full_0_ar_bits_addr),
		.m_axi_ar_bits_len(io_internal_vss_axi_full_0_ar_bits_len),
		.m_axi_ar_bits_size(io_internal_vss_axi_full_0_ar_bits_size),
		.m_axi_ar_bits_burst(io_internal_vss_axi_full_0_ar_bits_burst),
		.m_axi_ar_bits_lock(io_internal_vss_axi_full_0_ar_bits_lock),
		.m_axi_ar_bits_cache(io_internal_vss_axi_full_0_ar_bits_cache),
		.m_axi_ar_bits_prot(io_internal_vss_axi_full_0_ar_bits_prot),
		.m_axi_ar_bits_qos(io_internal_vss_axi_full_0_ar_bits_qos),
		.m_axi_ar_bits_region(io_internal_vss_axi_full_0_ar_bits_region),
		.m_axi_r_ready(io_internal_vss_axi_full_0_r_ready),
		.m_axi_r_valid(io_internal_vss_axi_full_0_r_valid),
		.m_axi_r_bits_data(io_internal_vss_axi_full_0_r_bits_data),
		.m_axi_aw_ready(io_internal_vss_axi_full_0_aw_ready),
		.m_axi_aw_valid(io_internal_vss_axi_full_0_aw_valid),
		.m_axi_aw_bits_addr(io_internal_vss_axi_full_0_aw_bits_addr),
		.m_axi_aw_bits_len(io_internal_vss_axi_full_0_aw_bits_len),
		.m_axi_aw_bits_size(io_internal_vss_axi_full_0_aw_bits_size),
		.m_axi_aw_bits_burst(io_internal_vss_axi_full_0_aw_bits_burst),
		.m_axi_aw_bits_lock(io_internal_vss_axi_full_0_aw_bits_lock),
		.m_axi_aw_bits_cache(io_internal_vss_axi_full_0_aw_bits_cache),
		.m_axi_aw_bits_prot(io_internal_vss_axi_full_0_aw_bits_prot),
		.m_axi_aw_bits_qos(io_internal_vss_axi_full_0_aw_bits_qos),
		.m_axi_aw_bits_region(io_internal_vss_axi_full_0_aw_bits_region),
		.m_axi_w_ready(io_internal_vss_axi_full_0_w_ready),
		.m_axi_w_valid(io_internal_vss_axi_full_0_w_valid),
		.m_axi_w_bits_data(io_internal_vss_axi_full_0_w_bits_data),
		.m_axi_w_bits_last(io_internal_vss_axi_full_0_w_bits_last),
		.m_axi_b_valid(io_internal_vss_axi_full_0_b_valid)
	);
	AxisDataWidthConverter axis_stream_converters_out_0(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_0_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_0_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_1(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_1_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_1_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_2(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_2_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_2_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_3(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_3_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_3_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_4(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_4_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_4_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_5(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_5_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_5_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_6(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_6_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_6_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_7(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_7_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_7_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_8(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_8_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_8_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_9(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_9_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_9_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_10(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_10_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_10_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_11(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_11_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_11_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_12(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_12_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_12_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_13(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_13_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_13_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_14(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_14_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_14_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_15(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_15_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_15_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_16(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_16_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_16_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_16_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_17(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_17_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_17_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_17_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_18(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_18_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_18_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_18_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_19(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_19_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_19_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_19_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_20(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_20_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_20_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_20_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_21(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_21_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_21_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_21_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_22(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_22_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_22_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_22_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_23(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_23_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_23_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_23_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_24(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_24_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_24_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_24_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_25(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_25_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_25_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_25_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_26(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_26_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_26_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_26_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_27(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_27_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_27_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_27_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_28(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_28_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_28_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_28_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_29(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_29_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_29_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_29_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_30(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_30_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_30_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_30_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_31(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_31_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_31_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_31_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_32(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_32_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_32_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_32_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_33(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_33_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_33_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_33_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_34(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_34_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_34_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_34_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_35(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_35_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_35_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_35_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_36(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_36_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_36_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_36_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_37(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_37_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_37_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_37_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_38(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_38_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_38_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_38_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_39(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_39_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_39_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_39_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_40(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_40_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_40_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_40_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_41(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_41_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_41_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_41_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_42(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_42_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_42_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_42_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_43(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_43_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_43_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_43_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_44(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_44_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_44_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_44_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_45(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_45_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_45_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_45_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_46(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_46_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_46_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_46_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_47(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_47_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_47_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_47_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_48(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_48_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_48_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_48_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_49(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_49_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_49_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_49_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_50(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_50_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_50_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_50_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_51(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_51_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_51_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_51_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_52(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_52_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_52_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_52_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_53(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_53_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_53_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_53_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_54(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_54_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_54_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_54_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_55(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_55_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_55_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_55_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_56(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_56_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_56_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_56_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_57(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_57_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_57_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_57_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_58(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_58_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_58_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_58_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_59(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_59_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_59_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_59_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_60(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_60_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_60_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_60_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_61(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_61_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_61_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_61_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_62(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_62_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_62_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_62_TVALID)
	);
	AxisDataWidthConverter axis_stream_converters_out_63(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_63_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_63_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_63_TVALID)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_0(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_0_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_0_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_0_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_0_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_0_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_1(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_1_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_1_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_1_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_1_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_1_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_2(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_2_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_2_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_2_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_2_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_2_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_3(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_3_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_3_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_3_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_3_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_3_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_4(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_4_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_4_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_4_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_4_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_4_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_5(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_5_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_5_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_5_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_5_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_5_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_6(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_6_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_6_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_6_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_6_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_6_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_7(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_7_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_7_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_7_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_7_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_7_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_8(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_8_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_8_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_8_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_8_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_8_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_9(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_9_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_9_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_9_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_9_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_9_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_10(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_10_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_10_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_10_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_10_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_10_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_11(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_11_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_11_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_11_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_11_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_11_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_12(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_12_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_12_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_12_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_12_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_12_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_13(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_13_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_13_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_13_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_13_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_13_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_14(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_14_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_14_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_14_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_14_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_14_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_15(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_15_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_15_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_15_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_15_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_15_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_16(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_16_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_16_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_16_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_16_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_16_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_17(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_17_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_17_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_17_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_17_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_17_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_18(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_18_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_18_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_18_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_18_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_18_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_19(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_19_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_19_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_19_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_19_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_19_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_20(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_20_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_20_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_20_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_20_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_20_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_21(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_21_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_21_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_21_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_21_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_21_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_22(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_22_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_22_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_22_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_22_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_22_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_23(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_23_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_23_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_23_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_23_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_23_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_24(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_24_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_24_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_24_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_24_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_24_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_25(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_25_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_25_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_25_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_25_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_25_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_26(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_26_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_26_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_26_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_26_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_26_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_27(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_27_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_27_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_27_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_27_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_27_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_28(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_28_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_28_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_28_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_28_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_28_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_29(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_29_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_29_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_29_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_29_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_29_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_30(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_30_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_30_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_30_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_30_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_30_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_31(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_31_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_31_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_31_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_31_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_31_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_32(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_32_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_32_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_32_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_32_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_32_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_33(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_33_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_33_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_33_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_33_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_33_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_34(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_34_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_34_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_34_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_34_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_34_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_35(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_35_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_35_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_35_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_35_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_35_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_36(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_36_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_36_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_36_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_36_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_36_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_37(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_37_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_37_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_37_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_37_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_37_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_38(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_38_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_38_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_38_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_38_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_38_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_39(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_39_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_39_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_39_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_39_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_39_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_40(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_40_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_40_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_40_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_40_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_40_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_41(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_41_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_41_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_41_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_41_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_41_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_42(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_42_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_42_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_42_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_42_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_42_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_43(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_43_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_43_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_43_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_43_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_43_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_44(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_44_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_44_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_44_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_44_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_44_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_45(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_45_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_45_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_45_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_45_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_45_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_46(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_46_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_46_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_46_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_46_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_46_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_47(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_47_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_47_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_47_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_47_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_47_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_48(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_48_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_48_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_48_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_48_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_48_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_49(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_49_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_49_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_49_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_49_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_49_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_50(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_50_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_50_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_50_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_50_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_50_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_51(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_51_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_51_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_51_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_51_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_51_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_52(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_52_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_52_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_52_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_52_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_52_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_53(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_53_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_53_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_53_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_53_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_53_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_54(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_54_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_54_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_54_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_54_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_54_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_55(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_55_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_55_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_55_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_55_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_55_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_56(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_56_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_56_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_56_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_56_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_56_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_57(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_57_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_57_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_57_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_57_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_57_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_58(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_58_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_58_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_58_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_58_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_58_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_59(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_59_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_59_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_59_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_59_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_59_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_60(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_60_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_60_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_60_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_60_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_60_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_61(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_61_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_61_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_61_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_61_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_61_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_62(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_62_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_62_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_62_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_62_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_62_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_64 axis_stream_converters_in_63(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_export_taskIn_63_TREADY),
		.io_dataIn_TVALID(io_export_taskIn_63_TVALID),
		.io_dataIn_TDATA(io_export_taskIn_63_TDATA),
		.io_dataOut_TREADY(_stealNW_TQ_io_connPE_63_push_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_63_io_dataOut_TDATA)
	);
endmodule
module SchedulerNetworkDataUnit_65 (
	clock,
	reset,
	io_taskIn,
	io_taskOut,
	io_validIn,
	io_validOut,
	io_connSS_availableTask_ready,
	io_connSS_availableTask_valid,
	io_connSS_availableTask_bits,
	io_connSS_qOutTask_ready,
	io_connSS_qOutTask_valid,
	io_connSS_qOutTask_bits,
	io_occupied
);
	input clock;
	input reset;
	input [127:0] io_taskIn;
	output wire [127:0] io_taskOut;
	input io_validIn;
	output wire io_validOut;
	input io_connSS_availableTask_ready;
	output wire io_connSS_availableTask_valid;
	output wire [127:0] io_connSS_availableTask_bits;
	output wire io_connSS_qOutTask_ready;
	input io_connSS_qOutTask_valid;
	input [127:0] io_connSS_qOutTask_bits;
	output wire io_occupied;
	reg [127:0] taskReg;
	reg validReg;
	wire io_connSS_availableTask_valid_0 = io_connSS_availableTask_ready & io_validIn;
	wire _GEN = io_connSS_qOutTask_valid & ~io_validIn;
	always @(posedge clock)
		if (reset) begin
			taskReg <= 128'h00000000000000000000000000000000;
			validReg <= 1'h0;
		end
		else begin
			taskReg <= (io_connSS_availableTask_valid_0 ? 128'h00000000000000000000000000000000 : (_GEN ? io_connSS_qOutTask_bits : (io_validIn ? io_taskIn : 128'h00000000000000000000000000000000)));
			validReg <= ~io_connSS_availableTask_valid_0 & (_GEN | io_validIn);
		end
	assign io_taskOut = taskReg;
	assign io_validOut = validReg;
	assign io_connSS_availableTask_valid = io_connSS_availableTask_valid_0;
	assign io_connSS_availableTask_bits = (io_connSS_availableTask_valid_0 ? io_taskIn : 128'h00000000000000000000000000000000);
	assign io_connSS_qOutTask_ready = ~io_connSS_availableTask_valid_0 & _GEN;
	assign io_occupied = validReg;
endmodule
module SchedulerNetwork_1 (
	clock,
	reset,
	io_connSS_0_ctrl_serveStealReq_valid,
	io_connSS_0_ctrl_serveStealReq_ready,
	io_connSS_0_data_availableTask_ready,
	io_connSS_0_data_availableTask_valid,
	io_connSS_0_data_availableTask_bits,
	io_connSS_0_data_qOutTask_ready,
	io_connSS_0_data_qOutTask_valid,
	io_connSS_0_data_qOutTask_bits,
	io_connSS_1_ctrl_serveStealReq_valid,
	io_connSS_1_ctrl_serveStealReq_ready,
	io_connSS_1_data_qOutTask_ready,
	io_connSS_1_data_qOutTask_valid,
	io_connSS_1_data_qOutTask_bits,
	io_connSS_2_ctrl_serveStealReq_valid,
	io_connSS_2_ctrl_serveStealReq_ready,
	io_connSS_2_data_qOutTask_ready,
	io_connSS_2_data_qOutTask_valid,
	io_connSS_2_data_qOutTask_bits,
	io_connSS_3_ctrl_serveStealReq_valid,
	io_connSS_3_ctrl_serveStealReq_ready,
	io_connSS_3_data_qOutTask_ready,
	io_connSS_3_data_qOutTask_valid,
	io_connSS_3_data_qOutTask_bits,
	io_connSS_4_ctrl_serveStealReq_valid,
	io_connSS_4_ctrl_serveStealReq_ready,
	io_connSS_4_data_qOutTask_ready,
	io_connSS_4_data_qOutTask_valid,
	io_connSS_4_data_qOutTask_bits,
	io_connSS_5_ctrl_serveStealReq_valid,
	io_connSS_5_ctrl_serveStealReq_ready,
	io_connSS_5_data_qOutTask_ready,
	io_connSS_5_data_qOutTask_valid,
	io_connSS_5_data_qOutTask_bits,
	io_connSS_6_ctrl_serveStealReq_valid,
	io_connSS_6_ctrl_serveStealReq_ready,
	io_connSS_6_data_qOutTask_ready,
	io_connSS_6_data_qOutTask_valid,
	io_connSS_6_data_qOutTask_bits,
	io_connSS_7_ctrl_serveStealReq_valid,
	io_connSS_7_ctrl_serveStealReq_ready,
	io_connSS_7_data_qOutTask_ready,
	io_connSS_7_data_qOutTask_valid,
	io_connSS_7_data_qOutTask_bits,
	io_connSS_8_ctrl_serveStealReq_valid,
	io_connSS_8_ctrl_serveStealReq_ready,
	io_connSS_8_data_qOutTask_ready,
	io_connSS_8_data_qOutTask_valid,
	io_connSS_8_data_qOutTask_bits,
	io_connSS_9_ctrl_serveStealReq_valid,
	io_connSS_9_ctrl_serveStealReq_ready,
	io_connSS_9_data_qOutTask_ready,
	io_connSS_9_data_qOutTask_valid,
	io_connSS_9_data_qOutTask_bits,
	io_connSS_10_ctrl_serveStealReq_valid,
	io_connSS_10_ctrl_serveStealReq_ready,
	io_connSS_10_data_qOutTask_ready,
	io_connSS_10_data_qOutTask_valid,
	io_connSS_10_data_qOutTask_bits,
	io_connSS_11_ctrl_serveStealReq_valid,
	io_connSS_11_ctrl_serveStealReq_ready,
	io_connSS_11_data_qOutTask_ready,
	io_connSS_11_data_qOutTask_valid,
	io_connSS_11_data_qOutTask_bits,
	io_connSS_12_ctrl_serveStealReq_valid,
	io_connSS_12_ctrl_serveStealReq_ready,
	io_connSS_12_data_qOutTask_ready,
	io_connSS_12_data_qOutTask_valid,
	io_connSS_12_data_qOutTask_bits,
	io_connSS_13_ctrl_serveStealReq_valid,
	io_connSS_13_ctrl_serveStealReq_ready,
	io_connSS_13_data_qOutTask_ready,
	io_connSS_13_data_qOutTask_valid,
	io_connSS_13_data_qOutTask_bits,
	io_connSS_14_ctrl_serveStealReq_valid,
	io_connSS_14_ctrl_serveStealReq_ready,
	io_connSS_14_data_qOutTask_ready,
	io_connSS_14_data_qOutTask_valid,
	io_connSS_14_data_qOutTask_bits,
	io_connSS_15_ctrl_serveStealReq_valid,
	io_connSS_15_ctrl_serveStealReq_ready,
	io_connSS_15_data_qOutTask_ready,
	io_connSS_15_data_qOutTask_valid,
	io_connSS_15_data_qOutTask_bits,
	io_connSS_16_ctrl_serveStealReq_valid,
	io_connSS_16_ctrl_serveStealReq_ready,
	io_connSS_16_data_qOutTask_ready,
	io_connSS_16_data_qOutTask_valid,
	io_connSS_16_data_qOutTask_bits,
	io_connSS_17_ctrl_serveStealReq_valid,
	io_connSS_17_ctrl_serveStealReq_ready,
	io_connSS_17_ctrl_stealReq_valid,
	io_connSS_17_ctrl_stealReq_ready,
	io_connSS_17_data_availableTask_ready,
	io_connSS_17_data_availableTask_valid,
	io_connSS_17_data_availableTask_bits,
	io_connSS_17_data_qOutTask_ready,
	io_connSS_17_data_qOutTask_valid,
	io_connSS_17_data_qOutTask_bits,
	io_connSS_18_ctrl_serveStealReq_valid,
	io_connSS_18_ctrl_serveStealReq_ready,
	io_connSS_18_ctrl_stealReq_valid,
	io_connSS_18_ctrl_stealReq_ready,
	io_connSS_18_data_availableTask_ready,
	io_connSS_18_data_availableTask_valid,
	io_connSS_18_data_availableTask_bits,
	io_connSS_18_data_qOutTask_ready,
	io_connSS_18_data_qOutTask_valid,
	io_connSS_18_data_qOutTask_bits,
	io_connSS_19_ctrl_serveStealReq_valid,
	io_connSS_19_ctrl_serveStealReq_ready,
	io_connSS_19_ctrl_stealReq_valid,
	io_connSS_19_ctrl_stealReq_ready,
	io_connSS_19_data_availableTask_ready,
	io_connSS_19_data_availableTask_valid,
	io_connSS_19_data_availableTask_bits,
	io_connSS_19_data_qOutTask_ready,
	io_connSS_19_data_qOutTask_valid,
	io_connSS_19_data_qOutTask_bits,
	io_connSS_20_ctrl_serveStealReq_valid,
	io_connSS_20_ctrl_serveStealReq_ready,
	io_connSS_20_ctrl_stealReq_valid,
	io_connSS_20_ctrl_stealReq_ready,
	io_connSS_20_data_availableTask_ready,
	io_connSS_20_data_availableTask_valid,
	io_connSS_20_data_availableTask_bits,
	io_connSS_20_data_qOutTask_ready,
	io_connSS_20_data_qOutTask_valid,
	io_connSS_20_data_qOutTask_bits,
	io_connSS_21_ctrl_serveStealReq_valid,
	io_connSS_21_ctrl_serveStealReq_ready,
	io_connSS_21_ctrl_stealReq_valid,
	io_connSS_21_ctrl_stealReq_ready,
	io_connSS_21_data_availableTask_ready,
	io_connSS_21_data_availableTask_valid,
	io_connSS_21_data_availableTask_bits,
	io_connSS_21_data_qOutTask_ready,
	io_connSS_21_data_qOutTask_valid,
	io_connSS_21_data_qOutTask_bits,
	io_connSS_22_ctrl_serveStealReq_valid,
	io_connSS_22_ctrl_serveStealReq_ready,
	io_connSS_22_ctrl_stealReq_valid,
	io_connSS_22_ctrl_stealReq_ready,
	io_connSS_22_data_availableTask_ready,
	io_connSS_22_data_availableTask_valid,
	io_connSS_22_data_availableTask_bits,
	io_connSS_22_data_qOutTask_ready,
	io_connSS_22_data_qOutTask_valid,
	io_connSS_22_data_qOutTask_bits,
	io_connSS_23_ctrl_serveStealReq_valid,
	io_connSS_23_ctrl_serveStealReq_ready,
	io_connSS_23_ctrl_stealReq_valid,
	io_connSS_23_ctrl_stealReq_ready,
	io_connSS_23_data_availableTask_ready,
	io_connSS_23_data_availableTask_valid,
	io_connSS_23_data_availableTask_bits,
	io_connSS_23_data_qOutTask_ready,
	io_connSS_23_data_qOutTask_valid,
	io_connSS_23_data_qOutTask_bits,
	io_connSS_24_ctrl_serveStealReq_valid,
	io_connSS_24_ctrl_serveStealReq_ready,
	io_connSS_24_ctrl_stealReq_valid,
	io_connSS_24_ctrl_stealReq_ready,
	io_connSS_24_data_availableTask_ready,
	io_connSS_24_data_availableTask_valid,
	io_connSS_24_data_availableTask_bits,
	io_connSS_24_data_qOutTask_ready,
	io_connSS_24_data_qOutTask_valid,
	io_connSS_24_data_qOutTask_bits,
	io_connSS_25_ctrl_serveStealReq_valid,
	io_connSS_25_ctrl_serveStealReq_ready,
	io_connSS_25_ctrl_stealReq_valid,
	io_connSS_25_ctrl_stealReq_ready,
	io_connSS_25_data_availableTask_ready,
	io_connSS_25_data_availableTask_valid,
	io_connSS_25_data_availableTask_bits,
	io_connSS_25_data_qOutTask_ready,
	io_connSS_25_data_qOutTask_valid,
	io_connSS_25_data_qOutTask_bits,
	io_connSS_26_ctrl_serveStealReq_valid,
	io_connSS_26_ctrl_serveStealReq_ready,
	io_connSS_26_ctrl_stealReq_valid,
	io_connSS_26_ctrl_stealReq_ready,
	io_connSS_26_data_availableTask_ready,
	io_connSS_26_data_availableTask_valid,
	io_connSS_26_data_availableTask_bits,
	io_connSS_26_data_qOutTask_ready,
	io_connSS_26_data_qOutTask_valid,
	io_connSS_26_data_qOutTask_bits,
	io_connSS_27_ctrl_serveStealReq_valid,
	io_connSS_27_ctrl_serveStealReq_ready,
	io_connSS_27_ctrl_stealReq_valid,
	io_connSS_27_ctrl_stealReq_ready,
	io_connSS_27_data_availableTask_ready,
	io_connSS_27_data_availableTask_valid,
	io_connSS_27_data_availableTask_bits,
	io_connSS_27_data_qOutTask_ready,
	io_connSS_27_data_qOutTask_valid,
	io_connSS_27_data_qOutTask_bits,
	io_connSS_28_ctrl_serveStealReq_valid,
	io_connSS_28_ctrl_serveStealReq_ready,
	io_connSS_28_ctrl_stealReq_valid,
	io_connSS_28_ctrl_stealReq_ready,
	io_connSS_28_data_availableTask_ready,
	io_connSS_28_data_availableTask_valid,
	io_connSS_28_data_availableTask_bits,
	io_connSS_28_data_qOutTask_ready,
	io_connSS_28_data_qOutTask_valid,
	io_connSS_28_data_qOutTask_bits,
	io_connSS_29_ctrl_serveStealReq_valid,
	io_connSS_29_ctrl_serveStealReq_ready,
	io_connSS_29_ctrl_stealReq_valid,
	io_connSS_29_ctrl_stealReq_ready,
	io_connSS_29_data_availableTask_ready,
	io_connSS_29_data_availableTask_valid,
	io_connSS_29_data_availableTask_bits,
	io_connSS_29_data_qOutTask_ready,
	io_connSS_29_data_qOutTask_valid,
	io_connSS_29_data_qOutTask_bits,
	io_connSS_30_ctrl_serveStealReq_valid,
	io_connSS_30_ctrl_serveStealReq_ready,
	io_connSS_30_ctrl_stealReq_valid,
	io_connSS_30_ctrl_stealReq_ready,
	io_connSS_30_data_availableTask_ready,
	io_connSS_30_data_availableTask_valid,
	io_connSS_30_data_availableTask_bits,
	io_connSS_30_data_qOutTask_ready,
	io_connSS_30_data_qOutTask_valid,
	io_connSS_30_data_qOutTask_bits,
	io_connSS_31_ctrl_serveStealReq_valid,
	io_connSS_31_ctrl_serveStealReq_ready,
	io_connSS_31_ctrl_stealReq_valid,
	io_connSS_31_ctrl_stealReq_ready,
	io_connSS_31_data_availableTask_ready,
	io_connSS_31_data_availableTask_valid,
	io_connSS_31_data_availableTask_bits,
	io_connSS_31_data_qOutTask_ready,
	io_connSS_31_data_qOutTask_valid,
	io_connSS_31_data_qOutTask_bits,
	io_connSS_32_ctrl_serveStealReq_valid,
	io_connSS_32_ctrl_serveStealReq_ready,
	io_connSS_32_ctrl_stealReq_valid,
	io_connSS_32_ctrl_stealReq_ready,
	io_connSS_32_data_availableTask_ready,
	io_connSS_32_data_availableTask_valid,
	io_connSS_32_data_availableTask_bits,
	io_connSS_32_data_qOutTask_ready,
	io_connSS_32_data_qOutTask_valid,
	io_connSS_32_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0
);
	input clock;
	input reset;
	input io_connSS_0_ctrl_serveStealReq_valid;
	output wire io_connSS_0_ctrl_serveStealReq_ready;
	input io_connSS_0_data_availableTask_ready;
	output wire io_connSS_0_data_availableTask_valid;
	output wire [127:0] io_connSS_0_data_availableTask_bits;
	output wire io_connSS_0_data_qOutTask_ready;
	input io_connSS_0_data_qOutTask_valid;
	input [127:0] io_connSS_0_data_qOutTask_bits;
	input io_connSS_1_ctrl_serveStealReq_valid;
	output wire io_connSS_1_ctrl_serveStealReq_ready;
	output wire io_connSS_1_data_qOutTask_ready;
	input io_connSS_1_data_qOutTask_valid;
	input [127:0] io_connSS_1_data_qOutTask_bits;
	input io_connSS_2_ctrl_serveStealReq_valid;
	output wire io_connSS_2_ctrl_serveStealReq_ready;
	output wire io_connSS_2_data_qOutTask_ready;
	input io_connSS_2_data_qOutTask_valid;
	input [127:0] io_connSS_2_data_qOutTask_bits;
	input io_connSS_3_ctrl_serveStealReq_valid;
	output wire io_connSS_3_ctrl_serveStealReq_ready;
	output wire io_connSS_3_data_qOutTask_ready;
	input io_connSS_3_data_qOutTask_valid;
	input [127:0] io_connSS_3_data_qOutTask_bits;
	input io_connSS_4_ctrl_serveStealReq_valid;
	output wire io_connSS_4_ctrl_serveStealReq_ready;
	output wire io_connSS_4_data_qOutTask_ready;
	input io_connSS_4_data_qOutTask_valid;
	input [127:0] io_connSS_4_data_qOutTask_bits;
	input io_connSS_5_ctrl_serveStealReq_valid;
	output wire io_connSS_5_ctrl_serveStealReq_ready;
	output wire io_connSS_5_data_qOutTask_ready;
	input io_connSS_5_data_qOutTask_valid;
	input [127:0] io_connSS_5_data_qOutTask_bits;
	input io_connSS_6_ctrl_serveStealReq_valid;
	output wire io_connSS_6_ctrl_serveStealReq_ready;
	output wire io_connSS_6_data_qOutTask_ready;
	input io_connSS_6_data_qOutTask_valid;
	input [127:0] io_connSS_6_data_qOutTask_bits;
	input io_connSS_7_ctrl_serveStealReq_valid;
	output wire io_connSS_7_ctrl_serveStealReq_ready;
	output wire io_connSS_7_data_qOutTask_ready;
	input io_connSS_7_data_qOutTask_valid;
	input [127:0] io_connSS_7_data_qOutTask_bits;
	input io_connSS_8_ctrl_serveStealReq_valid;
	output wire io_connSS_8_ctrl_serveStealReq_ready;
	output wire io_connSS_8_data_qOutTask_ready;
	input io_connSS_8_data_qOutTask_valid;
	input [127:0] io_connSS_8_data_qOutTask_bits;
	input io_connSS_9_ctrl_serveStealReq_valid;
	output wire io_connSS_9_ctrl_serveStealReq_ready;
	output wire io_connSS_9_data_qOutTask_ready;
	input io_connSS_9_data_qOutTask_valid;
	input [127:0] io_connSS_9_data_qOutTask_bits;
	input io_connSS_10_ctrl_serveStealReq_valid;
	output wire io_connSS_10_ctrl_serveStealReq_ready;
	output wire io_connSS_10_data_qOutTask_ready;
	input io_connSS_10_data_qOutTask_valid;
	input [127:0] io_connSS_10_data_qOutTask_bits;
	input io_connSS_11_ctrl_serveStealReq_valid;
	output wire io_connSS_11_ctrl_serveStealReq_ready;
	output wire io_connSS_11_data_qOutTask_ready;
	input io_connSS_11_data_qOutTask_valid;
	input [127:0] io_connSS_11_data_qOutTask_bits;
	input io_connSS_12_ctrl_serveStealReq_valid;
	output wire io_connSS_12_ctrl_serveStealReq_ready;
	output wire io_connSS_12_data_qOutTask_ready;
	input io_connSS_12_data_qOutTask_valid;
	input [127:0] io_connSS_12_data_qOutTask_bits;
	input io_connSS_13_ctrl_serveStealReq_valid;
	output wire io_connSS_13_ctrl_serveStealReq_ready;
	output wire io_connSS_13_data_qOutTask_ready;
	input io_connSS_13_data_qOutTask_valid;
	input [127:0] io_connSS_13_data_qOutTask_bits;
	input io_connSS_14_ctrl_serveStealReq_valid;
	output wire io_connSS_14_ctrl_serveStealReq_ready;
	output wire io_connSS_14_data_qOutTask_ready;
	input io_connSS_14_data_qOutTask_valid;
	input [127:0] io_connSS_14_data_qOutTask_bits;
	input io_connSS_15_ctrl_serveStealReq_valid;
	output wire io_connSS_15_ctrl_serveStealReq_ready;
	output wire io_connSS_15_data_qOutTask_ready;
	input io_connSS_15_data_qOutTask_valid;
	input [127:0] io_connSS_15_data_qOutTask_bits;
	input io_connSS_16_ctrl_serveStealReq_valid;
	output wire io_connSS_16_ctrl_serveStealReq_ready;
	output wire io_connSS_16_data_qOutTask_ready;
	input io_connSS_16_data_qOutTask_valid;
	input [127:0] io_connSS_16_data_qOutTask_bits;
	input io_connSS_17_ctrl_serveStealReq_valid;
	output wire io_connSS_17_ctrl_serveStealReq_ready;
	input io_connSS_17_ctrl_stealReq_valid;
	output wire io_connSS_17_ctrl_stealReq_ready;
	input io_connSS_17_data_availableTask_ready;
	output wire io_connSS_17_data_availableTask_valid;
	output wire [127:0] io_connSS_17_data_availableTask_bits;
	output wire io_connSS_17_data_qOutTask_ready;
	input io_connSS_17_data_qOutTask_valid;
	input [127:0] io_connSS_17_data_qOutTask_bits;
	input io_connSS_18_ctrl_serveStealReq_valid;
	output wire io_connSS_18_ctrl_serveStealReq_ready;
	input io_connSS_18_ctrl_stealReq_valid;
	output wire io_connSS_18_ctrl_stealReq_ready;
	input io_connSS_18_data_availableTask_ready;
	output wire io_connSS_18_data_availableTask_valid;
	output wire [127:0] io_connSS_18_data_availableTask_bits;
	output wire io_connSS_18_data_qOutTask_ready;
	input io_connSS_18_data_qOutTask_valid;
	input [127:0] io_connSS_18_data_qOutTask_bits;
	input io_connSS_19_ctrl_serveStealReq_valid;
	output wire io_connSS_19_ctrl_serveStealReq_ready;
	input io_connSS_19_ctrl_stealReq_valid;
	output wire io_connSS_19_ctrl_stealReq_ready;
	input io_connSS_19_data_availableTask_ready;
	output wire io_connSS_19_data_availableTask_valid;
	output wire [127:0] io_connSS_19_data_availableTask_bits;
	output wire io_connSS_19_data_qOutTask_ready;
	input io_connSS_19_data_qOutTask_valid;
	input [127:0] io_connSS_19_data_qOutTask_bits;
	input io_connSS_20_ctrl_serveStealReq_valid;
	output wire io_connSS_20_ctrl_serveStealReq_ready;
	input io_connSS_20_ctrl_stealReq_valid;
	output wire io_connSS_20_ctrl_stealReq_ready;
	input io_connSS_20_data_availableTask_ready;
	output wire io_connSS_20_data_availableTask_valid;
	output wire [127:0] io_connSS_20_data_availableTask_bits;
	output wire io_connSS_20_data_qOutTask_ready;
	input io_connSS_20_data_qOutTask_valid;
	input [127:0] io_connSS_20_data_qOutTask_bits;
	input io_connSS_21_ctrl_serveStealReq_valid;
	output wire io_connSS_21_ctrl_serveStealReq_ready;
	input io_connSS_21_ctrl_stealReq_valid;
	output wire io_connSS_21_ctrl_stealReq_ready;
	input io_connSS_21_data_availableTask_ready;
	output wire io_connSS_21_data_availableTask_valid;
	output wire [127:0] io_connSS_21_data_availableTask_bits;
	output wire io_connSS_21_data_qOutTask_ready;
	input io_connSS_21_data_qOutTask_valid;
	input [127:0] io_connSS_21_data_qOutTask_bits;
	input io_connSS_22_ctrl_serveStealReq_valid;
	output wire io_connSS_22_ctrl_serveStealReq_ready;
	input io_connSS_22_ctrl_stealReq_valid;
	output wire io_connSS_22_ctrl_stealReq_ready;
	input io_connSS_22_data_availableTask_ready;
	output wire io_connSS_22_data_availableTask_valid;
	output wire [127:0] io_connSS_22_data_availableTask_bits;
	output wire io_connSS_22_data_qOutTask_ready;
	input io_connSS_22_data_qOutTask_valid;
	input [127:0] io_connSS_22_data_qOutTask_bits;
	input io_connSS_23_ctrl_serveStealReq_valid;
	output wire io_connSS_23_ctrl_serveStealReq_ready;
	input io_connSS_23_ctrl_stealReq_valid;
	output wire io_connSS_23_ctrl_stealReq_ready;
	input io_connSS_23_data_availableTask_ready;
	output wire io_connSS_23_data_availableTask_valid;
	output wire [127:0] io_connSS_23_data_availableTask_bits;
	output wire io_connSS_23_data_qOutTask_ready;
	input io_connSS_23_data_qOutTask_valid;
	input [127:0] io_connSS_23_data_qOutTask_bits;
	input io_connSS_24_ctrl_serveStealReq_valid;
	output wire io_connSS_24_ctrl_serveStealReq_ready;
	input io_connSS_24_ctrl_stealReq_valid;
	output wire io_connSS_24_ctrl_stealReq_ready;
	input io_connSS_24_data_availableTask_ready;
	output wire io_connSS_24_data_availableTask_valid;
	output wire [127:0] io_connSS_24_data_availableTask_bits;
	output wire io_connSS_24_data_qOutTask_ready;
	input io_connSS_24_data_qOutTask_valid;
	input [127:0] io_connSS_24_data_qOutTask_bits;
	input io_connSS_25_ctrl_serveStealReq_valid;
	output wire io_connSS_25_ctrl_serveStealReq_ready;
	input io_connSS_25_ctrl_stealReq_valid;
	output wire io_connSS_25_ctrl_stealReq_ready;
	input io_connSS_25_data_availableTask_ready;
	output wire io_connSS_25_data_availableTask_valid;
	output wire [127:0] io_connSS_25_data_availableTask_bits;
	output wire io_connSS_25_data_qOutTask_ready;
	input io_connSS_25_data_qOutTask_valid;
	input [127:0] io_connSS_25_data_qOutTask_bits;
	input io_connSS_26_ctrl_serveStealReq_valid;
	output wire io_connSS_26_ctrl_serveStealReq_ready;
	input io_connSS_26_ctrl_stealReq_valid;
	output wire io_connSS_26_ctrl_stealReq_ready;
	input io_connSS_26_data_availableTask_ready;
	output wire io_connSS_26_data_availableTask_valid;
	output wire [127:0] io_connSS_26_data_availableTask_bits;
	output wire io_connSS_26_data_qOutTask_ready;
	input io_connSS_26_data_qOutTask_valid;
	input [127:0] io_connSS_26_data_qOutTask_bits;
	input io_connSS_27_ctrl_serveStealReq_valid;
	output wire io_connSS_27_ctrl_serveStealReq_ready;
	input io_connSS_27_ctrl_stealReq_valid;
	output wire io_connSS_27_ctrl_stealReq_ready;
	input io_connSS_27_data_availableTask_ready;
	output wire io_connSS_27_data_availableTask_valid;
	output wire [127:0] io_connSS_27_data_availableTask_bits;
	output wire io_connSS_27_data_qOutTask_ready;
	input io_connSS_27_data_qOutTask_valid;
	input [127:0] io_connSS_27_data_qOutTask_bits;
	input io_connSS_28_ctrl_serveStealReq_valid;
	output wire io_connSS_28_ctrl_serveStealReq_ready;
	input io_connSS_28_ctrl_stealReq_valid;
	output wire io_connSS_28_ctrl_stealReq_ready;
	input io_connSS_28_data_availableTask_ready;
	output wire io_connSS_28_data_availableTask_valid;
	output wire [127:0] io_connSS_28_data_availableTask_bits;
	output wire io_connSS_28_data_qOutTask_ready;
	input io_connSS_28_data_qOutTask_valid;
	input [127:0] io_connSS_28_data_qOutTask_bits;
	input io_connSS_29_ctrl_serveStealReq_valid;
	output wire io_connSS_29_ctrl_serveStealReq_ready;
	input io_connSS_29_ctrl_stealReq_valid;
	output wire io_connSS_29_ctrl_stealReq_ready;
	input io_connSS_29_data_availableTask_ready;
	output wire io_connSS_29_data_availableTask_valid;
	output wire [127:0] io_connSS_29_data_availableTask_bits;
	output wire io_connSS_29_data_qOutTask_ready;
	input io_connSS_29_data_qOutTask_valid;
	input [127:0] io_connSS_29_data_qOutTask_bits;
	input io_connSS_30_ctrl_serveStealReq_valid;
	output wire io_connSS_30_ctrl_serveStealReq_ready;
	input io_connSS_30_ctrl_stealReq_valid;
	output wire io_connSS_30_ctrl_stealReq_ready;
	input io_connSS_30_data_availableTask_ready;
	output wire io_connSS_30_data_availableTask_valid;
	output wire [127:0] io_connSS_30_data_availableTask_bits;
	output wire io_connSS_30_data_qOutTask_ready;
	input io_connSS_30_data_qOutTask_valid;
	input [127:0] io_connSS_30_data_qOutTask_bits;
	input io_connSS_31_ctrl_serveStealReq_valid;
	output wire io_connSS_31_ctrl_serveStealReq_ready;
	input io_connSS_31_ctrl_stealReq_valid;
	output wire io_connSS_31_ctrl_stealReq_ready;
	input io_connSS_31_data_availableTask_ready;
	output wire io_connSS_31_data_availableTask_valid;
	output wire [127:0] io_connSS_31_data_availableTask_bits;
	output wire io_connSS_31_data_qOutTask_ready;
	input io_connSS_31_data_qOutTask_valid;
	input [127:0] io_connSS_31_data_qOutTask_bits;
	input io_connSS_32_ctrl_serveStealReq_valid;
	output wire io_connSS_32_ctrl_serveStealReq_ready;
	input io_connSS_32_ctrl_stealReq_valid;
	output wire io_connSS_32_ctrl_stealReq_ready;
	input io_connSS_32_data_availableTask_ready;
	output wire io_connSS_32_data_availableTask_valid;
	output wire [127:0] io_connSS_32_data_availableTask_bits;
	output wire io_connSS_32_data_qOutTask_ready;
	input io_connSS_32_data_qOutTask_valid;
	input [127:0] io_connSS_32_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	wire _ctrlunits_32_io_reqTaskOut;
	wire _ctrlunits_31_io_reqTaskOut;
	wire _ctrlunits_30_io_reqTaskOut;
	wire _ctrlunits_29_io_reqTaskOut;
	wire _ctrlunits_28_io_reqTaskOut;
	wire _ctrlunits_27_io_reqTaskOut;
	wire _ctrlunits_26_io_reqTaskOut;
	wire _ctrlunits_25_io_reqTaskOut;
	wire _ctrlunits_24_io_reqTaskOut;
	wire _ctrlunits_23_io_reqTaskOut;
	wire _ctrlunits_22_io_reqTaskOut;
	wire _ctrlunits_21_io_reqTaskOut;
	wire _ctrlunits_20_io_reqTaskOut;
	wire _ctrlunits_19_io_reqTaskOut;
	wire _ctrlunits_18_io_reqTaskOut;
	wire _ctrlunits_17_io_reqTaskOut;
	wire _ctrlunits_16_io_reqTaskOut;
	wire _ctrlunits_15_io_reqTaskOut;
	wire _ctrlunits_14_io_reqTaskOut;
	wire _ctrlunits_13_io_reqTaskOut;
	wire _ctrlunits_12_io_reqTaskOut;
	wire _ctrlunits_11_io_reqTaskOut;
	wire _ctrlunits_10_io_reqTaskOut;
	wire _ctrlunits_9_io_reqTaskOut;
	wire _ctrlunits_8_io_reqTaskOut;
	wire _ctrlunits_7_io_reqTaskOut;
	wire _ctrlunits_6_io_reqTaskOut;
	wire _ctrlunits_5_io_reqTaskOut;
	wire _ctrlunits_4_io_reqTaskOut;
	wire _ctrlunits_3_io_reqTaskOut;
	wire _ctrlunits_2_io_reqTaskOut;
	wire _ctrlunits_1_io_reqTaskOut;
	wire _ctrlunits_0_io_reqTaskOut;
	wire [127:0] _dataUnits_32_io_taskOut;
	wire _dataUnits_32_io_validOut;
	wire [127:0] _dataUnits_31_io_taskOut;
	wire _dataUnits_31_io_validOut;
	wire [127:0] _dataUnits_30_io_taskOut;
	wire _dataUnits_30_io_validOut;
	wire [127:0] _dataUnits_29_io_taskOut;
	wire _dataUnits_29_io_validOut;
	wire [127:0] _dataUnits_28_io_taskOut;
	wire _dataUnits_28_io_validOut;
	wire [127:0] _dataUnits_27_io_taskOut;
	wire _dataUnits_27_io_validOut;
	wire [127:0] _dataUnits_26_io_taskOut;
	wire _dataUnits_26_io_validOut;
	wire [127:0] _dataUnits_25_io_taskOut;
	wire _dataUnits_25_io_validOut;
	wire [127:0] _dataUnits_24_io_taskOut;
	wire _dataUnits_24_io_validOut;
	wire [127:0] _dataUnits_23_io_taskOut;
	wire _dataUnits_23_io_validOut;
	wire [127:0] _dataUnits_22_io_taskOut;
	wire _dataUnits_22_io_validOut;
	wire [127:0] _dataUnits_21_io_taskOut;
	wire _dataUnits_21_io_validOut;
	wire [127:0] _dataUnits_20_io_taskOut;
	wire _dataUnits_20_io_validOut;
	wire [127:0] _dataUnits_19_io_taskOut;
	wire _dataUnits_19_io_validOut;
	wire [127:0] _dataUnits_18_io_taskOut;
	wire _dataUnits_18_io_validOut;
	wire [127:0] _dataUnits_17_io_taskOut;
	wire _dataUnits_17_io_validOut;
	wire [127:0] _dataUnits_16_io_taskOut;
	wire _dataUnits_16_io_validOut;
	wire [127:0] _dataUnits_15_io_taskOut;
	wire _dataUnits_15_io_validOut;
	wire [127:0] _dataUnits_14_io_taskOut;
	wire _dataUnits_14_io_validOut;
	wire [127:0] _dataUnits_13_io_taskOut;
	wire _dataUnits_13_io_validOut;
	wire [127:0] _dataUnits_12_io_taskOut;
	wire _dataUnits_12_io_validOut;
	wire [127:0] _dataUnits_11_io_taskOut;
	wire _dataUnits_11_io_validOut;
	wire [127:0] _dataUnits_10_io_taskOut;
	wire _dataUnits_10_io_validOut;
	wire [127:0] _dataUnits_9_io_taskOut;
	wire _dataUnits_9_io_validOut;
	wire [127:0] _dataUnits_8_io_taskOut;
	wire _dataUnits_8_io_validOut;
	wire [127:0] _dataUnits_7_io_taskOut;
	wire _dataUnits_7_io_validOut;
	wire [127:0] _dataUnits_6_io_taskOut;
	wire _dataUnits_6_io_validOut;
	wire [127:0] _dataUnits_5_io_taskOut;
	wire _dataUnits_5_io_validOut;
	wire [127:0] _dataUnits_4_io_taskOut;
	wire _dataUnits_4_io_validOut;
	wire [127:0] _dataUnits_3_io_taskOut;
	wire _dataUnits_3_io_validOut;
	wire [127:0] _dataUnits_2_io_taskOut;
	wire _dataUnits_2_io_validOut;
	wire [127:0] _dataUnits_1_io_taskOut;
	wire _dataUnits_1_io_validOut;
	wire [127:0] _dataUnits_0_io_taskOut;
	wire _dataUnits_0_io_validOut;
	SchedulerNetworkDataUnit_65 dataUnits_0(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_32_io_taskOut),
		.io_taskOut(_dataUnits_0_io_taskOut),
		.io_validIn(_dataUnits_32_io_validOut),
		.io_validOut(_dataUnits_0_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_0_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_0_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_0_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_0_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_0_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_0_data_qOutTask_bits),
		.io_occupied(io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerNetworkDataUnit_65 dataUnits_1(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_0_io_taskOut),
		.io_taskOut(_dataUnits_1_io_taskOut),
		.io_validIn(_dataUnits_0_io_validOut),
		.io_validOut(_dataUnits_1_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_1_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_1_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_1_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_2(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_1_io_taskOut),
		.io_taskOut(_dataUnits_2_io_taskOut),
		.io_validIn(_dataUnits_1_io_validOut),
		.io_validOut(_dataUnits_2_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_2_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_2_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_2_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_3(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_2_io_taskOut),
		.io_taskOut(_dataUnits_3_io_taskOut),
		.io_validIn(_dataUnits_2_io_validOut),
		.io_validOut(_dataUnits_3_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_3_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_3_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_3_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_4(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_3_io_taskOut),
		.io_taskOut(_dataUnits_4_io_taskOut),
		.io_validIn(_dataUnits_3_io_validOut),
		.io_validOut(_dataUnits_4_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_4_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_4_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_4_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_5(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_4_io_taskOut),
		.io_taskOut(_dataUnits_5_io_taskOut),
		.io_validIn(_dataUnits_4_io_validOut),
		.io_validOut(_dataUnits_5_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_5_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_5_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_5_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_6(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_5_io_taskOut),
		.io_taskOut(_dataUnits_6_io_taskOut),
		.io_validIn(_dataUnits_5_io_validOut),
		.io_validOut(_dataUnits_6_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_6_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_6_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_6_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_7(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_6_io_taskOut),
		.io_taskOut(_dataUnits_7_io_taskOut),
		.io_validIn(_dataUnits_6_io_validOut),
		.io_validOut(_dataUnits_7_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_7_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_7_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_7_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_8(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_7_io_taskOut),
		.io_taskOut(_dataUnits_8_io_taskOut),
		.io_validIn(_dataUnits_7_io_validOut),
		.io_validOut(_dataUnits_8_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_8_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_8_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_8_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_9(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_8_io_taskOut),
		.io_taskOut(_dataUnits_9_io_taskOut),
		.io_validIn(_dataUnits_8_io_validOut),
		.io_validOut(_dataUnits_9_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_9_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_9_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_9_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_10(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_9_io_taskOut),
		.io_taskOut(_dataUnits_10_io_taskOut),
		.io_validIn(_dataUnits_9_io_validOut),
		.io_validOut(_dataUnits_10_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_10_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_10_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_10_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_11(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_10_io_taskOut),
		.io_taskOut(_dataUnits_11_io_taskOut),
		.io_validIn(_dataUnits_10_io_validOut),
		.io_validOut(_dataUnits_11_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_11_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_11_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_11_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_12(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_11_io_taskOut),
		.io_taskOut(_dataUnits_12_io_taskOut),
		.io_validIn(_dataUnits_11_io_validOut),
		.io_validOut(_dataUnits_12_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_12_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_12_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_12_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_13(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_12_io_taskOut),
		.io_taskOut(_dataUnits_13_io_taskOut),
		.io_validIn(_dataUnits_12_io_validOut),
		.io_validOut(_dataUnits_13_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_13_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_13_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_13_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_14(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_13_io_taskOut),
		.io_taskOut(_dataUnits_14_io_taskOut),
		.io_validIn(_dataUnits_13_io_validOut),
		.io_validOut(_dataUnits_14_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_14_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_14_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_14_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_15(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_14_io_taskOut),
		.io_taskOut(_dataUnits_15_io_taskOut),
		.io_validIn(_dataUnits_14_io_validOut),
		.io_validOut(_dataUnits_15_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_15_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_15_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_15_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_16(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_15_io_taskOut),
		.io_taskOut(_dataUnits_16_io_taskOut),
		.io_validIn(_dataUnits_15_io_validOut),
		.io_validOut(_dataUnits_16_io_validOut),
		.io_connSS_availableTask_ready(1'h0),
		.io_connSS_availableTask_valid(),
		.io_connSS_availableTask_bits(),
		.io_connSS_qOutTask_ready(io_connSS_16_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_16_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_16_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_17(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_16_io_taskOut),
		.io_taskOut(_dataUnits_17_io_taskOut),
		.io_validIn(_dataUnits_16_io_validOut),
		.io_validOut(_dataUnits_17_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_17_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_17_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_17_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_17_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_17_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_17_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_18(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_17_io_taskOut),
		.io_taskOut(_dataUnits_18_io_taskOut),
		.io_validIn(_dataUnits_17_io_validOut),
		.io_validOut(_dataUnits_18_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_18_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_18_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_18_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_18_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_18_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_18_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_19(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_18_io_taskOut),
		.io_taskOut(_dataUnits_19_io_taskOut),
		.io_validIn(_dataUnits_18_io_validOut),
		.io_validOut(_dataUnits_19_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_19_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_19_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_19_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_19_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_19_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_19_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_20(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_19_io_taskOut),
		.io_taskOut(_dataUnits_20_io_taskOut),
		.io_validIn(_dataUnits_19_io_validOut),
		.io_validOut(_dataUnits_20_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_20_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_20_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_20_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_20_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_20_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_20_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_21(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_20_io_taskOut),
		.io_taskOut(_dataUnits_21_io_taskOut),
		.io_validIn(_dataUnits_20_io_validOut),
		.io_validOut(_dataUnits_21_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_21_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_21_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_21_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_21_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_21_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_21_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_22(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_21_io_taskOut),
		.io_taskOut(_dataUnits_22_io_taskOut),
		.io_validIn(_dataUnits_21_io_validOut),
		.io_validOut(_dataUnits_22_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_22_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_22_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_22_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_22_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_22_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_22_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_23(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_22_io_taskOut),
		.io_taskOut(_dataUnits_23_io_taskOut),
		.io_validIn(_dataUnits_22_io_validOut),
		.io_validOut(_dataUnits_23_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_23_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_23_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_23_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_23_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_23_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_23_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_24(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_23_io_taskOut),
		.io_taskOut(_dataUnits_24_io_taskOut),
		.io_validIn(_dataUnits_23_io_validOut),
		.io_validOut(_dataUnits_24_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_24_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_24_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_24_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_24_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_24_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_24_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_25(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_24_io_taskOut),
		.io_taskOut(_dataUnits_25_io_taskOut),
		.io_validIn(_dataUnits_24_io_validOut),
		.io_validOut(_dataUnits_25_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_25_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_25_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_25_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_25_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_25_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_25_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_26(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_25_io_taskOut),
		.io_taskOut(_dataUnits_26_io_taskOut),
		.io_validIn(_dataUnits_25_io_validOut),
		.io_validOut(_dataUnits_26_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_26_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_26_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_26_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_26_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_26_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_26_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_27(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_26_io_taskOut),
		.io_taskOut(_dataUnits_27_io_taskOut),
		.io_validIn(_dataUnits_26_io_validOut),
		.io_validOut(_dataUnits_27_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_27_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_27_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_27_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_27_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_27_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_27_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_28(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_27_io_taskOut),
		.io_taskOut(_dataUnits_28_io_taskOut),
		.io_validIn(_dataUnits_27_io_validOut),
		.io_validOut(_dataUnits_28_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_28_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_28_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_28_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_28_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_28_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_28_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_29(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_28_io_taskOut),
		.io_taskOut(_dataUnits_29_io_taskOut),
		.io_validIn(_dataUnits_28_io_validOut),
		.io_validOut(_dataUnits_29_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_29_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_29_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_29_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_29_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_29_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_29_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_30(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_29_io_taskOut),
		.io_taskOut(_dataUnits_30_io_taskOut),
		.io_validIn(_dataUnits_29_io_validOut),
		.io_validOut(_dataUnits_30_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_30_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_30_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_30_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_30_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_30_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_30_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_31(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_30_io_taskOut),
		.io_taskOut(_dataUnits_31_io_taskOut),
		.io_validIn(_dataUnits_30_io_validOut),
		.io_validOut(_dataUnits_31_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_31_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_31_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_31_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_31_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_31_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_31_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkDataUnit_65 dataUnits_32(
		.clock(clock),
		.reset(reset),
		.io_taskIn(_dataUnits_31_io_taskOut),
		.io_taskOut(_dataUnits_32_io_taskOut),
		.io_validIn(_dataUnits_31_io_validOut),
		.io_validOut(_dataUnits_32_io_validOut),
		.io_connSS_availableTask_ready(io_connSS_32_data_availableTask_ready),
		.io_connSS_availableTask_valid(io_connSS_32_data_availableTask_valid),
		.io_connSS_availableTask_bits(io_connSS_32_data_availableTask_bits),
		.io_connSS_qOutTask_ready(io_connSS_32_data_qOutTask_ready),
		.io_connSS_qOutTask_valid(io_connSS_32_data_qOutTask_valid),
		.io_connSS_qOutTask_bits(io_connSS_32_data_qOutTask_bits),
		.io_occupied()
	);
	SchedulerNetworkControlUnit ctrlunits_0(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_1_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_0_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_0_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_0_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_1(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_2_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_1_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_1_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_1_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_2(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_3_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_2_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_2_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_2_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_3(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_4_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_3_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_3_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_3_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_4(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_5_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_4_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_4_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_4_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_5(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_6_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_5_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_5_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_5_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_6(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_7_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_6_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_6_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_6_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_7(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_8_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_7_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_7_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_7_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_8(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_9_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_8_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_8_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_8_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_9(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_10_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_9_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_9_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_9_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_10(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_11_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_10_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_10_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_10_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_11(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_12_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_11_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_11_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_11_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_12(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_13_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_12_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_12_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_12_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_13(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_14_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_13_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_13_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_13_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_14(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_15_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_14_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_14_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_14_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_15(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_16_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_15_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_15_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_15_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_16(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_17_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_16_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_16_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_16_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(1'h0),
		.io_connSS_stealReq_ready()
	);
	SchedulerNetworkControlUnit ctrlunits_17(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_18_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_17_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_17_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_17_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_17_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_18(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_19_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_18_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_18_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_18_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_18_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_19(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_20_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_19_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_19_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_19_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_19_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_20(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_21_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_20_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_20_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_20_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_20_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_21(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_22_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_21_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_21_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_21_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_21_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_22(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_23_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_22_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_22_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_22_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_22_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_23(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_24_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_23_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_23_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_23_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_23_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_24(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_25_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_24_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_24_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_24_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_24_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_25(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_26_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_25_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_25_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_25_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_25_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_26(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_27_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_26_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_26_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_26_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_26_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_27(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_28_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_27_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_27_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_27_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_27_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_28(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_29_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_28_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_28_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_28_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_28_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_29(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_30_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_29_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_29_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_29_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_29_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_30(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_31_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_30_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_30_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_30_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_30_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_31(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_32_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_31_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_31_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_31_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_31_ctrl_stealReq_ready)
	);
	SchedulerNetworkControlUnit ctrlunits_32(
		.clock(clock),
		.reset(reset),
		.io_reqTaskIn(_ctrlunits_0_io_reqTaskOut),
		.io_reqTaskOut(_ctrlunits_32_io_reqTaskOut),
		.io_connSS_serveStealReq_valid(io_connSS_32_ctrl_serveStealReq_valid),
		.io_connSS_serveStealReq_ready(io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_stealReq_valid(io_connSS_32_ctrl_stealReq_valid),
		.io_connSS_stealReq_ready(io_connSS_32_ctrl_stealReq_ready)
	);
endmodule
module SchedulerClient_64 (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_ctrl_stealReq_valid,
	io_connNetwork_ctrl_stealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_connQ_currLength,
	io_connQ_push_ready,
	io_connQ_push_valid,
	io_connQ_push_bits,
	io_connQ_pop_ready,
	io_connQ_pop_valid,
	io_connQ_pop_bits
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_ctrl_stealReq_valid;
	input io_connNetwork_ctrl_stealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [127:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [127:0] io_connNetwork_data_qOutTask_bits;
	input [7:0] io_connQ_currLength;
	input io_connQ_push_ready;
	output wire io_connQ_push_valid;
	output wire [127:0] io_connQ_push_bits;
	output wire io_connQ_pop_ready;
	input io_connQ_pop_valid;
	input [127:0] io_connQ_pop_bits;
	reg [2:0] stateReg;
	reg [127:0] stolenTaskReg;
	reg [127:0] giveTaskReg;
	reg [31:0] requestKilledCount;
	reg [31:0] requestTaskCount;
	wire _GEN = stateReg == 3'h0;
	wire _GEN_0 = io_connQ_currLength < 8'h66;
	wire _GEN_1 = stateReg == 3'h2;
	wire _GEN_2 = requestKilledCount == 32'h00000000;
	wire _GEN_3 = stateReg == 3'h3;
	wire _GEN_4 = _GEN | _GEN_1;
	wire _GEN_5 = stateReg == 3'h4;
	wire _GEN_6 = io_connQ_currLength == 8'h00;
	wire _GEN_7 = stateReg == 3'h5;
	wire _GEN_8 = ((_GEN | _GEN_1) | _GEN_3) | _GEN_5;
	wire _GEN_9 = stateReg == 3'h6;
	wire io_connNetwork_ctrl_stealReq_valid_0 = ((|requestTaskCount & ~(_GEN_9 & _GEN_0)) & ~(_GEN_5 & _GEN_6)) & ~(_GEN_1 & _GEN_2);
	always @(posedge clock)
		if (reset) begin
			stateReg <= 3'h0;
			stolenTaskReg <= 128'h00000000000000000000000000000000;
			giveTaskReg <= 128'h00000000000000000000000000000000;
			requestKilledCount <= 32'h00000021;
			requestTaskCount <= 32'h00000000;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_10;
			reg _GEN_11;
			reg _GEN_12;
			reg _GEN_13;
			reg _GEN_14;
			reg _GEN_15;
			reg [23:0] _GEN_16;
			_GEN_10 = io_connQ_currLength > 8'h65;
			_GEN_11 = io_connQ_currLength > 8'h7e;
			_GEN_12 = io_connQ_pop_valid | ~_GEN_6;
			_GEN_13 = io_connQ_currLength[7] | (io_connNetwork_ctrl_serveStealReq_ready & _GEN_10);
			_GEN_14 = _GEN_0 & io_connNetwork_ctrl_serveStealReq_ready;
			_GEN_15 = _GEN_14 | _GEN_0;
			_GEN_16 = {stateReg, (_GEN_13 ? 3'h4 : {~_GEN_15, 2'h2}), (io_connNetwork_data_qOutTask_ready ? 3'h0 : 3'h5), (io_connQ_pop_valid ? 3'h5 : (_GEN_6 ? 3'h2 : 3'h4)), (io_connQ_push_ready ? 3'h0 : (_GEN_11 ? 3'h5 : 3'h3)), (io_connNetwork_data_availableTask_valid ? 3'h3 : (_GEN_10 ? 3'h0 : (_GEN_2 ? stateReg : 3'h2))), stateReg, (_GEN_0 ? 3'h2 : (io_connQ_currLength[7] ? 3'h4 : (io_connQ_currLength > 8'h66 ? 3'h6 : 3'h0)))};
			stateReg <= _GEN_16[stateReg * 3+:3];
			if (_GEN | ~(_GEN_1 & io_connNetwork_data_availableTask_valid))
				;
			else
				stolenTaskReg <= io_connNetwork_data_availableTask_bits;
			if (~_GEN_4) begin
				if (_GEN_3) begin
					if (io_connQ_push_ready | ~_GEN_11)
						;
					else
						giveTaskReg <= stolenTaskReg;
				end
				else if (_GEN_5 & io_connQ_pop_valid)
					giveTaskReg <= io_connQ_pop_bits;
			end
			if (_GEN) begin
				if (_GEN_0)
					requestKilledCount <= 32'h00000023;
			end
			else if (_GEN_1) begin
				if (io_connNetwork_ctrl_serveStealReq_ready)
					requestKilledCount <= 32'h00000023;
				else
					requestKilledCount <= requestKilledCount - 32'h00000001;
			end
			else if (_GEN_3 | (_GEN_5 ? _GEN_12 : ((_GEN_7 | ~_GEN_9) | _GEN_13) | ~_GEN_15))
				;
			else
				requestKilledCount <= 32'h00000023;
			if (io_connNetwork_ctrl_stealReq_valid_0 & io_connNetwork_ctrl_stealReq_ready)
				requestTaskCount <= requestTaskCount - 32'h00000001;
			else begin : sv2v_autoblock_2
				reg [31:0] _GEN_17;
				reg [255:0] _GEN_18;
				_GEN_17 = ((_GEN_7 | ~_GEN_9) | _GEN_13 ? requestTaskCount : (_GEN_14 ? requestTaskCount + 32'h00000002 : (_GEN_0 ? requestTaskCount + 32'h00000001 : requestTaskCount)));
				_GEN_18 = {_GEN_17, _GEN_17, requestTaskCount, (_GEN_12 ? requestTaskCount : requestTaskCount + 32'h00000001), requestTaskCount, ((io_connNetwork_data_availableTask_valid | _GEN_10) | ~_GEN_2 ? requestTaskCount : requestTaskCount + 32'h00000001), _GEN_17, (_GEN_0 ? requestTaskCount + 32'h00000001 : requestTaskCount)};
				requestTaskCount <= _GEN_18[stateReg * 32+:32];
			end
		end
	assign io_connNetwork_ctrl_serveStealReq_valid = ~((((_GEN | _GEN_1) | _GEN_3) | _GEN_5) | _GEN_7) & _GEN_9;
	assign io_connNetwork_ctrl_stealReq_valid = io_connNetwork_ctrl_stealReq_valid_0;
	assign io_connNetwork_data_availableTask_ready = ~_GEN & _GEN_1;
	assign io_connNetwork_data_qOutTask_valid = ~_GEN_8 & _GEN_7;
	assign io_connNetwork_data_qOutTask_bits = (_GEN_8 | ~_GEN_7 ? 128'h00000000000000000000000000000000 : giveTaskReg);
	assign io_connQ_push_valid = ~_GEN_4 & _GEN_3;
	assign io_connQ_push_bits = (_GEN_4 | ~_GEN_3 ? 128'h00000000000000000000000000000000 : stolenTaskReg);
	assign io_connQ_pop_ready = ~((_GEN | _GEN_1) | _GEN_3) & _GEN_5;
endmodule
module hw_deque_64 (
	clock,
	reset,
	io_connVec_0_pop_ready,
	io_connVec_0_pop_valid,
	io_connVec_1_currLength,
	io_connVec_1_push_ready,
	io_connVec_1_push_valid,
	io_connVec_1_push_bits,
	io_connVec_1_pop_ready,
	io_connVec_1_pop_valid,
	io_connVec_1_pop_bits
);
	input clock;
	input reset;
	input io_connVec_0_pop_ready;
	output wire io_connVec_0_pop_valid;
	output wire [8:0] io_connVec_1_currLength;
	output wire io_connVec_1_push_ready;
	input io_connVec_1_push_valid;
	input [127:0] io_connVec_1_push_bits;
	input io_connVec_1_pop_ready;
	output wire io_connVec_1_pop_valid;
	output wire [127:0] io_connVec_1_pop_bits;
	wire [127:0] _bramMem_b_dout;
	reg [8:0] sideReg_0;
	reg [8:0] sideReg_1;
	reg readLatency_0;
	reg readLatency_1;
	reg writeLatency_0;
	reg writeLatency_1;
	reg [2:0] stateRegs_0;
	reg [2:0] stateRegs_1;
	wire _GEN = stateRegs_0 == 3'h0;
	wire _GEN_0 = stateRegs_1 == 3'h0;
	wire _GEN_1 = stateRegs_0 == 3'h1;
	wire _GEN_2 = stateRegs_0 == 3'h2;
	wire _GEN_3 = sideReg_0 == 9'h081;
	wire _GEN_4 = stateRegs_0 == 3'h4;
	wire [8:0] _bramMem_io_a_addr_T_2 = sideReg_0 + 9'h001;
	wire _GEN_5 = (_GEN | _GEN_1) | _GEN_2;
	wire _GEN_6 = stateRegs_1 == 3'h1;
	wire _GEN_7 = stateRegs_1 == 3'h2;
	wire _GEN_8 = sideReg_1 == 9'h000;
	wire _GEN_9 = stateRegs_1 == 3'h4;
	wire [8:0] _bramMem_io_b_addr_T_6 = sideReg_1 - 9'h001;
	wire _GEN_10 = (_GEN_0 | _GEN_6) | _GEN_7;
	wire _GEN_11 = stateRegs_1 == 3'h3;
	wire [8:0] currLen = (sideReg_0 > sideReg_1 ? ((sideReg_1 + 9'h082) - sideReg_0) - 9'h001 : (sideReg_1 - sideReg_0) - 9'h001);
	always @(posedge clock)
		if (reset) begin
			sideReg_0 <= 9'h000;
			sideReg_1 <= 9'h001;
			readLatency_0 <= 1'h0;
			readLatency_1 <= 1'h0;
			writeLatency_0 <= 1'h0;
			writeLatency_1 <= 1'h0;
			stateRegs_0 <= 3'h0;
			stateRegs_1 <= 3'h0;
		end
		else begin : sv2v_autoblock_1
			reg [23:0] _GEN_12;
			reg [23:0] _GEN_13;
			_GEN_12 = {stateRegs_0, stateRegs_0, stateRegs_0, 6'h00, (readLatency_0 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_0, 2'h2, (io_connVec_0_pop_ready & |currLen[8:1]) | ((io_connVec_0_pop_ready & _GEN_0) & |currLen), 1'h0};
			_GEN_13 = {stateRegs_1, stateRegs_1, stateRegs_1, 6'h00, (readLatency_1 ? 3'h2 : 3'h4), 1'h0, ~writeLatency_1, 1'h1, (io_connVec_1_push_valid & (currLen < 9'h081) ? 3'h1 : {1'h0, (io_connVec_1_pop_ready & |currLen[8:1]) | (((io_connVec_1_pop_ready & ~io_connVec_0_pop_ready) & |currLen) & (stateRegs_0 != 3'h4)), 1'h0})};
			if (~_GEN_5) begin
				if (_GEN_4) begin
					if (_GEN_3)
						sideReg_0 <= 9'h000;
					else
						sideReg_0 <= _bramMem_io_a_addr_T_2;
				end
				else if (stateRegs_0 == 3'h3) begin
					if (sideReg_0 == 9'h000)
						sideReg_0 <= 9'h081;
					else
						sideReg_0 <= sideReg_0 - 9'h001;
				end
			end
			if (~_GEN_10) begin
				if (_GEN_9) begin
					if (_GEN_8)
						sideReg_1 <= 9'h081;
					else
						sideReg_1 <= _bramMem_io_b_addr_T_6;
				end
				else if (_GEN_11) begin
					if (sideReg_1 == 9'h081)
						sideReg_1 <= 9'h000;
					else
						sideReg_1 <= sideReg_1 + 9'h001;
				end
			end
			readLatency_0 <= (((_GEN | _GEN_1) | ~_GEN_2) | (readLatency_0 - 1'h1)) & readLatency_0;
			readLatency_1 <= (((_GEN_0 | _GEN_6) | ~_GEN_7) | (readLatency_1 - 1'h1)) & readLatency_1;
			writeLatency_0 <= ((_GEN | ~_GEN_1) | (writeLatency_0 - 1'h1)) & writeLatency_0;
			writeLatency_1 <= ((_GEN_0 | ~_GEN_6) | (writeLatency_1 - 1'h1)) & writeLatency_1;
			stateRegs_0 <= _GEN_12[stateRegs_0 * 3+:3];
			stateRegs_1 <= _GEN_13[stateRegs_1 * 3+:3];
		end
	DualPortBRAM #(
		.ADDR(10),
		.DATA(128)
	) bramMem(
		.clk(clock),
		.rst(reset),
		.a_addr((_GEN ? 10'h3ff : (_GEN_1 ? {1'h0, sideReg_0} : (_GEN_2 ? (_GEN_3 ? 10'h000 : {1'h0, sideReg_0 + 9'h001}) : (_GEN_4 ? (_GEN_3 ? 10'h000 : {1'h0, _bramMem_io_a_addr_T_2}) : 10'h3ff))))),
		.a_din(128'h00000000000000000000000000000000),
		.a_wr(~_GEN & _GEN_1),
		.a_dout(),
		.b_addr((_GEN_0 ? 10'h3ff : (_GEN_6 ? {1'h0, sideReg_1} : (_GEN_7 ? (_GEN_8 ? 10'h081 : {1'h0, sideReg_1 - 9'h001}) : (_GEN_9 ? (_GEN_8 ? 10'h081 : {1'h0, _bramMem_io_b_addr_T_6}) : 10'h3ff))))),
		.b_din(io_connVec_1_push_bits),
		.b_wr(~_GEN_0 & _GEN_6),
		.b_dout(_bramMem_b_dout)
	);
	assign io_connVec_0_pop_valid = ~_GEN_5 & _GEN_4;
	assign io_connVec_1_currLength = currLen;
	assign io_connVec_1_push_ready = ~(((_GEN_0 | _GEN_6) | _GEN_7) | _GEN_9) & _GEN_11;
	assign io_connVec_1_pop_valid = ~_GEN_10 & _GEN_9;
	assign io_connVec_1_pop_bits = (_GEN_10 | ~_GEN_9 ? 128'h00000000000000000000000000000000 : _bramMem_b_dout);
endmodule
module SchedulerLocalNetwork_1 (
	clock,
	reset,
	io_connPE_0_pop_ready,
	io_connPE_0_pop_valid,
	io_connPE_1_pop_ready,
	io_connPE_1_pop_valid,
	io_connPE_2_pop_ready,
	io_connPE_2_pop_valid,
	io_connPE_3_pop_ready,
	io_connPE_3_pop_valid,
	io_connPE_4_pop_ready,
	io_connPE_4_pop_valid,
	io_connPE_5_pop_ready,
	io_connPE_5_pop_valid,
	io_connPE_6_pop_ready,
	io_connPE_6_pop_valid,
	io_connPE_7_pop_ready,
	io_connPE_7_pop_valid,
	io_connPE_8_pop_ready,
	io_connPE_8_pop_valid,
	io_connPE_9_pop_ready,
	io_connPE_9_pop_valid,
	io_connPE_10_pop_ready,
	io_connPE_10_pop_valid,
	io_connPE_11_pop_ready,
	io_connPE_11_pop_valid,
	io_connPE_12_pop_ready,
	io_connPE_12_pop_valid,
	io_connPE_13_pop_ready,
	io_connPE_13_pop_valid,
	io_connPE_14_pop_ready,
	io_connPE_14_pop_valid,
	io_connPE_15_pop_ready,
	io_connPE_15_pop_valid,
	io_connVSS_0_ctrl_serveStealReq_valid,
	io_connVSS_0_ctrl_serveStealReq_ready,
	io_connVSS_0_data_availableTask_ready,
	io_connVSS_0_data_availableTask_valid,
	io_connVSS_0_data_availableTask_bits,
	io_connVSS_0_data_qOutTask_ready,
	io_connVSS_0_data_qOutTask_valid,
	io_connVSS_0_data_qOutTask_bits,
	io_connVAS_0_ctrl_serveStealReq_valid,
	io_connVAS_0_ctrl_serveStealReq_ready,
	io_connVAS_0_data_qOutTask_ready,
	io_connVAS_0_data_qOutTask_valid,
	io_connVAS_0_data_qOutTask_bits,
	io_connVAS_1_ctrl_serveStealReq_valid,
	io_connVAS_1_ctrl_serveStealReq_ready,
	io_connVAS_1_data_qOutTask_ready,
	io_connVAS_1_data_qOutTask_valid,
	io_connVAS_1_data_qOutTask_bits,
	io_connVAS_2_ctrl_serveStealReq_valid,
	io_connVAS_2_ctrl_serveStealReq_ready,
	io_connVAS_2_data_qOutTask_ready,
	io_connVAS_2_data_qOutTask_valid,
	io_connVAS_2_data_qOutTask_bits,
	io_connVAS_3_ctrl_serveStealReq_valid,
	io_connVAS_3_ctrl_serveStealReq_ready,
	io_connVAS_3_data_qOutTask_ready,
	io_connVAS_3_data_qOutTask_valid,
	io_connVAS_3_data_qOutTask_bits,
	io_connVAS_4_ctrl_serveStealReq_valid,
	io_connVAS_4_ctrl_serveStealReq_ready,
	io_connVAS_4_data_qOutTask_ready,
	io_connVAS_4_data_qOutTask_valid,
	io_connVAS_4_data_qOutTask_bits,
	io_connVAS_5_ctrl_serveStealReq_valid,
	io_connVAS_5_ctrl_serveStealReq_ready,
	io_connVAS_5_data_qOutTask_ready,
	io_connVAS_5_data_qOutTask_valid,
	io_connVAS_5_data_qOutTask_bits,
	io_connVAS_6_ctrl_serveStealReq_valid,
	io_connVAS_6_ctrl_serveStealReq_ready,
	io_connVAS_6_data_qOutTask_ready,
	io_connVAS_6_data_qOutTask_valid,
	io_connVAS_6_data_qOutTask_bits,
	io_connVAS_7_ctrl_serveStealReq_valid,
	io_connVAS_7_ctrl_serveStealReq_ready,
	io_connVAS_7_data_qOutTask_ready,
	io_connVAS_7_data_qOutTask_valid,
	io_connVAS_7_data_qOutTask_bits,
	io_connVAS_8_ctrl_serveStealReq_valid,
	io_connVAS_8_ctrl_serveStealReq_ready,
	io_connVAS_8_data_qOutTask_ready,
	io_connVAS_8_data_qOutTask_valid,
	io_connVAS_8_data_qOutTask_bits,
	io_connVAS_9_ctrl_serveStealReq_valid,
	io_connVAS_9_ctrl_serveStealReq_ready,
	io_connVAS_9_data_qOutTask_ready,
	io_connVAS_9_data_qOutTask_valid,
	io_connVAS_9_data_qOutTask_bits,
	io_connVAS_10_ctrl_serveStealReq_valid,
	io_connVAS_10_ctrl_serveStealReq_ready,
	io_connVAS_10_data_qOutTask_ready,
	io_connVAS_10_data_qOutTask_valid,
	io_connVAS_10_data_qOutTask_bits,
	io_connVAS_11_ctrl_serveStealReq_valid,
	io_connVAS_11_ctrl_serveStealReq_ready,
	io_connVAS_11_data_qOutTask_ready,
	io_connVAS_11_data_qOutTask_valid,
	io_connVAS_11_data_qOutTask_bits,
	io_connVAS_12_ctrl_serveStealReq_valid,
	io_connVAS_12_ctrl_serveStealReq_ready,
	io_connVAS_12_data_qOutTask_ready,
	io_connVAS_12_data_qOutTask_valid,
	io_connVAS_12_data_qOutTask_bits,
	io_connVAS_13_ctrl_serveStealReq_valid,
	io_connVAS_13_ctrl_serveStealReq_ready,
	io_connVAS_13_data_qOutTask_ready,
	io_connVAS_13_data_qOutTask_valid,
	io_connVAS_13_data_qOutTask_bits,
	io_connVAS_14_ctrl_serveStealReq_valid,
	io_connVAS_14_ctrl_serveStealReq_ready,
	io_connVAS_14_data_qOutTask_ready,
	io_connVAS_14_data_qOutTask_valid,
	io_connVAS_14_data_qOutTask_bits,
	io_connVAS_15_ctrl_serveStealReq_valid,
	io_connVAS_15_ctrl_serveStealReq_ready,
	io_connVAS_15_data_qOutTask_ready,
	io_connVAS_15_data_qOutTask_valid,
	io_connVAS_15_data_qOutTask_bits,
	io_ntwDataUnitOccupancyVSS_0
);
	input clock;
	input reset;
	input io_connPE_0_pop_ready;
	output wire io_connPE_0_pop_valid;
	input io_connPE_1_pop_ready;
	output wire io_connPE_1_pop_valid;
	input io_connPE_2_pop_ready;
	output wire io_connPE_2_pop_valid;
	input io_connPE_3_pop_ready;
	output wire io_connPE_3_pop_valid;
	input io_connPE_4_pop_ready;
	output wire io_connPE_4_pop_valid;
	input io_connPE_5_pop_ready;
	output wire io_connPE_5_pop_valid;
	input io_connPE_6_pop_ready;
	output wire io_connPE_6_pop_valid;
	input io_connPE_7_pop_ready;
	output wire io_connPE_7_pop_valid;
	input io_connPE_8_pop_ready;
	output wire io_connPE_8_pop_valid;
	input io_connPE_9_pop_ready;
	output wire io_connPE_9_pop_valid;
	input io_connPE_10_pop_ready;
	output wire io_connPE_10_pop_valid;
	input io_connPE_11_pop_ready;
	output wire io_connPE_11_pop_valid;
	input io_connPE_12_pop_ready;
	output wire io_connPE_12_pop_valid;
	input io_connPE_13_pop_ready;
	output wire io_connPE_13_pop_valid;
	input io_connPE_14_pop_ready;
	output wire io_connPE_14_pop_valid;
	input io_connPE_15_pop_ready;
	output wire io_connPE_15_pop_valid;
	input io_connVSS_0_ctrl_serveStealReq_valid;
	output wire io_connVSS_0_ctrl_serveStealReq_ready;
	input io_connVSS_0_data_availableTask_ready;
	output wire io_connVSS_0_data_availableTask_valid;
	output wire [127:0] io_connVSS_0_data_availableTask_bits;
	output wire io_connVSS_0_data_qOutTask_ready;
	input io_connVSS_0_data_qOutTask_valid;
	input [127:0] io_connVSS_0_data_qOutTask_bits;
	input io_connVAS_0_ctrl_serveStealReq_valid;
	output wire io_connVAS_0_ctrl_serveStealReq_ready;
	output wire io_connVAS_0_data_qOutTask_ready;
	input io_connVAS_0_data_qOutTask_valid;
	input [127:0] io_connVAS_0_data_qOutTask_bits;
	input io_connVAS_1_ctrl_serveStealReq_valid;
	output wire io_connVAS_1_ctrl_serveStealReq_ready;
	output wire io_connVAS_1_data_qOutTask_ready;
	input io_connVAS_1_data_qOutTask_valid;
	input [127:0] io_connVAS_1_data_qOutTask_bits;
	input io_connVAS_2_ctrl_serveStealReq_valid;
	output wire io_connVAS_2_ctrl_serveStealReq_ready;
	output wire io_connVAS_2_data_qOutTask_ready;
	input io_connVAS_2_data_qOutTask_valid;
	input [127:0] io_connVAS_2_data_qOutTask_bits;
	input io_connVAS_3_ctrl_serveStealReq_valid;
	output wire io_connVAS_3_ctrl_serveStealReq_ready;
	output wire io_connVAS_3_data_qOutTask_ready;
	input io_connVAS_3_data_qOutTask_valid;
	input [127:0] io_connVAS_3_data_qOutTask_bits;
	input io_connVAS_4_ctrl_serveStealReq_valid;
	output wire io_connVAS_4_ctrl_serveStealReq_ready;
	output wire io_connVAS_4_data_qOutTask_ready;
	input io_connVAS_4_data_qOutTask_valid;
	input [127:0] io_connVAS_4_data_qOutTask_bits;
	input io_connVAS_5_ctrl_serveStealReq_valid;
	output wire io_connVAS_5_ctrl_serveStealReq_ready;
	output wire io_connVAS_5_data_qOutTask_ready;
	input io_connVAS_5_data_qOutTask_valid;
	input [127:0] io_connVAS_5_data_qOutTask_bits;
	input io_connVAS_6_ctrl_serveStealReq_valid;
	output wire io_connVAS_6_ctrl_serveStealReq_ready;
	output wire io_connVAS_6_data_qOutTask_ready;
	input io_connVAS_6_data_qOutTask_valid;
	input [127:0] io_connVAS_6_data_qOutTask_bits;
	input io_connVAS_7_ctrl_serveStealReq_valid;
	output wire io_connVAS_7_ctrl_serveStealReq_ready;
	output wire io_connVAS_7_data_qOutTask_ready;
	input io_connVAS_7_data_qOutTask_valid;
	input [127:0] io_connVAS_7_data_qOutTask_bits;
	input io_connVAS_8_ctrl_serveStealReq_valid;
	output wire io_connVAS_8_ctrl_serveStealReq_ready;
	output wire io_connVAS_8_data_qOutTask_ready;
	input io_connVAS_8_data_qOutTask_valid;
	input [127:0] io_connVAS_8_data_qOutTask_bits;
	input io_connVAS_9_ctrl_serveStealReq_valid;
	output wire io_connVAS_9_ctrl_serveStealReq_ready;
	output wire io_connVAS_9_data_qOutTask_ready;
	input io_connVAS_9_data_qOutTask_valid;
	input [127:0] io_connVAS_9_data_qOutTask_bits;
	input io_connVAS_10_ctrl_serveStealReq_valid;
	output wire io_connVAS_10_ctrl_serveStealReq_ready;
	output wire io_connVAS_10_data_qOutTask_ready;
	input io_connVAS_10_data_qOutTask_valid;
	input [127:0] io_connVAS_10_data_qOutTask_bits;
	input io_connVAS_11_ctrl_serveStealReq_valid;
	output wire io_connVAS_11_ctrl_serveStealReq_ready;
	output wire io_connVAS_11_data_qOutTask_ready;
	input io_connVAS_11_data_qOutTask_valid;
	input [127:0] io_connVAS_11_data_qOutTask_bits;
	input io_connVAS_12_ctrl_serveStealReq_valid;
	output wire io_connVAS_12_ctrl_serveStealReq_ready;
	output wire io_connVAS_12_data_qOutTask_ready;
	input io_connVAS_12_data_qOutTask_valid;
	input [127:0] io_connVAS_12_data_qOutTask_bits;
	input io_connVAS_13_ctrl_serveStealReq_valid;
	output wire io_connVAS_13_ctrl_serveStealReq_ready;
	output wire io_connVAS_13_data_qOutTask_ready;
	input io_connVAS_13_data_qOutTask_valid;
	input [127:0] io_connVAS_13_data_qOutTask_bits;
	input io_connVAS_14_ctrl_serveStealReq_valid;
	output wire io_connVAS_14_ctrl_serveStealReq_ready;
	output wire io_connVAS_14_data_qOutTask_ready;
	input io_connVAS_14_data_qOutTask_valid;
	input [127:0] io_connVAS_14_data_qOutTask_bits;
	input io_connVAS_15_ctrl_serveStealReq_valid;
	output wire io_connVAS_15_ctrl_serveStealReq_ready;
	output wire io_connVAS_15_data_qOutTask_ready;
	input io_connVAS_15_data_qOutTask_valid;
	input [127:0] io_connVAS_15_data_qOutTask_bits;
	output wire io_ntwDataUnitOccupancyVSS_0;
	wire [8:0] _taskQueues_15_io_connVec_1_currLength;
	wire _taskQueues_15_io_connVec_1_push_ready;
	wire _taskQueues_15_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_15_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_14_io_connVec_1_currLength;
	wire _taskQueues_14_io_connVec_1_push_ready;
	wire _taskQueues_14_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_14_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_13_io_connVec_1_currLength;
	wire _taskQueues_13_io_connVec_1_push_ready;
	wire _taskQueues_13_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_13_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_12_io_connVec_1_currLength;
	wire _taskQueues_12_io_connVec_1_push_ready;
	wire _taskQueues_12_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_12_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_11_io_connVec_1_currLength;
	wire _taskQueues_11_io_connVec_1_push_ready;
	wire _taskQueues_11_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_11_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_10_io_connVec_1_currLength;
	wire _taskQueues_10_io_connVec_1_push_ready;
	wire _taskQueues_10_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_10_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_9_io_connVec_1_currLength;
	wire _taskQueues_9_io_connVec_1_push_ready;
	wire _taskQueues_9_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_9_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_8_io_connVec_1_currLength;
	wire _taskQueues_8_io_connVec_1_push_ready;
	wire _taskQueues_8_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_8_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_7_io_connVec_1_currLength;
	wire _taskQueues_7_io_connVec_1_push_ready;
	wire _taskQueues_7_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_7_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_6_io_connVec_1_currLength;
	wire _taskQueues_6_io_connVec_1_push_ready;
	wire _taskQueues_6_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_6_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_5_io_connVec_1_currLength;
	wire _taskQueues_5_io_connVec_1_push_ready;
	wire _taskQueues_5_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_5_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_4_io_connVec_1_currLength;
	wire _taskQueues_4_io_connVec_1_push_ready;
	wire _taskQueues_4_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_4_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_3_io_connVec_1_currLength;
	wire _taskQueues_3_io_connVec_1_push_ready;
	wire _taskQueues_3_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_3_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_2_io_connVec_1_currLength;
	wire _taskQueues_2_io_connVec_1_push_ready;
	wire _taskQueues_2_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_2_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_1_io_connVec_1_currLength;
	wire _taskQueues_1_io_connVec_1_push_ready;
	wire _taskQueues_1_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_1_io_connVec_1_pop_bits;
	wire [8:0] _taskQueues_0_io_connVec_1_currLength;
	wire _taskQueues_0_io_connVec_1_push_ready;
	wire _taskQueues_0_io_connVec_1_pop_valid;
	wire [127:0] _taskQueues_0_io_connVec_1_pop_bits;
	wire _stealServers_15_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_15_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_15_io_connNetwork_data_availableTask_ready;
	wire _stealServers_15_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_15_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_15_io_connQ_push_valid;
	wire [127:0] _stealServers_15_io_connQ_push_bits;
	wire _stealServers_15_io_connQ_pop_ready;
	wire _stealServers_14_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_14_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_14_io_connNetwork_data_availableTask_ready;
	wire _stealServers_14_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_14_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_14_io_connQ_push_valid;
	wire [127:0] _stealServers_14_io_connQ_push_bits;
	wire _stealServers_14_io_connQ_pop_ready;
	wire _stealServers_13_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_13_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_13_io_connNetwork_data_availableTask_ready;
	wire _stealServers_13_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_13_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_13_io_connQ_push_valid;
	wire [127:0] _stealServers_13_io_connQ_push_bits;
	wire _stealServers_13_io_connQ_pop_ready;
	wire _stealServers_12_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_12_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_12_io_connNetwork_data_availableTask_ready;
	wire _stealServers_12_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_12_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_12_io_connQ_push_valid;
	wire [127:0] _stealServers_12_io_connQ_push_bits;
	wire _stealServers_12_io_connQ_pop_ready;
	wire _stealServers_11_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_11_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_11_io_connNetwork_data_availableTask_ready;
	wire _stealServers_11_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_11_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_11_io_connQ_push_valid;
	wire [127:0] _stealServers_11_io_connQ_push_bits;
	wire _stealServers_11_io_connQ_pop_ready;
	wire _stealServers_10_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_10_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_10_io_connNetwork_data_availableTask_ready;
	wire _stealServers_10_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_10_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_10_io_connQ_push_valid;
	wire [127:0] _stealServers_10_io_connQ_push_bits;
	wire _stealServers_10_io_connQ_pop_ready;
	wire _stealServers_9_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_9_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_9_io_connNetwork_data_availableTask_ready;
	wire _stealServers_9_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_9_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_9_io_connQ_push_valid;
	wire [127:0] _stealServers_9_io_connQ_push_bits;
	wire _stealServers_9_io_connQ_pop_ready;
	wire _stealServers_8_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_8_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_8_io_connNetwork_data_availableTask_ready;
	wire _stealServers_8_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_8_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_8_io_connQ_push_valid;
	wire [127:0] _stealServers_8_io_connQ_push_bits;
	wire _stealServers_8_io_connQ_pop_ready;
	wire _stealServers_7_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_7_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_7_io_connNetwork_data_availableTask_ready;
	wire _stealServers_7_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_7_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_7_io_connQ_push_valid;
	wire [127:0] _stealServers_7_io_connQ_push_bits;
	wire _stealServers_7_io_connQ_pop_ready;
	wire _stealServers_6_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_6_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_6_io_connNetwork_data_availableTask_ready;
	wire _stealServers_6_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_6_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_6_io_connQ_push_valid;
	wire [127:0] _stealServers_6_io_connQ_push_bits;
	wire _stealServers_6_io_connQ_pop_ready;
	wire _stealServers_5_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_5_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_5_io_connNetwork_data_availableTask_ready;
	wire _stealServers_5_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_5_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_5_io_connQ_push_valid;
	wire [127:0] _stealServers_5_io_connQ_push_bits;
	wire _stealServers_5_io_connQ_pop_ready;
	wire _stealServers_4_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_4_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_4_io_connNetwork_data_availableTask_ready;
	wire _stealServers_4_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_4_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_4_io_connQ_push_valid;
	wire [127:0] _stealServers_4_io_connQ_push_bits;
	wire _stealServers_4_io_connQ_pop_ready;
	wire _stealServers_3_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_3_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_3_io_connNetwork_data_availableTask_ready;
	wire _stealServers_3_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_3_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_3_io_connQ_push_valid;
	wire [127:0] _stealServers_3_io_connQ_push_bits;
	wire _stealServers_3_io_connQ_pop_ready;
	wire _stealServers_2_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_2_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_2_io_connNetwork_data_availableTask_ready;
	wire _stealServers_2_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_2_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_2_io_connQ_push_valid;
	wire [127:0] _stealServers_2_io_connQ_push_bits;
	wire _stealServers_2_io_connQ_pop_ready;
	wire _stealServers_1_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_1_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_1_io_connNetwork_data_availableTask_ready;
	wire _stealServers_1_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_1_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_1_io_connQ_push_valid;
	wire [127:0] _stealServers_1_io_connQ_push_bits;
	wire _stealServers_1_io_connQ_pop_ready;
	wire _stealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _stealServers_0_io_connNetwork_ctrl_stealReq_valid;
	wire _stealServers_0_io_connNetwork_data_availableTask_ready;
	wire _stealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _stealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _stealServers_0_io_connQ_push_valid;
	wire [127:0] _stealServers_0_io_connQ_push_bits;
	wire _stealServers_0_io_connQ_pop_ready;
	wire _stealNet_io_connSS_17_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_17_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_17_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_17_data_availableTask_bits;
	wire _stealNet_io_connSS_17_data_qOutTask_ready;
	wire _stealNet_io_connSS_18_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_18_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_18_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_18_data_availableTask_bits;
	wire _stealNet_io_connSS_18_data_qOutTask_ready;
	wire _stealNet_io_connSS_19_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_19_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_19_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_19_data_availableTask_bits;
	wire _stealNet_io_connSS_19_data_qOutTask_ready;
	wire _stealNet_io_connSS_20_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_20_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_20_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_20_data_availableTask_bits;
	wire _stealNet_io_connSS_20_data_qOutTask_ready;
	wire _stealNet_io_connSS_21_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_21_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_21_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_21_data_availableTask_bits;
	wire _stealNet_io_connSS_21_data_qOutTask_ready;
	wire _stealNet_io_connSS_22_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_22_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_22_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_22_data_availableTask_bits;
	wire _stealNet_io_connSS_22_data_qOutTask_ready;
	wire _stealNet_io_connSS_23_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_23_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_23_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_23_data_availableTask_bits;
	wire _stealNet_io_connSS_23_data_qOutTask_ready;
	wire _stealNet_io_connSS_24_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_24_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_24_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_24_data_availableTask_bits;
	wire _stealNet_io_connSS_24_data_qOutTask_ready;
	wire _stealNet_io_connSS_25_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_25_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_25_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_25_data_availableTask_bits;
	wire _stealNet_io_connSS_25_data_qOutTask_ready;
	wire _stealNet_io_connSS_26_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_26_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_26_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_26_data_availableTask_bits;
	wire _stealNet_io_connSS_26_data_qOutTask_ready;
	wire _stealNet_io_connSS_27_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_27_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_27_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_27_data_availableTask_bits;
	wire _stealNet_io_connSS_27_data_qOutTask_ready;
	wire _stealNet_io_connSS_28_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_28_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_28_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_28_data_availableTask_bits;
	wire _stealNet_io_connSS_28_data_qOutTask_ready;
	wire _stealNet_io_connSS_29_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_29_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_29_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_29_data_availableTask_bits;
	wire _stealNet_io_connSS_29_data_qOutTask_ready;
	wire _stealNet_io_connSS_30_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_30_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_30_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_30_data_availableTask_bits;
	wire _stealNet_io_connSS_30_data_qOutTask_ready;
	wire _stealNet_io_connSS_31_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_31_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_31_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_31_data_availableTask_bits;
	wire _stealNet_io_connSS_31_data_qOutTask_ready;
	wire _stealNet_io_connSS_32_ctrl_serveStealReq_ready;
	wire _stealNet_io_connSS_32_ctrl_stealReq_ready;
	wire _stealNet_io_connSS_32_data_availableTask_valid;
	wire [127:0] _stealNet_io_connSS_32_data_availableTask_bits;
	wire _stealNet_io_connSS_32_data_qOutTask_ready;
	SchedulerNetwork_1 stealNet(
		.clock(clock),
		.reset(reset),
		.io_connSS_0_ctrl_serveStealReq_valid(io_connVAS_0_ctrl_serveStealReq_valid),
		.io_connSS_0_ctrl_serveStealReq_ready(io_connVAS_0_ctrl_serveStealReq_ready),
		.io_connSS_0_data_availableTask_ready(io_connVSS_0_data_availableTask_ready),
		.io_connSS_0_data_availableTask_valid(io_connVSS_0_data_availableTask_valid),
		.io_connSS_0_data_availableTask_bits(io_connVSS_0_data_availableTask_bits),
		.io_connSS_0_data_qOutTask_ready(io_connVSS_0_data_qOutTask_ready),
		.io_connSS_0_data_qOutTask_valid(io_connVSS_0_data_qOutTask_valid),
		.io_connSS_0_data_qOutTask_bits(io_connVSS_0_data_qOutTask_bits),
		.io_connSS_1_ctrl_serveStealReq_valid(io_connVAS_1_ctrl_serveStealReq_valid),
		.io_connSS_1_ctrl_serveStealReq_ready(io_connVAS_1_ctrl_serveStealReq_ready),
		.io_connSS_1_data_qOutTask_ready(io_connVAS_0_data_qOutTask_ready),
		.io_connSS_1_data_qOutTask_valid(io_connVAS_0_data_qOutTask_valid),
		.io_connSS_1_data_qOutTask_bits(io_connVAS_0_data_qOutTask_bits),
		.io_connSS_2_ctrl_serveStealReq_valid(io_connVAS_2_ctrl_serveStealReq_valid),
		.io_connSS_2_ctrl_serveStealReq_ready(io_connVAS_2_ctrl_serveStealReq_ready),
		.io_connSS_2_data_qOutTask_ready(io_connVAS_1_data_qOutTask_ready),
		.io_connSS_2_data_qOutTask_valid(io_connVAS_1_data_qOutTask_valid),
		.io_connSS_2_data_qOutTask_bits(io_connVAS_1_data_qOutTask_bits),
		.io_connSS_3_ctrl_serveStealReq_valid(io_connVAS_3_ctrl_serveStealReq_valid),
		.io_connSS_3_ctrl_serveStealReq_ready(io_connVAS_3_ctrl_serveStealReq_ready),
		.io_connSS_3_data_qOutTask_ready(io_connVAS_2_data_qOutTask_ready),
		.io_connSS_3_data_qOutTask_valid(io_connVAS_2_data_qOutTask_valid),
		.io_connSS_3_data_qOutTask_bits(io_connVAS_2_data_qOutTask_bits),
		.io_connSS_4_ctrl_serveStealReq_valid(io_connVAS_4_ctrl_serveStealReq_valid),
		.io_connSS_4_ctrl_serveStealReq_ready(io_connVAS_4_ctrl_serveStealReq_ready),
		.io_connSS_4_data_qOutTask_ready(io_connVAS_3_data_qOutTask_ready),
		.io_connSS_4_data_qOutTask_valid(io_connVAS_3_data_qOutTask_valid),
		.io_connSS_4_data_qOutTask_bits(io_connVAS_3_data_qOutTask_bits),
		.io_connSS_5_ctrl_serveStealReq_valid(io_connVAS_5_ctrl_serveStealReq_valid),
		.io_connSS_5_ctrl_serveStealReq_ready(io_connVAS_5_ctrl_serveStealReq_ready),
		.io_connSS_5_data_qOutTask_ready(io_connVAS_4_data_qOutTask_ready),
		.io_connSS_5_data_qOutTask_valid(io_connVAS_4_data_qOutTask_valid),
		.io_connSS_5_data_qOutTask_bits(io_connVAS_4_data_qOutTask_bits),
		.io_connSS_6_ctrl_serveStealReq_valid(io_connVAS_6_ctrl_serveStealReq_valid),
		.io_connSS_6_ctrl_serveStealReq_ready(io_connVAS_6_ctrl_serveStealReq_ready),
		.io_connSS_6_data_qOutTask_ready(io_connVAS_5_data_qOutTask_ready),
		.io_connSS_6_data_qOutTask_valid(io_connVAS_5_data_qOutTask_valid),
		.io_connSS_6_data_qOutTask_bits(io_connVAS_5_data_qOutTask_bits),
		.io_connSS_7_ctrl_serveStealReq_valid(io_connVAS_7_ctrl_serveStealReq_valid),
		.io_connSS_7_ctrl_serveStealReq_ready(io_connVAS_7_ctrl_serveStealReq_ready),
		.io_connSS_7_data_qOutTask_ready(io_connVAS_6_data_qOutTask_ready),
		.io_connSS_7_data_qOutTask_valid(io_connVAS_6_data_qOutTask_valid),
		.io_connSS_7_data_qOutTask_bits(io_connVAS_6_data_qOutTask_bits),
		.io_connSS_8_ctrl_serveStealReq_valid(io_connVAS_8_ctrl_serveStealReq_valid),
		.io_connSS_8_ctrl_serveStealReq_ready(io_connVAS_8_ctrl_serveStealReq_ready),
		.io_connSS_8_data_qOutTask_ready(io_connVAS_7_data_qOutTask_ready),
		.io_connSS_8_data_qOutTask_valid(io_connVAS_7_data_qOutTask_valid),
		.io_connSS_8_data_qOutTask_bits(io_connVAS_7_data_qOutTask_bits),
		.io_connSS_9_ctrl_serveStealReq_valid(io_connVAS_9_ctrl_serveStealReq_valid),
		.io_connSS_9_ctrl_serveStealReq_ready(io_connVAS_9_ctrl_serveStealReq_ready),
		.io_connSS_9_data_qOutTask_ready(io_connVAS_8_data_qOutTask_ready),
		.io_connSS_9_data_qOutTask_valid(io_connVAS_8_data_qOutTask_valid),
		.io_connSS_9_data_qOutTask_bits(io_connVAS_8_data_qOutTask_bits),
		.io_connSS_10_ctrl_serveStealReq_valid(io_connVAS_10_ctrl_serveStealReq_valid),
		.io_connSS_10_ctrl_serveStealReq_ready(io_connVAS_10_ctrl_serveStealReq_ready),
		.io_connSS_10_data_qOutTask_ready(io_connVAS_9_data_qOutTask_ready),
		.io_connSS_10_data_qOutTask_valid(io_connVAS_9_data_qOutTask_valid),
		.io_connSS_10_data_qOutTask_bits(io_connVAS_9_data_qOutTask_bits),
		.io_connSS_11_ctrl_serveStealReq_valid(io_connVAS_11_ctrl_serveStealReq_valid),
		.io_connSS_11_ctrl_serveStealReq_ready(io_connVAS_11_ctrl_serveStealReq_ready),
		.io_connSS_11_data_qOutTask_ready(io_connVAS_10_data_qOutTask_ready),
		.io_connSS_11_data_qOutTask_valid(io_connVAS_10_data_qOutTask_valid),
		.io_connSS_11_data_qOutTask_bits(io_connVAS_10_data_qOutTask_bits),
		.io_connSS_12_ctrl_serveStealReq_valid(io_connVAS_12_ctrl_serveStealReq_valid),
		.io_connSS_12_ctrl_serveStealReq_ready(io_connVAS_12_ctrl_serveStealReq_ready),
		.io_connSS_12_data_qOutTask_ready(io_connVAS_11_data_qOutTask_ready),
		.io_connSS_12_data_qOutTask_valid(io_connVAS_11_data_qOutTask_valid),
		.io_connSS_12_data_qOutTask_bits(io_connVAS_11_data_qOutTask_bits),
		.io_connSS_13_ctrl_serveStealReq_valid(io_connVAS_13_ctrl_serveStealReq_valid),
		.io_connSS_13_ctrl_serveStealReq_ready(io_connVAS_13_ctrl_serveStealReq_ready),
		.io_connSS_13_data_qOutTask_ready(io_connVAS_12_data_qOutTask_ready),
		.io_connSS_13_data_qOutTask_valid(io_connVAS_12_data_qOutTask_valid),
		.io_connSS_13_data_qOutTask_bits(io_connVAS_12_data_qOutTask_bits),
		.io_connSS_14_ctrl_serveStealReq_valid(io_connVAS_14_ctrl_serveStealReq_valid),
		.io_connSS_14_ctrl_serveStealReq_ready(io_connVAS_14_ctrl_serveStealReq_ready),
		.io_connSS_14_data_qOutTask_ready(io_connVAS_13_data_qOutTask_ready),
		.io_connSS_14_data_qOutTask_valid(io_connVAS_13_data_qOutTask_valid),
		.io_connSS_14_data_qOutTask_bits(io_connVAS_13_data_qOutTask_bits),
		.io_connSS_15_ctrl_serveStealReq_valid(io_connVAS_15_ctrl_serveStealReq_valid),
		.io_connSS_15_ctrl_serveStealReq_ready(io_connVAS_15_ctrl_serveStealReq_ready),
		.io_connSS_15_data_qOutTask_ready(io_connVAS_14_data_qOutTask_ready),
		.io_connSS_15_data_qOutTask_valid(io_connVAS_14_data_qOutTask_valid),
		.io_connSS_15_data_qOutTask_bits(io_connVAS_14_data_qOutTask_bits),
		.io_connSS_16_ctrl_serveStealReq_valid(io_connVSS_0_ctrl_serveStealReq_valid),
		.io_connSS_16_ctrl_serveStealReq_ready(io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connSS_16_data_qOutTask_ready(io_connVAS_15_data_qOutTask_ready),
		.io_connSS_16_data_qOutTask_valid(io_connVAS_15_data_qOutTask_valid),
		.io_connSS_16_data_qOutTask_bits(io_connVAS_15_data_qOutTask_bits),
		.io_connSS_17_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_17_ctrl_serveStealReq_ready(_stealNet_io_connSS_17_ctrl_serveStealReq_ready),
		.io_connSS_17_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_17_ctrl_stealReq_ready(_stealNet_io_connSS_17_ctrl_stealReq_ready),
		.io_connSS_17_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connSS_17_data_availableTask_valid(_stealNet_io_connSS_17_data_availableTask_valid),
		.io_connSS_17_data_availableTask_bits(_stealNet_io_connSS_17_data_availableTask_bits),
		.io_connSS_17_data_qOutTask_ready(_stealNet_io_connSS_17_data_qOutTask_ready),
		.io_connSS_17_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connSS_17_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connSS_18_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_18_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connSS_18_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_18_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connSS_18_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connSS_18_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connSS_18_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connSS_18_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connSS_18_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connSS_18_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connSS_19_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_19_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connSS_19_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_19_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connSS_19_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connSS_19_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connSS_19_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connSS_19_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connSS_19_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connSS_19_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connSS_20_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_20_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connSS_20_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_20_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connSS_20_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connSS_20_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connSS_20_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connSS_20_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connSS_20_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connSS_20_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connSS_21_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_21_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connSS_21_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_21_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connSS_21_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connSS_21_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connSS_21_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connSS_21_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connSS_21_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connSS_21_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connSS_22_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_22_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connSS_22_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_22_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connSS_22_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connSS_22_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connSS_22_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connSS_22_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connSS_22_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connSS_22_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connSS_23_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_23_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connSS_23_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_23_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connSS_23_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connSS_23_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connSS_23_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connSS_23_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connSS_23_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connSS_23_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connSS_24_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_24_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connSS_24_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_24_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connSS_24_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connSS_24_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connSS_24_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connSS_24_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connSS_24_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connSS_24_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connSS_25_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_25_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connSS_25_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_25_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connSS_25_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connSS_25_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connSS_25_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connSS_25_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connSS_25_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connSS_25_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connSS_26_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_26_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connSS_26_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_26_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connSS_26_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connSS_26_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connSS_26_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connSS_26_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connSS_26_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connSS_26_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connSS_27_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_27_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connSS_27_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_27_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connSS_27_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connSS_27_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connSS_27_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connSS_27_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connSS_27_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connSS_27_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connSS_28_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_28_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connSS_28_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_28_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connSS_28_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connSS_28_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connSS_28_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connSS_28_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connSS_28_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connSS_28_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connSS_29_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_29_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connSS_29_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_29_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connSS_29_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connSS_29_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connSS_29_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connSS_29_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connSS_29_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connSS_29_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connSS_30_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_30_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connSS_30_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_30_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connSS_30_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connSS_30_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connSS_30_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connSS_30_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connSS_30_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connSS_30_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connSS_31_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_31_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connSS_31_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_31_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connSS_31_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connSS_31_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connSS_31_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connSS_31_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connSS_31_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connSS_31_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connSS_32_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connSS_32_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connSS_32_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connSS_32_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connSS_32_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connSS_32_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connSS_32_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connSS_32_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connSS_32_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connSS_32_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerClient_64 stealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_17_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_0_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_17_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_17_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_17_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_17_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_0_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_1_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_18_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_1_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_18_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_1_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_18_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_18_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_18_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_1_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_1_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_1_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_2(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_2_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_19_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_2_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_19_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_2_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_19_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_19_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_19_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_2_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_2_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_2_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_3(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_3_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_20_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_3_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_20_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_3_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_20_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_20_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_20_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_3_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_3_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_3_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_4(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_4_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_21_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_4_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_21_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_4_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_21_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_21_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_21_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_4_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_4_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_4_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_5(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_5_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_22_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_5_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_22_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_5_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_22_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_22_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_22_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_5_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_5_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_5_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_6(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_6_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_23_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_6_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_23_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_6_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_23_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_23_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_23_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_6_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_6_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_6_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_7(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_7_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_24_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_7_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_24_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_7_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_24_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_24_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_24_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_7_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_7_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_7_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_8(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_8_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_25_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_8_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_25_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_8_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_25_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_25_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_25_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_8_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_8_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_8_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_9(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_9_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_26_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_9_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_26_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_9_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_26_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_26_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_26_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_9_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_9_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_9_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_10(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_10_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_27_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_10_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_27_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_10_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_27_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_27_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_27_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_10_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_10_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_10_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_11(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_11_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_28_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_11_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_28_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_11_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_28_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_28_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_28_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_11_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_11_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_11_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_12(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_12_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_29_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_12_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_29_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_12_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_29_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_29_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_29_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_12_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_12_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_12_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_13(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_13_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_30_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_13_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_30_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_13_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_30_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_30_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_30_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_13_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_13_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_13_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_14(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_14_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_31_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_14_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_31_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_14_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_31_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_31_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_31_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_14_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_14_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_14_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	SchedulerClient_64 stealServers_15(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_stealServers_15_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNet_io_connSS_32_ctrl_serveStealReq_ready),
		.io_connNetwork_ctrl_stealReq_valid(_stealServers_15_io_connNetwork_ctrl_stealReq_valid),
		.io_connNetwork_ctrl_stealReq_ready(_stealNet_io_connSS_32_ctrl_stealReq_ready),
		.io_connNetwork_data_availableTask_ready(_stealServers_15_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNet_io_connSS_32_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNet_io_connSS_32_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNet_io_connSS_32_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_stealServers_15_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_stealServers_15_io_connNetwork_data_qOutTask_bits),
		.io_connQ_currLength(_taskQueues_15_io_connVec_1_currLength[7:0]),
		.io_connQ_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connQ_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connQ_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connQ_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connQ_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connQ_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_0(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_0_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_0_pop_valid),
		.io_connVec_1_currLength(_taskQueues_0_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_0_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_0_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_0_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_0_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_0_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_0_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_1(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_1_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_1_pop_valid),
		.io_connVec_1_currLength(_taskQueues_1_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_1_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_1_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_1_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_1_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_1_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_1_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_2(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_2_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_2_pop_valid),
		.io_connVec_1_currLength(_taskQueues_2_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_2_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_2_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_2_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_2_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_2_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_2_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_3(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_3_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_3_pop_valid),
		.io_connVec_1_currLength(_taskQueues_3_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_3_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_3_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_3_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_3_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_3_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_3_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_4(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_4_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_4_pop_valid),
		.io_connVec_1_currLength(_taskQueues_4_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_4_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_4_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_4_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_4_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_4_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_4_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_5(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_5_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_5_pop_valid),
		.io_connVec_1_currLength(_taskQueues_5_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_5_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_5_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_5_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_5_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_5_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_5_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_6(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_6_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_6_pop_valid),
		.io_connVec_1_currLength(_taskQueues_6_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_6_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_6_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_6_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_6_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_6_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_6_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_7(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_7_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_7_pop_valid),
		.io_connVec_1_currLength(_taskQueues_7_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_7_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_7_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_7_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_7_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_7_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_7_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_8(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_8_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_8_pop_valid),
		.io_connVec_1_currLength(_taskQueues_8_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_8_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_8_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_8_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_8_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_8_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_8_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_9(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_9_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_9_pop_valid),
		.io_connVec_1_currLength(_taskQueues_9_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_9_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_9_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_9_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_9_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_9_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_9_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_10(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_10_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_10_pop_valid),
		.io_connVec_1_currLength(_taskQueues_10_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_10_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_10_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_10_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_10_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_10_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_10_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_11(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_11_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_11_pop_valid),
		.io_connVec_1_currLength(_taskQueues_11_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_11_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_11_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_11_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_11_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_11_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_11_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_12(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_12_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_12_pop_valid),
		.io_connVec_1_currLength(_taskQueues_12_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_12_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_12_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_12_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_12_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_12_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_12_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_13(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_13_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_13_pop_valid),
		.io_connVec_1_currLength(_taskQueues_13_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_13_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_13_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_13_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_13_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_13_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_13_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_14(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_14_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_14_pop_valid),
		.io_connVec_1_currLength(_taskQueues_14_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_14_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_14_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_14_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_14_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_14_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_14_io_connVec_1_pop_bits)
	);
	hw_deque_64 taskQueues_15(
		.clock(clock),
		.reset(reset),
		.io_connVec_0_pop_ready(io_connPE_15_pop_ready),
		.io_connVec_0_pop_valid(io_connPE_15_pop_valid),
		.io_connVec_1_currLength(_taskQueues_15_io_connVec_1_currLength),
		.io_connVec_1_push_ready(_taskQueues_15_io_connVec_1_push_ready),
		.io_connVec_1_push_valid(_stealServers_15_io_connQ_push_valid),
		.io_connVec_1_push_bits(_stealServers_15_io_connQ_push_bits),
		.io_connVec_1_pop_ready(_stealServers_15_io_connQ_pop_ready),
		.io_connVec_1_pop_valid(_taskQueues_15_io_connVec_1_pop_valid),
		.io_connVec_1_pop_bits(_taskQueues_15_io_connVec_1_pop_bits)
	);
endmodule
module Queue1_UInt_1 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_bits,
	io_count
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [127:0] io_enq_bits;
	input io_deq_ready;
	output wire [127:0] io_deq_bits;
	output wire io_count;
	reg [127:0] ram;
	reg full;
	always @(posedge clock) begin : sv2v_autoblock_1
		reg do_enq;
		do_enq = ~full & io_enq_valid;
		if (do_enq)
			ram <= io_enq_bits;
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == (io_deq_ready & full)))
			full <= do_enq;
	end
	assign io_enq_ready = ~full;
	assign io_deq_bits = ram;
	assign io_count = full;
endmodule
module SchedulerServer_1 (
	clock,
	reset,
	io_connNetwork_ctrl_serveStealReq_valid,
	io_connNetwork_ctrl_serveStealReq_ready,
	io_connNetwork_data_availableTask_ready,
	io_connNetwork_data_availableTask_valid,
	io_connNetwork_data_availableTask_bits,
	io_connNetwork_data_qOutTask_ready,
	io_connNetwork_data_qOutTask_valid,
	io_connNetwork_data_qOutTask_bits,
	io_axi_mgmt_ar_ready,
	io_axi_mgmt_ar_valid,
	io_axi_mgmt_ar_bits_addr,
	io_axi_mgmt_ar_bits_prot,
	io_axi_mgmt_r_ready,
	io_axi_mgmt_r_valid,
	io_axi_mgmt_r_bits_data,
	io_axi_mgmt_r_bits_resp,
	io_axi_mgmt_aw_ready,
	io_axi_mgmt_aw_valid,
	io_axi_mgmt_aw_bits_addr,
	io_axi_mgmt_aw_bits_prot,
	io_axi_mgmt_w_ready,
	io_axi_mgmt_w_valid,
	io_axi_mgmt_w_bits_data,
	io_axi_mgmt_w_bits_strb,
	io_axi_mgmt_b_ready,
	io_axi_mgmt_b_valid,
	io_axi_mgmt_b_bits_resp,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_read_burst_len,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_write_last,
	io_ntwDataUnitOccupancy
);
	input clock;
	input reset;
	output wire io_connNetwork_ctrl_serveStealReq_valid;
	input io_connNetwork_ctrl_serveStealReq_ready;
	output wire io_connNetwork_data_availableTask_ready;
	input io_connNetwork_data_availableTask_valid;
	input [127:0] io_connNetwork_data_availableTask_bits;
	input io_connNetwork_data_qOutTask_ready;
	output wire io_connNetwork_data_qOutTask_valid;
	output wire [127:0] io_connNetwork_data_qOutTask_bits;
	output wire io_axi_mgmt_ar_ready;
	input io_axi_mgmt_ar_valid;
	input [5:0] io_axi_mgmt_ar_bits_addr;
	input [2:0] io_axi_mgmt_ar_bits_prot;
	input io_axi_mgmt_r_ready;
	output wire io_axi_mgmt_r_valid;
	output wire [63:0] io_axi_mgmt_r_bits_data;
	output wire [1:0] io_axi_mgmt_r_bits_resp;
	output wire io_axi_mgmt_aw_ready;
	input io_axi_mgmt_aw_valid;
	input [5:0] io_axi_mgmt_aw_bits_addr;
	input [2:0] io_axi_mgmt_aw_bits_prot;
	output wire io_axi_mgmt_w_ready;
	input io_axi_mgmt_w_valid;
	input [63:0] io_axi_mgmt_w_bits_data;
	input [7:0] io_axi_mgmt_w_bits_strb;
	input io_axi_mgmt_b_ready;
	output wire io_axi_mgmt_b_valid;
	output wire [1:0] io_axi_mgmt_b_bits_resp;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [127:0] io_read_data_bits;
	output wire [3:0] io_read_burst_len;
	input io_write_address_ready;
	output wire io_write_address_valid;
	output wire [63:0] io_write_address_bits;
	input io_write_data_ready;
	output wire io_write_data_valid;
	output wire [127:0] io_write_data_bits;
	output wire io_write_last;
	input io_ntwDataUnitOccupancy;
	wire [63:0] currLen;
	wire _taskQueueBuffer_io_enq_ready;
	wire [127:0] _taskQueueBuffer_io_deq_bits;
	wire _taskQueueBuffer_io_count;
	wire _wrRespQueue__io_enq_ready;
	wire _wrRespQueue__io_deq_valid;
	wire _wrReqData__deq_q_io_enq_ready;
	wire _wrReqData__deq_q_io_deq_valid;
	wire [63:0] _wrReqData__deq_q_io_deq_bits_data;
	wire [7:0] _wrReqData__deq_q_io_deq_bits_strb;
	wire _wrReq__deq_q_io_enq_ready;
	wire _wrReq__deq_q_io_deq_valid;
	wire [5:0] _wrReq__deq_q_io_deq_bits_addr;
	wire _rdRespQueue__io_enq_ready;
	wire _rdRespQueue__io_deq_valid;
	wire [63:0] _rdRespQueue__io_deq_bits_data;
	wire [1:0] _rdRespQueue__io_deq_bits_resp;
	wire _rdReq__deq_q_io_enq_ready;
	wire _rdReq__deq_q_io_deq_valid;
	wire [5:0] _rdReq__deq_q_io_deq_bits_addr;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	wire rdReq = _rdReq__deq_q_io_deq_valid & _rdRespQueue__io_enq_ready;
	wire wrReq = (_wrReq__deq_q_io_deq_valid & _wrReqData__deq_q_io_deq_valid) & _wrRespQueue__io_enq_ready;
	reg [63:0] rAddr;
	reg [63:0] rPause;
	reg [63:0] procInterrupt;
	reg [63:0] maxLength;
	reg [3:0] stateReg;
	reg [63:0] contentionCounter;
	reg networkCongested;
	reg [63:0] fifoTailReg;
	reg [63:0] fifoHeadReg;
	reg popOrPush;
	reg [4:0] memDataCounter;
	wire _GEN = stateReg == 4'h2;
	wire _GEN_0 = stateReg == 4'h4;
	wire _GEN_1 = stateReg == 4'h3;
	wire _GEN_2 = memDataCounter == 5'h01;
	wire _GEN_3 = _GEN | _GEN_0;
	wire _GEN_4 = stateReg == 4'h6;
	wire _GEN_5 = stateReg == 4'h5;
	wire _GEN_6 = (_GEN_0 | _GEN_1) | _GEN_4;
	wire _GEN_7 = _GEN | _GEN_6;
	wire _GEN_8 = stateReg == 4'h7;
	wire _GEN_9 = (_GEN | _GEN_0) | _GEN_1;
	wire _GEN_10 = _GEN_4 | _GEN_5;
	reg [63:0] lengthHistroy;
	wire _GEN_11 = fifoTailReg > fifoHeadReg;
	wire [63:0] _currLen_T = fifoTailReg - fifoHeadReg;
	wire _GEN_12 = fifoTailReg < fifoHeadReg;
	wire [63:0] _currLen_T_4 = (maxLength - fifoHeadReg) + fifoTailReg;
	wire [63:0] _currLen_T_6 = lengthHistroy + 64'h0000000000000001;
	assign currLen = (_GEN_11 ? _currLen_T : (_GEN_12 ? _currLen_T_4 : (popOrPush ? 64'h0000000000000000 : _currLen_T_6)));
	wire [511:0] _GEN_13 = {128'hffffffffffffffffffffffffffffffff, procInterrupt, fifoHeadReg, fifoTailReg, maxLength, rAddr, rPause};
	always @(posedge clock)
		if (reset) begin
			rAddr <= 64'h0000000000000000;
			rPause <= 64'h0000000000000000;
			procInterrupt <= 64'h0000000000000000;
			maxLength <= 64'h0000000000000000;
			stateReg <= 4'h0;
			contentionCounter <= 64'h0000000000000000;
			networkCongested <= 1'h0;
			fifoTailReg <= 64'h0000000000000000;
			fifoHeadReg <= 64'h0000000000000000;
			popOrPush <= 1'h1;
			memDataCounter <= 5'h00;
			lengthHistroy <= 64'h0000000000000000;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_14;
			reg _GEN_15;
			reg _GEN_16;
			reg [63:0] _GEN_17;
			reg _GEN_18;
			reg _GEN_19;
			reg _GEN_20;
			reg [63:0] _GEN_21;
			_GEN_20 = rPause == 64'h0000000000000000;
			_GEN_14 = stateReg == 4'h0;
			_GEN_15 = ((currLen == maxLength) & networkCongested) | (maxLength < (currLen + 64'h0000000000000001));
			_GEN_16 = io_write_data_ready & _GEN_2;
			_GEN_17 = maxLength - 64'h0000000000000001;
			_GEN_18 = _GEN_14 | _GEN_3;
			_GEN_19 = io_read_data_valid & _GEN_2;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h1))
				rAddr <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rAddr[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rAddr[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rAddr[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rAddr[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rAddr[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rAddr[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rAddr[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rAddr[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h0))
				rPause <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rPause[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rPause[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rPause[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rPause[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rPause[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rPause[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rPause[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rPause[7:0])};
			else if (_GEN_14 & (|procInterrupt | _GEN_15))
				rPause <= 64'hffffffffffffffff;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h5))
				procInterrupt <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : procInterrupt[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : procInterrupt[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : procInterrupt[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : procInterrupt[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : procInterrupt[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : procInterrupt[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : procInterrupt[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : procInterrupt[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h2))
				maxLength <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : maxLength[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : maxLength[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : maxLength[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : maxLength[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : maxLength[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : maxLength[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : maxLength[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : maxLength[7:0])};
			_GEN_21 = {stateReg, stateReg, stateReg, stateReg, stateReg, (_GEN_20 ? 4'h0 : 4'ha), (_GEN_20 ? 4'h0 : 4'h9), (io_connNetwork_ctrl_serveStealReq_ready ? 4'h7 : (networkCongested | (|procInterrupt) ? 4'h0 : stateReg)), (io_connNetwork_data_qOutTask_ready | networkCongested ? 4'h0 : 4'h7), (io_read_address_ready ? 4'h5 : stateReg), (_GEN_19 ? 4'h8 : stateReg), (io_write_address_ready ? 4'h3 : stateReg), (_GEN_16 ? 4'h0 : stateReg), (~_taskQueueBuffer_io_count & io_connNetwork_data_availableTask_valid ? 4'h4 : (io_connNetwork_data_availableTask_valid & networkCongested ? 4'h2 : (networkCongested ? stateReg : 4'h0))), stateReg, (|procInterrupt ? 4'ha : (_GEN_15 ? 4'h9 : (networkCongested & _taskQueueBuffer_io_count ? 4'h4 : (networkCongested ? 4'h2 : ((~networkCongested & |currLen) & ~_taskQueueBuffer_io_count ? 4'h6 : (~networkCongested & _taskQueueBuffer_io_count ? 4'h7 : stateReg))))))};
			stateReg <= _GEN_21[stateReg * 4+:4];
			if (io_ntwDataUnitOccupancy & (contentionCounter != 64'h0000000000000020))
				contentionCounter <= contentionCounter + 64'h0000000000000001;
			else if (|contentionCounter & ~io_ntwDataUnitOccupancy)
				contentionCounter <= contentionCounter - 64'h0000000000000001;
			networkCongested <= (contentionCounter > 64'h000000000000001a) | ((contentionCounter > 64'h0000000000000018) & networkCongested);
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h3))
				fifoTailReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoTailReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoTailReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoTailReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoTailReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoTailReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoTailReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoTailReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoTailReg[7:0])};
			else if (_GEN_18 | ~_GEN_1)
				;
			else begin : sv2v_autoblock_2
				reg _GEN_22;
				_GEN_22 = fifoTailReg < _GEN_17;
				if (_GEN_16) begin
					if (_GEN_22)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
				else if (io_write_data_ready) begin
					if (_GEN_22)
						fifoTailReg <= fifoTailReg + 64'h0000000000000001;
					else
						fifoTailReg <= 64'h0000000000000000;
				end
			end
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h4))
				fifoHeadReg <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : fifoHeadReg[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : fifoHeadReg[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : fifoHeadReg[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : fifoHeadReg[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : fifoHeadReg[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : fifoHeadReg[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : fifoHeadReg[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : fifoHeadReg[7:0])};
			else if ((_GEN_14 | _GEN_7) | ~_GEN_5)
				;
			else begin : sv2v_autoblock_3
				reg _GEN_23;
				_GEN_23 = fifoHeadReg < _GEN_17;
				if (_GEN_19) begin
					if (_GEN_23)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
				else if (io_read_data_valid) begin
					if (_GEN_23)
						fifoHeadReg <= fifoHeadReg + 64'h0000000000000001;
					else
						fifoHeadReg <= 64'h0000000000000000;
				end
			end
			if (~_GEN_18) begin
				if (_GEN_1)
					popOrPush <= ~_GEN_16 & popOrPush;
				else
					popOrPush <= ((~_GEN_4 & _GEN_5) & _GEN_19) | popOrPush;
			end
			if (~(_GEN_14 | _GEN)) begin
				if (_GEN_0) begin
					if (io_write_address_ready)
						memDataCounter <= 5'h01;
				end
				else if (_GEN_1) begin
					if (_GEN_16 | ~io_write_data_ready)
						;
					else
						memDataCounter <= memDataCounter - 5'h01;
				end
				else if (_GEN_4) begin
					if (io_read_address_ready)
						memDataCounter <= (currLen == 64'h0000000000000000 ? currLen[4:0] : 5'h01);
				end
				else if ((~_GEN_5 | _GEN_19) | ~io_read_data_valid)
					;
				else
					memDataCounter <= memDataCounter - 5'h01;
			end
			if (_GEN_11 | _GEN_12) begin
				if (_GEN_11)
					lengthHistroy <= _currLen_T;
				else if (_GEN_12)
					lengthHistroy <= _currLen_T_4;
				else if (popOrPush)
					lengthHistroy <= 64'h0000000000000000;
				else
					lengthHistroy <= _currLen_T_6;
			end
		end
	Queue2_AddressChannel_2 s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_ar_ready),
		.io_enq_valid(io_axi_mgmt_ar_valid),
		.io_enq_bits_addr(io_axi_mgmt_ar_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_ar_bits_prot),
		.io_deq_ready(_rdReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_rdRespQueue__io_deq_valid),
		.io_enq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_enq_bits_resp(_rdRespQueue__io_deq_bits_resp),
		.io_deq_ready(io_axi_mgmt_r_ready),
		.io_deq_valid(io_axi_mgmt_r_valid),
		.io_deq_bits_data(io_axi_mgmt_r_bits_data),
		.io_deq_bits_resp(io_axi_mgmt_r_bits_resp)
	);
	Queue2_AddressChannel_2 s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_aw_ready),
		.io_enq_valid(io_axi_mgmt_aw_valid),
		.io_enq_bits_addr(io_axi_mgmt_aw_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_aw_bits_prot),
		.io_deq_ready(_wrReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_w_ready),
		.io_enq_valid(io_axi_mgmt_w_valid),
		.io_enq_bits_data(io_axi_mgmt_w_bits_data),
		.io_enq_bits_strb(io_axi_mgmt_w_bits_strb),
		.io_deq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_wrRespQueue__io_deq_valid),
		.io_enq_bits_resp(2'h0),
		.io_deq_ready(io_axi_mgmt_b_ready),
		.io_deq_valid(io_axi_mgmt_b_valid),
		.io_deq_bits_resp(io_axi_mgmt_b_bits_resp)
	);
	Queue1_AddressChannel rdReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_deq_ready(rdReq),
		.io_deq_valid(_rdReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_rdReq__deq_q_io_deq_bits_addr)
	);
	Queue1_ReadDataChannel rdRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdRespQueue__io_enq_ready),
		.io_enq_valid(rdReq),
		.io_enq_bits_data(_GEN_13[_rdReq__deq_q_io_deq_bits_addr[5:3] * 64+:64]),
		.io_deq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_deq_valid(_rdRespQueue__io_deq_valid),
		.io_deq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_deq_bits_resp(_rdRespQueue__io_deq_bits_resp)
	);
	Queue1_AddressChannel wrReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_wrReq__deq_q_io_deq_bits_addr)
	);
	Queue1_WriteDataChannel wrReqData__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_enq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_enq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReqData__deq_q_io_deq_valid),
		.io_deq_bits_data(_wrReqData__deq_q_io_deq_bits_data),
		.io_deq_bits_strb(_wrReqData__deq_q_io_deq_bits_strb)
	);
	Queue1_WriteResponseChannel wrRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrRespQueue__io_enq_ready),
		.io_enq_valid(wrReq),
		.io_deq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_deq_valid(_wrRespQueue__io_deq_valid)
	);
	Queue1_UInt_1 taskQueueBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_taskQueueBuffer_io_enq_ready),
		.io_enq_valid((_GEN ? io_connNetwork_data_availableTask_valid : (~_GEN_6 & _GEN_5) & io_read_data_valid)),
		.io_enq_bits((_GEN ? io_connNetwork_data_availableTask_bits : (_GEN_6 | ~_GEN_5 ? 128'h00000000000000000000000000000000 : io_read_data_bits))),
		.io_deq_ready(~_GEN_3 & (_GEN_1 ? io_write_data_ready : (~_GEN_10 & _GEN_8) & io_connNetwork_data_qOutTask_ready)),
		.io_deq_bits(_taskQueueBuffer_io_deq_bits),
		.io_count(_taskQueueBuffer_io_count)
	);
	assign io_connNetwork_ctrl_serveStealReq_valid = ~(((((_GEN | _GEN_0) | _GEN_1) | _GEN_4) | _GEN_5) | _GEN_8) & (stateReg == 4'h8);
	assign io_connNetwork_data_availableTask_ready = _GEN & _taskQueueBuffer_io_enq_ready;
	assign io_connNetwork_data_qOutTask_valid = ~(((_GEN | _GEN_0) | _GEN_1) | _GEN_10) & _GEN_8;
	assign io_connNetwork_data_qOutTask_bits = _taskQueueBuffer_io_deq_bits;
	assign io_read_address_valid = ~_GEN_9 & _GEN_4;
	assign io_read_address_bits = (_GEN_9 | ~_GEN_4 ? 64'h0000000000000000 : {fifoHeadReg[59:0], 4'h0} + rAddr);
	assign io_read_data_ready = ~_GEN_7 & _GEN_5;
	assign io_read_burst_len = (_GEN_9 | ~(_GEN_4 & (currLen == 64'h0000000000000000)) ? 4'h0 : currLen[3:0] - 4'h1);
	assign io_write_address_valid = ~_GEN & _GEN_0;
	assign io_write_address_bits = (_GEN | ~_GEN_0 ? 64'h0000000000000000 : {fifoTailReg[59:0], 4'h0} + rAddr);
	assign io_write_data_valid = ~_GEN_3 & _GEN_1;
	assign io_write_data_bits = _taskQueueBuffer_io_deq_bits;
	assign io_write_last = (~_GEN_3 & _GEN_1) & _GEN_2;
endmodule
module RVtoAXIBridge_1 (
	clock,
	reset,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_writeBurst_last,
	io_readBurst_len,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_ar_bits_len,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data,
	axi_aw_ready,
	axi_aw_valid,
	axi_aw_bits_addr,
	axi_w_ready,
	axi_w_valid,
	axi_w_bits_data,
	axi_w_bits_last,
	axi_b_valid
);
	input clock;
	input reset;
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [127:0] io_read_data_bits;
	output wire io_write_address_ready;
	input io_write_address_valid;
	input [63:0] io_write_address_bits;
	output wire io_write_data_ready;
	input io_write_data_valid;
	input [127:0] io_write_data_bits;
	input io_writeBurst_last;
	input [3:0] io_readBurst_len;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire [7:0] axi_ar_bits_len;
	output wire axi_r_ready;
	input axi_r_valid;
	input [127:0] axi_r_bits_data;
	input axi_aw_ready;
	output wire axi_aw_valid;
	output wire [63:0] axi_aw_bits_addr;
	input axi_w_ready;
	output wire axi_w_valid;
	output wire [127:0] axi_w_bits_data;
	output wire axi_w_bits_last;
	input axi_b_valid;
	reg writeHandshakeDetector;
	wire axi_w_valid_0 = (io_write_data_valid & axi_w_ready) & ~writeHandshakeDetector;
	always @(posedge clock)
		if (reset)
			writeHandshakeDetector <= 1'h0;
		else if (axi_w_valid_0)
			writeHandshakeDetector <= io_writeBurst_last | writeHandshakeDetector;
		else
			writeHandshakeDetector <= ~axi_b_valid & writeHandshakeDetector;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign io_write_address_ready = axi_aw_ready;
	assign io_write_data_ready = axi_w_ready & ~writeHandshakeDetector;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_ar_bits_len = {4'h0, io_readBurst_len};
	assign axi_r_ready = io_read_data_ready;
	assign axi_aw_valid = io_write_address_valid;
	assign axi_aw_bits_addr = io_write_address_bits;
	assign axi_w_valid = axi_w_valid_0;
	assign axi_w_bits_data = io_write_data_bits;
	assign axi_w_bits_last = io_writeBurst_last;
endmodule
module AxiWriteBuffer_1 (
	clock,
	reset,
	s_axi_ar_ready,
	s_axi_ar_valid,
	s_axi_ar_bits_addr,
	s_axi_ar_bits_len,
	s_axi_r_ready,
	s_axi_r_valid,
	s_axi_r_bits_data,
	s_axi_aw_ready,
	s_axi_aw_valid,
	s_axi_aw_bits_addr,
	s_axi_w_ready,
	s_axi_w_valid,
	s_axi_w_bits_data,
	s_axi_w_bits_last,
	s_axi_b_valid,
	m_axi_ar_ready,
	m_axi_ar_valid,
	m_axi_ar_bits_addr,
	m_axi_ar_bits_len,
	m_axi_ar_bits_size,
	m_axi_ar_bits_burst,
	m_axi_ar_bits_lock,
	m_axi_ar_bits_cache,
	m_axi_ar_bits_prot,
	m_axi_ar_bits_qos,
	m_axi_ar_bits_region,
	m_axi_r_ready,
	m_axi_r_valid,
	m_axi_r_bits_data,
	m_axi_aw_ready,
	m_axi_aw_valid,
	m_axi_aw_bits_addr,
	m_axi_aw_bits_len,
	m_axi_aw_bits_size,
	m_axi_aw_bits_burst,
	m_axi_aw_bits_lock,
	m_axi_aw_bits_cache,
	m_axi_aw_bits_prot,
	m_axi_aw_bits_qos,
	m_axi_aw_bits_region,
	m_axi_w_ready,
	m_axi_w_valid,
	m_axi_w_bits_data,
	m_axi_w_bits_last,
	m_axi_b_valid
);
	input clock;
	input reset;
	output wire s_axi_ar_ready;
	input s_axi_ar_valid;
	input [63:0] s_axi_ar_bits_addr;
	input [7:0] s_axi_ar_bits_len;
	input s_axi_r_ready;
	output wire s_axi_r_valid;
	output wire [127:0] s_axi_r_bits_data;
	output wire s_axi_aw_ready;
	input s_axi_aw_valid;
	input [63:0] s_axi_aw_bits_addr;
	output wire s_axi_w_ready;
	input s_axi_w_valid;
	input [127:0] s_axi_w_bits_data;
	input s_axi_w_bits_last;
	output wire s_axi_b_valid;
	input m_axi_ar_ready;
	output wire m_axi_ar_valid;
	output wire [63:0] m_axi_ar_bits_addr;
	output wire [7:0] m_axi_ar_bits_len;
	output wire [2:0] m_axi_ar_bits_size;
	output wire [1:0] m_axi_ar_bits_burst;
	output wire m_axi_ar_bits_lock;
	output wire [3:0] m_axi_ar_bits_cache;
	output wire [2:0] m_axi_ar_bits_prot;
	output wire [3:0] m_axi_ar_bits_qos;
	output wire [3:0] m_axi_ar_bits_region;
	output wire m_axi_r_ready;
	input m_axi_r_valid;
	input [127:0] m_axi_r_bits_data;
	input m_axi_aw_ready;
	output wire m_axi_aw_valid;
	output wire [63:0] m_axi_aw_bits_addr;
	output wire [7:0] m_axi_aw_bits_len;
	output wire [2:0] m_axi_aw_bits_size;
	output wire [1:0] m_axi_aw_bits_burst;
	output wire m_axi_aw_bits_lock;
	output wire [3:0] m_axi_aw_bits_cache;
	output wire [2:0] m_axi_aw_bits_prot;
	output wire [3:0] m_axi_aw_bits_qos;
	output wire [3:0] m_axi_aw_bits_region;
	input m_axi_w_ready;
	output wire m_axi_w_valid;
	output wire [127:0] m_axi_w_bits_data;
	output wire m_axi_w_bits_last;
	input m_axi_b_valid;
	wire s_axi_aw_ready_0;
	wire _sinkBuffered__sinkBuffer_1_io_enq_ready;
	wire _sinkBuffered__sinkBuffer_io_enq_ready;
	wire _counter_io_empty;
	wire _counter_io_full;
	wire _counter_io_incEn_T = s_axi_aw_ready_0 & s_axi_aw_valid;
	assign s_axi_aw_ready_0 = (_sinkBuffered__sinkBuffer_io_enq_ready & s_axi_aw_valid) & ~_counter_io_full;
	wire s_axi_ar_ready_0 = ((_sinkBuffered__sinkBuffer_1_io_enq_ready & s_axi_ar_valid) & _counter_io_empty) & ~_counter_io_incEn_T;
	Counter counter(
		.clock(clock),
		.reset(reset),
		.io_incEn(_counter_io_incEn_T),
		.io_decEn(m_axi_b_valid),
		.io_empty(_counter_io_empty),
		.io_full(_counter_io_full)
	);
	Queue2_WriteAddressChannel sinkBuffered__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_io_enq_ready),
		.io_enq_valid(s_axi_aw_ready_0),
		.io_enq_bits_addr(s_axi_aw_bits_addr),
		.io_enq_bits_size(3'h4),
		.io_deq_ready(m_axi_aw_ready),
		.io_deq_valid(m_axi_aw_valid),
		.io_deq_bits_addr(m_axi_aw_bits_addr),
		.io_deq_bits_len(m_axi_aw_bits_len),
		.io_deq_bits_size(m_axi_aw_bits_size),
		.io_deq_bits_burst(m_axi_aw_bits_burst),
		.io_deq_bits_lock(m_axi_aw_bits_lock),
		.io_deq_bits_cache(m_axi_aw_bits_cache),
		.io_deq_bits_prot(m_axi_aw_bits_prot),
		.io_deq_bits_qos(m_axi_aw_bits_qos),
		.io_deq_bits_region(m_axi_aw_bits_region)
	);
	Queue2_ReadAddressChannel sinkBuffered__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_sinkBuffered__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(s_axi_ar_ready_0),
		.io_enq_bits_addr(s_axi_ar_bits_addr),
		.io_enq_bits_len(s_axi_ar_bits_len),
		.io_enq_bits_size(3'h4),
		.io_deq_ready(m_axi_ar_ready),
		.io_deq_valid(m_axi_ar_valid),
		.io_deq_bits_addr(m_axi_ar_bits_addr),
		.io_deq_bits_len(m_axi_ar_bits_len),
		.io_deq_bits_size(m_axi_ar_bits_size),
		.io_deq_bits_burst(m_axi_ar_bits_burst),
		.io_deq_bits_lock(m_axi_ar_bits_lock),
		.io_deq_bits_cache(m_axi_ar_bits_cache),
		.io_deq_bits_prot(m_axi_ar_bits_prot),
		.io_deq_bits_qos(m_axi_ar_bits_qos),
		.io_deq_bits_region(m_axi_ar_bits_region)
	);
	assign s_axi_ar_ready = s_axi_ar_ready_0;
	assign s_axi_r_valid = m_axi_r_valid;
	assign s_axi_r_bits_data = m_axi_r_bits_data;
	assign s_axi_aw_ready = s_axi_aw_ready_0;
	assign s_axi_w_ready = m_axi_w_ready;
	assign s_axi_b_valid = m_axi_b_valid;
	assign m_axi_r_ready = s_axi_r_ready;
	assign m_axi_w_valid = s_axi_w_valid;
	assign m_axi_w_bits_data = s_axi_w_bits_data;
	assign m_axi_w_bits_last = s_axi_w_bits_last;
endmodule
module AxisDownscaler_64 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataOut_TREADY,
	io_dataOut_TVALID
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	reg writeCounter;
	always @(posedge clock)
		if (reset)
			writeCounter <= 1'h0;
		else
			writeCounter <= ~io_dataIn_TVALID & writeCounter;
	assign io_dataIn_TREADY = 1'h1;
	assign io_dataOut_TVALID = 1'h0;
endmodule
module AxisDataWidthConverter_128 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataOut_TREADY,
	io_dataOut_TVALID
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	AxisDownscaler_64 downScaler(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_dataIn_TREADY),
		.io_dataIn_TVALID(io_dataIn_TVALID),
		.io_dataOut_TREADY(io_dataOut_TREADY),
		.io_dataOut_TVALID(io_dataOut_TVALID)
	);
endmodule
module Scheduler_1 (
	clock,
	reset,
	io_export_taskOut_0_TREADY,
	io_export_taskOut_0_TVALID,
	io_export_taskOut_1_TREADY,
	io_export_taskOut_1_TVALID,
	io_export_taskOut_2_TREADY,
	io_export_taskOut_2_TVALID,
	io_export_taskOut_3_TREADY,
	io_export_taskOut_3_TVALID,
	io_export_taskOut_4_TREADY,
	io_export_taskOut_4_TVALID,
	io_export_taskOut_5_TREADY,
	io_export_taskOut_5_TVALID,
	io_export_taskOut_6_TREADY,
	io_export_taskOut_6_TVALID,
	io_export_taskOut_7_TREADY,
	io_export_taskOut_7_TVALID,
	io_export_taskOut_8_TREADY,
	io_export_taskOut_8_TVALID,
	io_export_taskOut_9_TREADY,
	io_export_taskOut_9_TVALID,
	io_export_taskOut_10_TREADY,
	io_export_taskOut_10_TVALID,
	io_export_taskOut_11_TREADY,
	io_export_taskOut_11_TVALID,
	io_export_taskOut_12_TREADY,
	io_export_taskOut_12_TVALID,
	io_export_taskOut_13_TREADY,
	io_export_taskOut_13_TVALID,
	io_export_taskOut_14_TREADY,
	io_export_taskOut_14_TVALID,
	io_export_taskOut_15_TREADY,
	io_export_taskOut_15_TVALID,
	io_internal_vss_axi_full_0_ar_ready,
	io_internal_vss_axi_full_0_ar_valid,
	io_internal_vss_axi_full_0_ar_bits_addr,
	io_internal_vss_axi_full_0_ar_bits_len,
	io_internal_vss_axi_full_0_ar_bits_size,
	io_internal_vss_axi_full_0_ar_bits_burst,
	io_internal_vss_axi_full_0_ar_bits_lock,
	io_internal_vss_axi_full_0_ar_bits_cache,
	io_internal_vss_axi_full_0_ar_bits_prot,
	io_internal_vss_axi_full_0_ar_bits_qos,
	io_internal_vss_axi_full_0_ar_bits_region,
	io_internal_vss_axi_full_0_r_ready,
	io_internal_vss_axi_full_0_r_valid,
	io_internal_vss_axi_full_0_r_bits_data,
	io_internal_vss_axi_full_0_aw_ready,
	io_internal_vss_axi_full_0_aw_valid,
	io_internal_vss_axi_full_0_aw_bits_addr,
	io_internal_vss_axi_full_0_aw_bits_len,
	io_internal_vss_axi_full_0_aw_bits_size,
	io_internal_vss_axi_full_0_aw_bits_burst,
	io_internal_vss_axi_full_0_aw_bits_lock,
	io_internal_vss_axi_full_0_aw_bits_cache,
	io_internal_vss_axi_full_0_aw_bits_prot,
	io_internal_vss_axi_full_0_aw_bits_qos,
	io_internal_vss_axi_full_0_aw_bits_region,
	io_internal_vss_axi_full_0_w_ready,
	io_internal_vss_axi_full_0_w_valid,
	io_internal_vss_axi_full_0_w_bits_data,
	io_internal_vss_axi_full_0_w_bits_last,
	io_internal_vss_axi_full_0_b_valid,
	io_internal_axi_mgmt_vss_0_ar_ready,
	io_internal_axi_mgmt_vss_0_ar_valid,
	io_internal_axi_mgmt_vss_0_ar_bits_addr,
	io_internal_axi_mgmt_vss_0_ar_bits_prot,
	io_internal_axi_mgmt_vss_0_r_ready,
	io_internal_axi_mgmt_vss_0_r_valid,
	io_internal_axi_mgmt_vss_0_r_bits_data,
	io_internal_axi_mgmt_vss_0_r_bits_resp,
	io_internal_axi_mgmt_vss_0_aw_ready,
	io_internal_axi_mgmt_vss_0_aw_valid,
	io_internal_axi_mgmt_vss_0_aw_bits_addr,
	io_internal_axi_mgmt_vss_0_aw_bits_prot,
	io_internal_axi_mgmt_vss_0_w_ready,
	io_internal_axi_mgmt_vss_0_w_valid,
	io_internal_axi_mgmt_vss_0_w_bits_data,
	io_internal_axi_mgmt_vss_0_w_bits_strb,
	io_internal_axi_mgmt_vss_0_b_ready,
	io_internal_axi_mgmt_vss_0_b_valid,
	io_internal_axi_mgmt_vss_0_b_bits_resp,
	connArgumentNotifier_0_ctrl_serveStealReq_valid,
	connArgumentNotifier_0_ctrl_serveStealReq_ready,
	connArgumentNotifier_0_data_qOutTask_ready,
	connArgumentNotifier_0_data_qOutTask_valid,
	connArgumentNotifier_0_data_qOutTask_bits,
	connArgumentNotifier_1_ctrl_serveStealReq_valid,
	connArgumentNotifier_1_ctrl_serveStealReq_ready,
	connArgumentNotifier_1_data_qOutTask_ready,
	connArgumentNotifier_1_data_qOutTask_valid,
	connArgumentNotifier_1_data_qOutTask_bits,
	connArgumentNotifier_2_ctrl_serveStealReq_valid,
	connArgumentNotifier_2_ctrl_serveStealReq_ready,
	connArgumentNotifier_2_data_qOutTask_ready,
	connArgumentNotifier_2_data_qOutTask_valid,
	connArgumentNotifier_2_data_qOutTask_bits,
	connArgumentNotifier_3_ctrl_serveStealReq_valid,
	connArgumentNotifier_3_ctrl_serveStealReq_ready,
	connArgumentNotifier_3_data_qOutTask_ready,
	connArgumentNotifier_3_data_qOutTask_valid,
	connArgumentNotifier_3_data_qOutTask_bits,
	connArgumentNotifier_4_ctrl_serveStealReq_valid,
	connArgumentNotifier_4_ctrl_serveStealReq_ready,
	connArgumentNotifier_4_data_qOutTask_ready,
	connArgumentNotifier_4_data_qOutTask_valid,
	connArgumentNotifier_4_data_qOutTask_bits,
	connArgumentNotifier_5_ctrl_serveStealReq_valid,
	connArgumentNotifier_5_ctrl_serveStealReq_ready,
	connArgumentNotifier_5_data_qOutTask_ready,
	connArgumentNotifier_5_data_qOutTask_valid,
	connArgumentNotifier_5_data_qOutTask_bits,
	connArgumentNotifier_6_ctrl_serveStealReq_valid,
	connArgumentNotifier_6_ctrl_serveStealReq_ready,
	connArgumentNotifier_6_data_qOutTask_ready,
	connArgumentNotifier_6_data_qOutTask_valid,
	connArgumentNotifier_6_data_qOutTask_bits,
	connArgumentNotifier_7_ctrl_serveStealReq_valid,
	connArgumentNotifier_7_ctrl_serveStealReq_ready,
	connArgumentNotifier_7_data_qOutTask_ready,
	connArgumentNotifier_7_data_qOutTask_valid,
	connArgumentNotifier_7_data_qOutTask_bits,
	connArgumentNotifier_8_ctrl_serveStealReq_valid,
	connArgumentNotifier_8_ctrl_serveStealReq_ready,
	connArgumentNotifier_8_data_qOutTask_ready,
	connArgumentNotifier_8_data_qOutTask_valid,
	connArgumentNotifier_8_data_qOutTask_bits,
	connArgumentNotifier_9_ctrl_serveStealReq_valid,
	connArgumentNotifier_9_ctrl_serveStealReq_ready,
	connArgumentNotifier_9_data_qOutTask_ready,
	connArgumentNotifier_9_data_qOutTask_valid,
	connArgumentNotifier_9_data_qOutTask_bits,
	connArgumentNotifier_10_ctrl_serveStealReq_valid,
	connArgumentNotifier_10_ctrl_serveStealReq_ready,
	connArgumentNotifier_10_data_qOutTask_ready,
	connArgumentNotifier_10_data_qOutTask_valid,
	connArgumentNotifier_10_data_qOutTask_bits,
	connArgumentNotifier_11_ctrl_serveStealReq_valid,
	connArgumentNotifier_11_ctrl_serveStealReq_ready,
	connArgumentNotifier_11_data_qOutTask_ready,
	connArgumentNotifier_11_data_qOutTask_valid,
	connArgumentNotifier_11_data_qOutTask_bits,
	connArgumentNotifier_12_ctrl_serveStealReq_valid,
	connArgumentNotifier_12_ctrl_serveStealReq_ready,
	connArgumentNotifier_12_data_qOutTask_ready,
	connArgumentNotifier_12_data_qOutTask_valid,
	connArgumentNotifier_12_data_qOutTask_bits,
	connArgumentNotifier_13_ctrl_serveStealReq_valid,
	connArgumentNotifier_13_ctrl_serveStealReq_ready,
	connArgumentNotifier_13_data_qOutTask_ready,
	connArgumentNotifier_13_data_qOutTask_valid,
	connArgumentNotifier_13_data_qOutTask_bits,
	connArgumentNotifier_14_ctrl_serveStealReq_valid,
	connArgumentNotifier_14_ctrl_serveStealReq_ready,
	connArgumentNotifier_14_data_qOutTask_ready,
	connArgumentNotifier_14_data_qOutTask_valid,
	connArgumentNotifier_14_data_qOutTask_bits,
	connArgumentNotifier_15_ctrl_serveStealReq_valid,
	connArgumentNotifier_15_ctrl_serveStealReq_ready,
	connArgumentNotifier_15_data_qOutTask_ready,
	connArgumentNotifier_15_data_qOutTask_valid,
	connArgumentNotifier_15_data_qOutTask_bits
);
	input clock;
	input reset;
	input io_export_taskOut_0_TREADY;
	output wire io_export_taskOut_0_TVALID;
	input io_export_taskOut_1_TREADY;
	output wire io_export_taskOut_1_TVALID;
	input io_export_taskOut_2_TREADY;
	output wire io_export_taskOut_2_TVALID;
	input io_export_taskOut_3_TREADY;
	output wire io_export_taskOut_3_TVALID;
	input io_export_taskOut_4_TREADY;
	output wire io_export_taskOut_4_TVALID;
	input io_export_taskOut_5_TREADY;
	output wire io_export_taskOut_5_TVALID;
	input io_export_taskOut_6_TREADY;
	output wire io_export_taskOut_6_TVALID;
	input io_export_taskOut_7_TREADY;
	output wire io_export_taskOut_7_TVALID;
	input io_export_taskOut_8_TREADY;
	output wire io_export_taskOut_8_TVALID;
	input io_export_taskOut_9_TREADY;
	output wire io_export_taskOut_9_TVALID;
	input io_export_taskOut_10_TREADY;
	output wire io_export_taskOut_10_TVALID;
	input io_export_taskOut_11_TREADY;
	output wire io_export_taskOut_11_TVALID;
	input io_export_taskOut_12_TREADY;
	output wire io_export_taskOut_12_TVALID;
	input io_export_taskOut_13_TREADY;
	output wire io_export_taskOut_13_TVALID;
	input io_export_taskOut_14_TREADY;
	output wire io_export_taskOut_14_TVALID;
	input io_export_taskOut_15_TREADY;
	output wire io_export_taskOut_15_TVALID;
	input io_internal_vss_axi_full_0_ar_ready;
	output wire io_internal_vss_axi_full_0_ar_valid;
	output wire [63:0] io_internal_vss_axi_full_0_ar_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_ar_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_ar_bits_burst;
	output wire io_internal_vss_axi_full_0_ar_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_ar_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_ar_bits_region;
	output wire io_internal_vss_axi_full_0_r_ready;
	input io_internal_vss_axi_full_0_r_valid;
	input [127:0] io_internal_vss_axi_full_0_r_bits_data;
	input io_internal_vss_axi_full_0_aw_ready;
	output wire io_internal_vss_axi_full_0_aw_valid;
	output wire [63:0] io_internal_vss_axi_full_0_aw_bits_addr;
	output wire [7:0] io_internal_vss_axi_full_0_aw_bits_len;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_size;
	output wire [1:0] io_internal_vss_axi_full_0_aw_bits_burst;
	output wire io_internal_vss_axi_full_0_aw_bits_lock;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_cache;
	output wire [2:0] io_internal_vss_axi_full_0_aw_bits_prot;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_qos;
	output wire [3:0] io_internal_vss_axi_full_0_aw_bits_region;
	input io_internal_vss_axi_full_0_w_ready;
	output wire io_internal_vss_axi_full_0_w_valid;
	output wire [127:0] io_internal_vss_axi_full_0_w_bits_data;
	output wire io_internal_vss_axi_full_0_w_bits_last;
	input io_internal_vss_axi_full_0_b_valid;
	output wire io_internal_axi_mgmt_vss_0_ar_ready;
	input io_internal_axi_mgmt_vss_0_ar_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_ar_bits_prot;
	input io_internal_axi_mgmt_vss_0_r_ready;
	output wire io_internal_axi_mgmt_vss_0_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vss_0_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vss_0_r_bits_resp;
	output wire io_internal_axi_mgmt_vss_0_aw_ready;
	input io_internal_axi_mgmt_vss_0_aw_valid;
	input [5:0] io_internal_axi_mgmt_vss_0_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vss_0_aw_bits_prot;
	output wire io_internal_axi_mgmt_vss_0_w_ready;
	input io_internal_axi_mgmt_vss_0_w_valid;
	input [63:0] io_internal_axi_mgmt_vss_0_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vss_0_w_bits_strb;
	input io_internal_axi_mgmt_vss_0_b_ready;
	output wire io_internal_axi_mgmt_vss_0_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vss_0_b_bits_resp;
	input connArgumentNotifier_0_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_0_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_0_data_qOutTask_ready;
	input connArgumentNotifier_0_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_0_data_qOutTask_bits;
	input connArgumentNotifier_1_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_1_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_1_data_qOutTask_ready;
	input connArgumentNotifier_1_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_1_data_qOutTask_bits;
	input connArgumentNotifier_2_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_2_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_2_data_qOutTask_ready;
	input connArgumentNotifier_2_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_2_data_qOutTask_bits;
	input connArgumentNotifier_3_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_3_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_3_data_qOutTask_ready;
	input connArgumentNotifier_3_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_3_data_qOutTask_bits;
	input connArgumentNotifier_4_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_4_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_4_data_qOutTask_ready;
	input connArgumentNotifier_4_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_4_data_qOutTask_bits;
	input connArgumentNotifier_5_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_5_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_5_data_qOutTask_ready;
	input connArgumentNotifier_5_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_5_data_qOutTask_bits;
	input connArgumentNotifier_6_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_6_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_6_data_qOutTask_ready;
	input connArgumentNotifier_6_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_6_data_qOutTask_bits;
	input connArgumentNotifier_7_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_7_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_7_data_qOutTask_ready;
	input connArgumentNotifier_7_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_7_data_qOutTask_bits;
	input connArgumentNotifier_8_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_8_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_8_data_qOutTask_ready;
	input connArgumentNotifier_8_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_8_data_qOutTask_bits;
	input connArgumentNotifier_9_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_9_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_9_data_qOutTask_ready;
	input connArgumentNotifier_9_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_9_data_qOutTask_bits;
	input connArgumentNotifier_10_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_10_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_10_data_qOutTask_ready;
	input connArgumentNotifier_10_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_10_data_qOutTask_bits;
	input connArgumentNotifier_11_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_11_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_11_data_qOutTask_ready;
	input connArgumentNotifier_11_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_11_data_qOutTask_bits;
	input connArgumentNotifier_12_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_12_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_12_data_qOutTask_ready;
	input connArgumentNotifier_12_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_12_data_qOutTask_bits;
	input connArgumentNotifier_13_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_13_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_13_data_qOutTask_ready;
	input connArgumentNotifier_13_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_13_data_qOutTask_bits;
	input connArgumentNotifier_14_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_14_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_14_data_qOutTask_ready;
	input connArgumentNotifier_14_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_14_data_qOutTask_bits;
	input connArgumentNotifier_15_ctrl_serveStealReq_valid;
	output wire connArgumentNotifier_15_ctrl_serveStealReq_ready;
	output wire connArgumentNotifier_15_data_qOutTask_ready;
	input connArgumentNotifier_15_data_qOutTask_valid;
	input [127:0] connArgumentNotifier_15_data_qOutTask_bits;
	wire _axis_stream_converters_out_15_io_dataIn_TREADY;
	wire _axis_stream_converters_out_14_io_dataIn_TREADY;
	wire _axis_stream_converters_out_13_io_dataIn_TREADY;
	wire _axis_stream_converters_out_12_io_dataIn_TREADY;
	wire _axis_stream_converters_out_11_io_dataIn_TREADY;
	wire _axis_stream_converters_out_10_io_dataIn_TREADY;
	wire _axis_stream_converters_out_9_io_dataIn_TREADY;
	wire _axis_stream_converters_out_8_io_dataIn_TREADY;
	wire _axis_stream_converters_out_7_io_dataIn_TREADY;
	wire _axis_stream_converters_out_6_io_dataIn_TREADY;
	wire _axis_stream_converters_out_5_io_dataIn_TREADY;
	wire _axis_stream_converters_out_4_io_dataIn_TREADY;
	wire _axis_stream_converters_out_3_io_dataIn_TREADY;
	wire _axis_stream_converters_out_2_io_dataIn_TREADY;
	wire _axis_stream_converters_out_1_io_dataIn_TREADY;
	wire _axis_stream_converters_out_0_io_dataIn_TREADY;
	wire _module_s_axi_ar_ready;
	wire _module_s_axi_r_valid;
	wire [127:0] _module_s_axi_r_bits_data;
	wire _module_s_axi_aw_ready;
	wire _module_s_axi_w_ready;
	wire _module_s_axi_b_valid;
	wire _vssRvm_0_io_read_address_ready;
	wire _vssRvm_0_io_read_data_valid;
	wire [127:0] _vssRvm_0_io_read_data_bits;
	wire _vssRvm_0_io_write_address_ready;
	wire _vssRvm_0_io_write_data_ready;
	wire _vssRvm_0_axi_ar_valid;
	wire [63:0] _vssRvm_0_axi_ar_bits_addr;
	wire [7:0] _vssRvm_0_axi_ar_bits_len;
	wire _vssRvm_0_axi_r_ready;
	wire _vssRvm_0_axi_aw_valid;
	wire [63:0] _vssRvm_0_axi_aw_bits_addr;
	wire _vssRvm_0_axi_w_valid;
	wire [127:0] _vssRvm_0_axi_w_bits_data;
	wire _vssRvm_0_axi_w_bits_last;
	wire _virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid;
	wire _virtualStealServers_0_io_connNetwork_data_availableTask_ready;
	wire _virtualStealServers_0_io_connNetwork_data_qOutTask_valid;
	wire [127:0] _virtualStealServers_0_io_connNetwork_data_qOutTask_bits;
	wire _virtualStealServers_0_io_read_address_valid;
	wire [63:0] _virtualStealServers_0_io_read_address_bits;
	wire _virtualStealServers_0_io_read_data_ready;
	wire [3:0] _virtualStealServers_0_io_read_burst_len;
	wire _virtualStealServers_0_io_write_address_valid;
	wire [63:0] _virtualStealServers_0_io_write_address_bits;
	wire _virtualStealServers_0_io_write_data_valid;
	wire [127:0] _virtualStealServers_0_io_write_data_bits;
	wire _virtualStealServers_0_io_write_last;
	wire _stealNW_TQ_io_connPE_0_pop_valid;
	wire _stealNW_TQ_io_connPE_1_pop_valid;
	wire _stealNW_TQ_io_connPE_2_pop_valid;
	wire _stealNW_TQ_io_connPE_3_pop_valid;
	wire _stealNW_TQ_io_connPE_4_pop_valid;
	wire _stealNW_TQ_io_connPE_5_pop_valid;
	wire _stealNW_TQ_io_connPE_6_pop_valid;
	wire _stealNW_TQ_io_connPE_7_pop_valid;
	wire _stealNW_TQ_io_connPE_8_pop_valid;
	wire _stealNW_TQ_io_connPE_9_pop_valid;
	wire _stealNW_TQ_io_connPE_10_pop_valid;
	wire _stealNW_TQ_io_connPE_11_pop_valid;
	wire _stealNW_TQ_io_connPE_12_pop_valid;
	wire _stealNW_TQ_io_connPE_13_pop_valid;
	wire _stealNW_TQ_io_connPE_14_pop_valid;
	wire _stealNW_TQ_io_connPE_15_pop_valid;
	wire _stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready;
	wire _stealNW_TQ_io_connVSS_0_data_availableTask_valid;
	wire [127:0] _stealNW_TQ_io_connVSS_0_data_availableTask_bits;
	wire _stealNW_TQ_io_connVSS_0_data_qOutTask_ready;
	wire _stealNW_TQ_io_ntwDataUnitOccupancyVSS_0;
	SchedulerLocalNetwork_1 stealNW_TQ(
		.clock(clock),
		.reset(reset),
		.io_connPE_0_pop_ready(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_connPE_0_pop_valid(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_connPE_1_pop_ready(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_connPE_1_pop_valid(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_connPE_2_pop_ready(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_connPE_2_pop_valid(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_connPE_3_pop_ready(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_connPE_3_pop_valid(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_connPE_4_pop_ready(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_connPE_4_pop_valid(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_connPE_5_pop_ready(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_connPE_5_pop_valid(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_connPE_6_pop_ready(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_connPE_6_pop_valid(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_connPE_7_pop_ready(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_connPE_7_pop_valid(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_connPE_8_pop_ready(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_connPE_8_pop_valid(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_connPE_9_pop_ready(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_connPE_9_pop_valid(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_connPE_10_pop_ready(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_connPE_10_pop_valid(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_connPE_11_pop_ready(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_connPE_11_pop_valid(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_connPE_12_pop_ready(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_connPE_12_pop_valid(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_connPE_13_pop_ready(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_connPE_13_pop_valid(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_connPE_14_pop_ready(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_connPE_14_pop_valid(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_connPE_15_pop_ready(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_connPE_15_pop_valid(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_connVSS_0_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connVSS_0_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connVSS_0_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connVSS_0_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connVSS_0_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connVSS_0_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connVSS_0_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connVSS_0_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_connVAS_0_ctrl_serveStealReq_valid(connArgumentNotifier_0_ctrl_serveStealReq_valid),
		.io_connVAS_0_ctrl_serveStealReq_ready(connArgumentNotifier_0_ctrl_serveStealReq_ready),
		.io_connVAS_0_data_qOutTask_ready(connArgumentNotifier_0_data_qOutTask_ready),
		.io_connVAS_0_data_qOutTask_valid(connArgumentNotifier_0_data_qOutTask_valid),
		.io_connVAS_0_data_qOutTask_bits(connArgumentNotifier_0_data_qOutTask_bits),
		.io_connVAS_1_ctrl_serveStealReq_valid(connArgumentNotifier_1_ctrl_serveStealReq_valid),
		.io_connVAS_1_ctrl_serveStealReq_ready(connArgumentNotifier_1_ctrl_serveStealReq_ready),
		.io_connVAS_1_data_qOutTask_ready(connArgumentNotifier_1_data_qOutTask_ready),
		.io_connVAS_1_data_qOutTask_valid(connArgumentNotifier_1_data_qOutTask_valid),
		.io_connVAS_1_data_qOutTask_bits(connArgumentNotifier_1_data_qOutTask_bits),
		.io_connVAS_2_ctrl_serveStealReq_valid(connArgumentNotifier_2_ctrl_serveStealReq_valid),
		.io_connVAS_2_ctrl_serveStealReq_ready(connArgumentNotifier_2_ctrl_serveStealReq_ready),
		.io_connVAS_2_data_qOutTask_ready(connArgumentNotifier_2_data_qOutTask_ready),
		.io_connVAS_2_data_qOutTask_valid(connArgumentNotifier_2_data_qOutTask_valid),
		.io_connVAS_2_data_qOutTask_bits(connArgumentNotifier_2_data_qOutTask_bits),
		.io_connVAS_3_ctrl_serveStealReq_valid(connArgumentNotifier_3_ctrl_serveStealReq_valid),
		.io_connVAS_3_ctrl_serveStealReq_ready(connArgumentNotifier_3_ctrl_serveStealReq_ready),
		.io_connVAS_3_data_qOutTask_ready(connArgumentNotifier_3_data_qOutTask_ready),
		.io_connVAS_3_data_qOutTask_valid(connArgumentNotifier_3_data_qOutTask_valid),
		.io_connVAS_3_data_qOutTask_bits(connArgumentNotifier_3_data_qOutTask_bits),
		.io_connVAS_4_ctrl_serveStealReq_valid(connArgumentNotifier_4_ctrl_serveStealReq_valid),
		.io_connVAS_4_ctrl_serveStealReq_ready(connArgumentNotifier_4_ctrl_serveStealReq_ready),
		.io_connVAS_4_data_qOutTask_ready(connArgumentNotifier_4_data_qOutTask_ready),
		.io_connVAS_4_data_qOutTask_valid(connArgumentNotifier_4_data_qOutTask_valid),
		.io_connVAS_4_data_qOutTask_bits(connArgumentNotifier_4_data_qOutTask_bits),
		.io_connVAS_5_ctrl_serveStealReq_valid(connArgumentNotifier_5_ctrl_serveStealReq_valid),
		.io_connVAS_5_ctrl_serveStealReq_ready(connArgumentNotifier_5_ctrl_serveStealReq_ready),
		.io_connVAS_5_data_qOutTask_ready(connArgumentNotifier_5_data_qOutTask_ready),
		.io_connVAS_5_data_qOutTask_valid(connArgumentNotifier_5_data_qOutTask_valid),
		.io_connVAS_5_data_qOutTask_bits(connArgumentNotifier_5_data_qOutTask_bits),
		.io_connVAS_6_ctrl_serveStealReq_valid(connArgumentNotifier_6_ctrl_serveStealReq_valid),
		.io_connVAS_6_ctrl_serveStealReq_ready(connArgumentNotifier_6_ctrl_serveStealReq_ready),
		.io_connVAS_6_data_qOutTask_ready(connArgumentNotifier_6_data_qOutTask_ready),
		.io_connVAS_6_data_qOutTask_valid(connArgumentNotifier_6_data_qOutTask_valid),
		.io_connVAS_6_data_qOutTask_bits(connArgumentNotifier_6_data_qOutTask_bits),
		.io_connVAS_7_ctrl_serveStealReq_valid(connArgumentNotifier_7_ctrl_serveStealReq_valid),
		.io_connVAS_7_ctrl_serveStealReq_ready(connArgumentNotifier_7_ctrl_serveStealReq_ready),
		.io_connVAS_7_data_qOutTask_ready(connArgumentNotifier_7_data_qOutTask_ready),
		.io_connVAS_7_data_qOutTask_valid(connArgumentNotifier_7_data_qOutTask_valid),
		.io_connVAS_7_data_qOutTask_bits(connArgumentNotifier_7_data_qOutTask_bits),
		.io_connVAS_8_ctrl_serveStealReq_valid(connArgumentNotifier_8_ctrl_serveStealReq_valid),
		.io_connVAS_8_ctrl_serveStealReq_ready(connArgumentNotifier_8_ctrl_serveStealReq_ready),
		.io_connVAS_8_data_qOutTask_ready(connArgumentNotifier_8_data_qOutTask_ready),
		.io_connVAS_8_data_qOutTask_valid(connArgumentNotifier_8_data_qOutTask_valid),
		.io_connVAS_8_data_qOutTask_bits(connArgumentNotifier_8_data_qOutTask_bits),
		.io_connVAS_9_ctrl_serveStealReq_valid(connArgumentNotifier_9_ctrl_serveStealReq_valid),
		.io_connVAS_9_ctrl_serveStealReq_ready(connArgumentNotifier_9_ctrl_serveStealReq_ready),
		.io_connVAS_9_data_qOutTask_ready(connArgumentNotifier_9_data_qOutTask_ready),
		.io_connVAS_9_data_qOutTask_valid(connArgumentNotifier_9_data_qOutTask_valid),
		.io_connVAS_9_data_qOutTask_bits(connArgumentNotifier_9_data_qOutTask_bits),
		.io_connVAS_10_ctrl_serveStealReq_valid(connArgumentNotifier_10_ctrl_serveStealReq_valid),
		.io_connVAS_10_ctrl_serveStealReq_ready(connArgumentNotifier_10_ctrl_serveStealReq_ready),
		.io_connVAS_10_data_qOutTask_ready(connArgumentNotifier_10_data_qOutTask_ready),
		.io_connVAS_10_data_qOutTask_valid(connArgumentNotifier_10_data_qOutTask_valid),
		.io_connVAS_10_data_qOutTask_bits(connArgumentNotifier_10_data_qOutTask_bits),
		.io_connVAS_11_ctrl_serveStealReq_valid(connArgumentNotifier_11_ctrl_serveStealReq_valid),
		.io_connVAS_11_ctrl_serveStealReq_ready(connArgumentNotifier_11_ctrl_serveStealReq_ready),
		.io_connVAS_11_data_qOutTask_ready(connArgumentNotifier_11_data_qOutTask_ready),
		.io_connVAS_11_data_qOutTask_valid(connArgumentNotifier_11_data_qOutTask_valid),
		.io_connVAS_11_data_qOutTask_bits(connArgumentNotifier_11_data_qOutTask_bits),
		.io_connVAS_12_ctrl_serveStealReq_valid(connArgumentNotifier_12_ctrl_serveStealReq_valid),
		.io_connVAS_12_ctrl_serveStealReq_ready(connArgumentNotifier_12_ctrl_serveStealReq_ready),
		.io_connVAS_12_data_qOutTask_ready(connArgumentNotifier_12_data_qOutTask_ready),
		.io_connVAS_12_data_qOutTask_valid(connArgumentNotifier_12_data_qOutTask_valid),
		.io_connVAS_12_data_qOutTask_bits(connArgumentNotifier_12_data_qOutTask_bits),
		.io_connVAS_13_ctrl_serveStealReq_valid(connArgumentNotifier_13_ctrl_serveStealReq_valid),
		.io_connVAS_13_ctrl_serveStealReq_ready(connArgumentNotifier_13_ctrl_serveStealReq_ready),
		.io_connVAS_13_data_qOutTask_ready(connArgumentNotifier_13_data_qOutTask_ready),
		.io_connVAS_13_data_qOutTask_valid(connArgumentNotifier_13_data_qOutTask_valid),
		.io_connVAS_13_data_qOutTask_bits(connArgumentNotifier_13_data_qOutTask_bits),
		.io_connVAS_14_ctrl_serveStealReq_valid(connArgumentNotifier_14_ctrl_serveStealReq_valid),
		.io_connVAS_14_ctrl_serveStealReq_ready(connArgumentNotifier_14_ctrl_serveStealReq_ready),
		.io_connVAS_14_data_qOutTask_ready(connArgumentNotifier_14_data_qOutTask_ready),
		.io_connVAS_14_data_qOutTask_valid(connArgumentNotifier_14_data_qOutTask_valid),
		.io_connVAS_14_data_qOutTask_bits(connArgumentNotifier_14_data_qOutTask_bits),
		.io_connVAS_15_ctrl_serveStealReq_valid(connArgumentNotifier_15_ctrl_serveStealReq_valid),
		.io_connVAS_15_ctrl_serveStealReq_ready(connArgumentNotifier_15_ctrl_serveStealReq_ready),
		.io_connVAS_15_data_qOutTask_ready(connArgumentNotifier_15_data_qOutTask_ready),
		.io_connVAS_15_data_qOutTask_valid(connArgumentNotifier_15_data_qOutTask_valid),
		.io_connVAS_15_data_qOutTask_bits(connArgumentNotifier_15_data_qOutTask_bits),
		.io_ntwDataUnitOccupancyVSS_0(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
	);
	SchedulerServer_1 virtualStealServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ctrl_serveStealReq_valid(_virtualStealServers_0_io_connNetwork_ctrl_serveStealReq_valid),
		.io_connNetwork_ctrl_serveStealReq_ready(_stealNW_TQ_io_connVSS_0_ctrl_serveStealReq_ready),
		.io_connNetwork_data_availableTask_ready(_virtualStealServers_0_io_connNetwork_data_availableTask_ready),
		.io_connNetwork_data_availableTask_valid(_stealNW_TQ_io_connVSS_0_data_availableTask_valid),
		.io_connNetwork_data_availableTask_bits(_stealNW_TQ_io_connVSS_0_data_availableTask_bits),
		.io_connNetwork_data_qOutTask_ready(_stealNW_TQ_io_connVSS_0_data_qOutTask_ready),
		.io_connNetwork_data_qOutTask_valid(_virtualStealServers_0_io_connNetwork_data_qOutTask_valid),
		.io_connNetwork_data_qOutTask_bits(_virtualStealServers_0_io_connNetwork_data_qOutTask_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vss_0_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vss_0_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vss_0_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vss_0_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vss_0_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vss_0_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vss_0_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vss_0_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vss_0_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vss_0_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vss_0_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vss_0_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vss_0_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vss_0_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vss_0_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vss_0_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vss_0_b_bits_resp),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_read_burst_len(_virtualStealServers_0_io_read_burst_len),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_write_last(_virtualStealServers_0_io_write_last),
		.io_ntwDataUnitOccupancy(_stealNW_TQ_io_ntwDataUnitOccupancyVSS_0)
	);
	RVtoAXIBridge_1 vssRvm_0(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_vssRvm_0_io_read_address_ready),
		.io_read_address_valid(_virtualStealServers_0_io_read_address_valid),
		.io_read_address_bits(_virtualStealServers_0_io_read_address_bits),
		.io_read_data_ready(_virtualStealServers_0_io_read_data_ready),
		.io_read_data_valid(_vssRvm_0_io_read_data_valid),
		.io_read_data_bits(_vssRvm_0_io_read_data_bits),
		.io_write_address_ready(_vssRvm_0_io_write_address_ready),
		.io_write_address_valid(_virtualStealServers_0_io_write_address_valid),
		.io_write_address_bits(_virtualStealServers_0_io_write_address_bits),
		.io_write_data_ready(_vssRvm_0_io_write_data_ready),
		.io_write_data_valid(_virtualStealServers_0_io_write_data_valid),
		.io_write_data_bits(_virtualStealServers_0_io_write_data_bits),
		.io_writeBurst_last(_virtualStealServers_0_io_write_last),
		.io_readBurst_len(_virtualStealServers_0_io_read_burst_len),
		.axi_ar_ready(_module_s_axi_ar_ready),
		.axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.axi_r_ready(_vssRvm_0_axi_r_ready),
		.axi_r_valid(_module_s_axi_r_valid),
		.axi_r_bits_data(_module_s_axi_r_bits_data),
		.axi_aw_ready(_module_s_axi_aw_ready),
		.axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.axi_w_ready(_module_s_axi_w_ready),
		.axi_w_valid(_vssRvm_0_axi_w_valid),
		.axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.axi_b_valid(_module_s_axi_b_valid)
	);
	AxiWriteBuffer_1 module_0(
		.clock(clock),
		.reset(reset),
		.s_axi_ar_ready(_module_s_axi_ar_ready),
		.s_axi_ar_valid(_vssRvm_0_axi_ar_valid),
		.s_axi_ar_bits_addr(_vssRvm_0_axi_ar_bits_addr),
		.s_axi_ar_bits_len(_vssRvm_0_axi_ar_bits_len),
		.s_axi_r_ready(_vssRvm_0_axi_r_ready),
		.s_axi_r_valid(_module_s_axi_r_valid),
		.s_axi_r_bits_data(_module_s_axi_r_bits_data),
		.s_axi_aw_ready(_module_s_axi_aw_ready),
		.s_axi_aw_valid(_vssRvm_0_axi_aw_valid),
		.s_axi_aw_bits_addr(_vssRvm_0_axi_aw_bits_addr),
		.s_axi_w_ready(_module_s_axi_w_ready),
		.s_axi_w_valid(_vssRvm_0_axi_w_valid),
		.s_axi_w_bits_data(_vssRvm_0_axi_w_bits_data),
		.s_axi_w_bits_last(_vssRvm_0_axi_w_bits_last),
		.s_axi_b_valid(_module_s_axi_b_valid),
		.m_axi_ar_ready(io_internal_vss_axi_full_0_ar_ready),
		.m_axi_ar_valid(io_internal_vss_axi_full_0_ar_valid),
		.m_axi_ar_bits_addr(io_internal_vss_axi_full_0_ar_bits_addr),
		.m_axi_ar_bits_len(io_internal_vss_axi_full_0_ar_bits_len),
		.m_axi_ar_bits_size(io_internal_vss_axi_full_0_ar_bits_size),
		.m_axi_ar_bits_burst(io_internal_vss_axi_full_0_ar_bits_burst),
		.m_axi_ar_bits_lock(io_internal_vss_axi_full_0_ar_bits_lock),
		.m_axi_ar_bits_cache(io_internal_vss_axi_full_0_ar_bits_cache),
		.m_axi_ar_bits_prot(io_internal_vss_axi_full_0_ar_bits_prot),
		.m_axi_ar_bits_qos(io_internal_vss_axi_full_0_ar_bits_qos),
		.m_axi_ar_bits_region(io_internal_vss_axi_full_0_ar_bits_region),
		.m_axi_r_ready(io_internal_vss_axi_full_0_r_ready),
		.m_axi_r_valid(io_internal_vss_axi_full_0_r_valid),
		.m_axi_r_bits_data(io_internal_vss_axi_full_0_r_bits_data),
		.m_axi_aw_ready(io_internal_vss_axi_full_0_aw_ready),
		.m_axi_aw_valid(io_internal_vss_axi_full_0_aw_valid),
		.m_axi_aw_bits_addr(io_internal_vss_axi_full_0_aw_bits_addr),
		.m_axi_aw_bits_len(io_internal_vss_axi_full_0_aw_bits_len),
		.m_axi_aw_bits_size(io_internal_vss_axi_full_0_aw_bits_size),
		.m_axi_aw_bits_burst(io_internal_vss_axi_full_0_aw_bits_burst),
		.m_axi_aw_bits_lock(io_internal_vss_axi_full_0_aw_bits_lock),
		.m_axi_aw_bits_cache(io_internal_vss_axi_full_0_aw_bits_cache),
		.m_axi_aw_bits_prot(io_internal_vss_axi_full_0_aw_bits_prot),
		.m_axi_aw_bits_qos(io_internal_vss_axi_full_0_aw_bits_qos),
		.m_axi_aw_bits_region(io_internal_vss_axi_full_0_aw_bits_region),
		.m_axi_w_ready(io_internal_vss_axi_full_0_w_ready),
		.m_axi_w_valid(io_internal_vss_axi_full_0_w_valid),
		.m_axi_w_bits_data(io_internal_vss_axi_full_0_w_bits_data),
		.m_axi_w_bits_last(io_internal_vss_axi_full_0_w_bits_last),
		.m_axi_b_valid(io_internal_vss_axi_full_0_b_valid)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_0(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_0_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_0_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_0_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_1(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_1_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_1_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_1_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_2(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_2_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_2_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_2_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_3(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_3_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_3_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_3_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_4(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_4_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_4_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_4_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_5(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_5_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_5_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_5_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_6(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_6_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_6_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_6_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_7(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_7_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_7_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_7_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_8(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_8_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_8_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_8_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_9(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_9_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_9_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_9_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_10(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_10_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_10_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_10_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_11(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_11_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_11_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_11_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_12(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_12_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_12_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_12_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_13(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_13_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_13_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_13_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_14(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_14_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_14_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_14_TVALID)
	);
	AxisDataWidthConverter_128 axis_stream_converters_out_15(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(_stealNW_TQ_io_connPE_15_pop_valid),
		.io_dataOut_TREADY(io_export_taskOut_15_TREADY),
		.io_dataOut_TVALID(io_export_taskOut_15_TVALID)
	);
endmodule
module AllocatorServerNetworkUnit (
	clock,
	reset,
	io_addressIn0_ready,
	io_addressIn0_valid,
	io_addressIn0_bits,
	io_addressIn1_ready,
	io_addressIn1_valid,
	io_addressIn1_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn0_ready;
	input io_addressIn0_valid;
	input [63:0] io_addressIn0_bits;
	output wire io_addressIn1_ready;
	input io_addressIn1_valid;
	input [63:0] io_addressIn1_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	reg priorityReg;
	wire io_addressIn0_ready_0 = stateReg == 2'h0;
	wire _GEN = stateReg == 2'h1;
	wire _GEN_0 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
			priorityReg <= 1'h1;
		end
		else if (io_addressIn0_ready_0) begin
			if (io_addressIn0_valid) begin
				stateReg <= 2'h2;
				addressReg <= io_addressIn0_bits;
				priorityReg <= ~priorityReg;
			end
			else begin
				if (io_addressIn1_valid)
					stateReg <= 2'h1;
				priorityReg <= io_addressIn1_valid ^ priorityReg;
			end
		end
		else begin
			if (_GEN) begin
				if (io_addressIn1_valid) begin
					stateReg <= 2'h2;
					priorityReg <= ~priorityReg;
				end
				else begin
					if (io_addressIn0_valid)
						stateReg <= 2'h0;
					priorityReg <= io_addressIn0_valid ^ priorityReg;
				end
			end
			else if (_GEN_0 & io_addressOut_ready)
				stateReg <= {1'h0, ~priorityReg};
			if (_GEN & io_addressIn1_valid)
				addressReg <= io_addressIn1_bits;
		end
	assign io_addressIn0_ready = io_addressIn0_ready_0;
	assign io_addressIn1_ready = ~io_addressIn0_ready_0 & _GEN;
	assign io_addressOut_valid = ~(io_addressIn0_ready_0 | _GEN) & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module AllocatorNetworkUnit (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits,
	io_casAddressOut_ready,
	io_casAddressOut_valid,
	io_casAddressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	input io_casAddressOut_ready;
	output wire io_casAddressOut_valid;
	output wire [63:0] io_casAddressOut_bits;
	reg stateReg;
	reg [63:0] addressReg;
	reg priorityReg;
	wire _GEN = io_addressOut_ready & io_casAddressOut_ready;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 1'h0;
			addressReg <= 64'h0000000000000000;
			priorityReg <= 1'h1;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_0;
			_GEN_0 = io_addressOut_ready | io_casAddressOut_ready;
			if (stateReg)
				stateReg <= stateReg & ~_GEN_0;
			else
				stateReg <= io_addressIn_valid | stateReg;
			if (~stateReg & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
			priorityReg <= (stateReg & _GEN_0) ^ priorityReg;
		end
	assign io_addressIn_ready = ~stateReg;
	assign io_addressOut_valid = stateReg & (_GEN ? ~priorityReg & io_addressOut_ready : ~io_casAddressOut_ready & io_addressOut_ready);
	assign io_addressOut_bits = addressReg;
	assign io_casAddressOut_valid = (stateReg & (~_GEN | priorityReg)) & io_casAddressOut_ready;
	assign io_casAddressOut_bits = addressReg;
endmodule
module AllocatorClient (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg stateReg;
	reg [63:0] addressReg;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 1'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (stateReg)
				stateReg <= stateReg & ~io_addressOut_ready;
			else
				stateReg <= io_addressIn_valid | stateReg;
			if (~stateReg & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = ~stateReg;
	assign io_addressOut_valid = stateReg;
	assign io_addressOut_bits = addressReg;
endmodule
module ram_32x64 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [4:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [63:0] R0_data;
	input [4:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [63:0] W0_data;
	reg [63:0] Memory [0:31];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue32_UInt (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits;
	reg [4:0] enq_ptr_value;
	reg [4:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 5'h00;
			deq_ptr_value <= 5'h00;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 5'h01;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 5'h01;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_32x64 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module AllocatorBuffer (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	Queue32_UInt q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_addressIn_ready),
		.io_enq_valid(io_addressIn_valid),
		.io_enq_bits(io_addressIn_bits),
		.io_deq_ready(io_addressOut_ready),
		.io_deq_valid(io_addressOut_valid),
		.io_deq_bits(io_addressOut_bits)
	);
endmodule
module AllocatorNetwork (
	clock,
	reset,
	io_connVCAS_0_ready,
	io_connVCAS_0_valid,
	io_connVCAS_0_bits,
	io_connVCAS_1_ready,
	io_connVCAS_1_valid,
	io_connVCAS_1_bits,
	io_connVCAS_2_ready,
	io_connVCAS_2_valid,
	io_connVCAS_2_bits,
	io_connVCAS_3_ready,
	io_connVCAS_3_valid,
	io_connVCAS_3_bits,
	io_connPE_0_ready,
	io_connPE_0_valid,
	io_connPE_1_ready,
	io_connPE_1_valid,
	io_connPE_2_ready,
	io_connPE_2_valid,
	io_connPE_3_ready,
	io_connPE_3_valid,
	io_connPE_4_ready,
	io_connPE_4_valid,
	io_connPE_5_ready,
	io_connPE_5_valid,
	io_connPE_6_ready,
	io_connPE_6_valid,
	io_connPE_7_ready,
	io_connPE_7_valid,
	io_connPE_8_ready,
	io_connPE_8_valid,
	io_connPE_9_ready,
	io_connPE_9_valid,
	io_connPE_10_ready,
	io_connPE_10_valid,
	io_connPE_11_ready,
	io_connPE_11_valid,
	io_connPE_12_ready,
	io_connPE_12_valid,
	io_connPE_13_ready,
	io_connPE_13_valid,
	io_connPE_14_ready,
	io_connPE_14_valid,
	io_connPE_15_ready,
	io_connPE_15_valid,
	io_connPE_16_ready,
	io_connPE_16_valid,
	io_connPE_17_ready,
	io_connPE_17_valid,
	io_connPE_18_ready,
	io_connPE_18_valid,
	io_connPE_19_ready,
	io_connPE_19_valid,
	io_connPE_20_ready,
	io_connPE_20_valid,
	io_connPE_21_ready,
	io_connPE_21_valid,
	io_connPE_22_ready,
	io_connPE_22_valid,
	io_connPE_23_ready,
	io_connPE_23_valid,
	io_connPE_24_ready,
	io_connPE_24_valid,
	io_connPE_25_ready,
	io_connPE_25_valid,
	io_connPE_26_ready,
	io_connPE_26_valid,
	io_connPE_27_ready,
	io_connPE_27_valid,
	io_connPE_28_ready,
	io_connPE_28_valid,
	io_connPE_29_ready,
	io_connPE_29_valid,
	io_connPE_30_ready,
	io_connPE_30_valid,
	io_connPE_31_ready,
	io_connPE_31_valid,
	io_connPE_32_ready,
	io_connPE_32_valid,
	io_connPE_33_ready,
	io_connPE_33_valid,
	io_connPE_34_ready,
	io_connPE_34_valid,
	io_connPE_35_ready,
	io_connPE_35_valid,
	io_connPE_36_ready,
	io_connPE_36_valid,
	io_connPE_37_ready,
	io_connPE_37_valid,
	io_connPE_38_ready,
	io_connPE_38_valid,
	io_connPE_39_ready,
	io_connPE_39_valid,
	io_connPE_40_ready,
	io_connPE_40_valid,
	io_connPE_41_ready,
	io_connPE_41_valid,
	io_connPE_42_ready,
	io_connPE_42_valid,
	io_connPE_43_ready,
	io_connPE_43_valid,
	io_connPE_44_ready,
	io_connPE_44_valid,
	io_connPE_45_ready,
	io_connPE_45_valid,
	io_connPE_46_ready,
	io_connPE_46_valid,
	io_connPE_47_ready,
	io_connPE_47_valid,
	io_connPE_48_ready,
	io_connPE_48_valid,
	io_connPE_49_ready,
	io_connPE_49_valid,
	io_connPE_50_ready,
	io_connPE_50_valid,
	io_connPE_51_ready,
	io_connPE_51_valid,
	io_connPE_52_ready,
	io_connPE_52_valid,
	io_connPE_53_ready,
	io_connPE_53_valid,
	io_connPE_54_ready,
	io_connPE_54_valid,
	io_connPE_55_ready,
	io_connPE_55_valid,
	io_connPE_56_ready,
	io_connPE_56_valid,
	io_connPE_57_ready,
	io_connPE_57_valid,
	io_connPE_58_ready,
	io_connPE_58_valid,
	io_connPE_59_ready,
	io_connPE_59_valid,
	io_connPE_60_ready,
	io_connPE_60_valid,
	io_connPE_61_ready,
	io_connPE_61_valid,
	io_connPE_62_ready,
	io_connPE_62_valid,
	io_connPE_63_ready,
	io_connPE_63_valid
);
	input clock;
	input reset;
	output wire io_connVCAS_0_ready;
	input io_connVCAS_0_valid;
	input [63:0] io_connVCAS_0_bits;
	output wire io_connVCAS_1_ready;
	input io_connVCAS_1_valid;
	input [63:0] io_connVCAS_1_bits;
	output wire io_connVCAS_2_ready;
	input io_connVCAS_2_valid;
	input [63:0] io_connVCAS_2_bits;
	output wire io_connVCAS_3_ready;
	input io_connVCAS_3_valid;
	input [63:0] io_connVCAS_3_bits;
	input io_connPE_0_ready;
	output wire io_connPE_0_valid;
	input io_connPE_1_ready;
	output wire io_connPE_1_valid;
	input io_connPE_2_ready;
	output wire io_connPE_2_valid;
	input io_connPE_3_ready;
	output wire io_connPE_3_valid;
	input io_connPE_4_ready;
	output wire io_connPE_4_valid;
	input io_connPE_5_ready;
	output wire io_connPE_5_valid;
	input io_connPE_6_ready;
	output wire io_connPE_6_valid;
	input io_connPE_7_ready;
	output wire io_connPE_7_valid;
	input io_connPE_8_ready;
	output wire io_connPE_8_valid;
	input io_connPE_9_ready;
	output wire io_connPE_9_valid;
	input io_connPE_10_ready;
	output wire io_connPE_10_valid;
	input io_connPE_11_ready;
	output wire io_connPE_11_valid;
	input io_connPE_12_ready;
	output wire io_connPE_12_valid;
	input io_connPE_13_ready;
	output wire io_connPE_13_valid;
	input io_connPE_14_ready;
	output wire io_connPE_14_valid;
	input io_connPE_15_ready;
	output wire io_connPE_15_valid;
	input io_connPE_16_ready;
	output wire io_connPE_16_valid;
	input io_connPE_17_ready;
	output wire io_connPE_17_valid;
	input io_connPE_18_ready;
	output wire io_connPE_18_valid;
	input io_connPE_19_ready;
	output wire io_connPE_19_valid;
	input io_connPE_20_ready;
	output wire io_connPE_20_valid;
	input io_connPE_21_ready;
	output wire io_connPE_21_valid;
	input io_connPE_22_ready;
	output wire io_connPE_22_valid;
	input io_connPE_23_ready;
	output wire io_connPE_23_valid;
	input io_connPE_24_ready;
	output wire io_connPE_24_valid;
	input io_connPE_25_ready;
	output wire io_connPE_25_valid;
	input io_connPE_26_ready;
	output wire io_connPE_26_valid;
	input io_connPE_27_ready;
	output wire io_connPE_27_valid;
	input io_connPE_28_ready;
	output wire io_connPE_28_valid;
	input io_connPE_29_ready;
	output wire io_connPE_29_valid;
	input io_connPE_30_ready;
	output wire io_connPE_30_valid;
	input io_connPE_31_ready;
	output wire io_connPE_31_valid;
	input io_connPE_32_ready;
	output wire io_connPE_32_valid;
	input io_connPE_33_ready;
	output wire io_connPE_33_valid;
	input io_connPE_34_ready;
	output wire io_connPE_34_valid;
	input io_connPE_35_ready;
	output wire io_connPE_35_valid;
	input io_connPE_36_ready;
	output wire io_connPE_36_valid;
	input io_connPE_37_ready;
	output wire io_connPE_37_valid;
	input io_connPE_38_ready;
	output wire io_connPE_38_valid;
	input io_connPE_39_ready;
	output wire io_connPE_39_valid;
	input io_connPE_40_ready;
	output wire io_connPE_40_valid;
	input io_connPE_41_ready;
	output wire io_connPE_41_valid;
	input io_connPE_42_ready;
	output wire io_connPE_42_valid;
	input io_connPE_43_ready;
	output wire io_connPE_43_valid;
	input io_connPE_44_ready;
	output wire io_connPE_44_valid;
	input io_connPE_45_ready;
	output wire io_connPE_45_valid;
	input io_connPE_46_ready;
	output wire io_connPE_46_valid;
	input io_connPE_47_ready;
	output wire io_connPE_47_valid;
	input io_connPE_48_ready;
	output wire io_connPE_48_valid;
	input io_connPE_49_ready;
	output wire io_connPE_49_valid;
	input io_connPE_50_ready;
	output wire io_connPE_50_valid;
	input io_connPE_51_ready;
	output wire io_connPE_51_valid;
	input io_connPE_52_ready;
	output wire io_connPE_52_valid;
	input io_connPE_53_ready;
	output wire io_connPE_53_valid;
	input io_connPE_54_ready;
	output wire io_connPE_54_valid;
	input io_connPE_55_ready;
	output wire io_connPE_55_valid;
	input io_connPE_56_ready;
	output wire io_connPE_56_valid;
	input io_connPE_57_ready;
	output wire io_connPE_57_valid;
	input io_connPE_58_ready;
	output wire io_connPE_58_valid;
	input io_connPE_59_ready;
	output wire io_connPE_59_valid;
	input io_connPE_60_ready;
	output wire io_connPE_60_valid;
	input io_connPE_61_ready;
	output wire io_connPE_61_valid;
	input io_connPE_62_ready;
	output wire io_connPE_62_valid;
	input io_connPE_63_ready;
	output wire io_connPE_63_valid;
	wire _queues_63_io_addressIn_ready;
	wire _queues_62_io_addressIn_ready;
	wire _queues_61_io_addressIn_ready;
	wire _queues_60_io_addressIn_ready;
	wire _queues_59_io_addressIn_ready;
	wire _queues_58_io_addressIn_ready;
	wire _queues_57_io_addressIn_ready;
	wire _queues_56_io_addressIn_ready;
	wire _queues_55_io_addressIn_ready;
	wire _queues_54_io_addressIn_ready;
	wire _queues_53_io_addressIn_ready;
	wire _queues_52_io_addressIn_ready;
	wire _queues_51_io_addressIn_ready;
	wire _queues_50_io_addressIn_ready;
	wire _queues_49_io_addressIn_ready;
	wire _queues_48_io_addressIn_ready;
	wire _queues_47_io_addressIn_ready;
	wire _queues_46_io_addressIn_ready;
	wire _queues_45_io_addressIn_ready;
	wire _queues_44_io_addressIn_ready;
	wire _queues_43_io_addressIn_ready;
	wire _queues_42_io_addressIn_ready;
	wire _queues_41_io_addressIn_ready;
	wire _queues_40_io_addressIn_ready;
	wire _queues_39_io_addressIn_ready;
	wire _queues_38_io_addressIn_ready;
	wire _queues_37_io_addressIn_ready;
	wire _queues_36_io_addressIn_ready;
	wire _queues_35_io_addressIn_ready;
	wire _queues_34_io_addressIn_ready;
	wire _queues_33_io_addressIn_ready;
	wire _queues_32_io_addressIn_ready;
	wire _queues_31_io_addressIn_ready;
	wire _queues_30_io_addressIn_ready;
	wire _queues_29_io_addressIn_ready;
	wire _queues_28_io_addressIn_ready;
	wire _queues_27_io_addressIn_ready;
	wire _queues_26_io_addressIn_ready;
	wire _queues_25_io_addressIn_ready;
	wire _queues_24_io_addressIn_ready;
	wire _queues_23_io_addressIn_ready;
	wire _queues_22_io_addressIn_ready;
	wire _queues_21_io_addressIn_ready;
	wire _queues_20_io_addressIn_ready;
	wire _queues_19_io_addressIn_ready;
	wire _queues_18_io_addressIn_ready;
	wire _queues_17_io_addressIn_ready;
	wire _queues_16_io_addressIn_ready;
	wire _queues_15_io_addressIn_ready;
	wire _queues_14_io_addressIn_ready;
	wire _queues_13_io_addressIn_ready;
	wire _queues_12_io_addressIn_ready;
	wire _queues_11_io_addressIn_ready;
	wire _queues_10_io_addressIn_ready;
	wire _queues_9_io_addressIn_ready;
	wire _queues_8_io_addressIn_ready;
	wire _queues_7_io_addressIn_ready;
	wire _queues_6_io_addressIn_ready;
	wire _queues_5_io_addressIn_ready;
	wire _queues_4_io_addressIn_ready;
	wire _queues_3_io_addressIn_ready;
	wire _queues_2_io_addressIn_ready;
	wire _queues_1_io_addressIn_ready;
	wire _queues_0_io_addressIn_ready;
	wire _casServers_63_io_addressIn_ready;
	wire _casServers_63_io_addressOut_valid;
	wire [63:0] _casServers_63_io_addressOut_bits;
	wire _casServers_62_io_addressIn_ready;
	wire _casServers_62_io_addressOut_valid;
	wire [63:0] _casServers_62_io_addressOut_bits;
	wire _casServers_61_io_addressIn_ready;
	wire _casServers_61_io_addressOut_valid;
	wire [63:0] _casServers_61_io_addressOut_bits;
	wire _casServers_60_io_addressIn_ready;
	wire _casServers_60_io_addressOut_valid;
	wire [63:0] _casServers_60_io_addressOut_bits;
	wire _casServers_59_io_addressIn_ready;
	wire _casServers_59_io_addressOut_valid;
	wire [63:0] _casServers_59_io_addressOut_bits;
	wire _casServers_58_io_addressIn_ready;
	wire _casServers_58_io_addressOut_valid;
	wire [63:0] _casServers_58_io_addressOut_bits;
	wire _casServers_57_io_addressIn_ready;
	wire _casServers_57_io_addressOut_valid;
	wire [63:0] _casServers_57_io_addressOut_bits;
	wire _casServers_56_io_addressIn_ready;
	wire _casServers_56_io_addressOut_valid;
	wire [63:0] _casServers_56_io_addressOut_bits;
	wire _casServers_55_io_addressIn_ready;
	wire _casServers_55_io_addressOut_valid;
	wire [63:0] _casServers_55_io_addressOut_bits;
	wire _casServers_54_io_addressIn_ready;
	wire _casServers_54_io_addressOut_valid;
	wire [63:0] _casServers_54_io_addressOut_bits;
	wire _casServers_53_io_addressIn_ready;
	wire _casServers_53_io_addressOut_valid;
	wire [63:0] _casServers_53_io_addressOut_bits;
	wire _casServers_52_io_addressIn_ready;
	wire _casServers_52_io_addressOut_valid;
	wire [63:0] _casServers_52_io_addressOut_bits;
	wire _casServers_51_io_addressIn_ready;
	wire _casServers_51_io_addressOut_valid;
	wire [63:0] _casServers_51_io_addressOut_bits;
	wire _casServers_50_io_addressIn_ready;
	wire _casServers_50_io_addressOut_valid;
	wire [63:0] _casServers_50_io_addressOut_bits;
	wire _casServers_49_io_addressIn_ready;
	wire _casServers_49_io_addressOut_valid;
	wire [63:0] _casServers_49_io_addressOut_bits;
	wire _casServers_48_io_addressIn_ready;
	wire _casServers_48_io_addressOut_valid;
	wire [63:0] _casServers_48_io_addressOut_bits;
	wire _casServers_47_io_addressIn_ready;
	wire _casServers_47_io_addressOut_valid;
	wire [63:0] _casServers_47_io_addressOut_bits;
	wire _casServers_46_io_addressIn_ready;
	wire _casServers_46_io_addressOut_valid;
	wire [63:0] _casServers_46_io_addressOut_bits;
	wire _casServers_45_io_addressIn_ready;
	wire _casServers_45_io_addressOut_valid;
	wire [63:0] _casServers_45_io_addressOut_bits;
	wire _casServers_44_io_addressIn_ready;
	wire _casServers_44_io_addressOut_valid;
	wire [63:0] _casServers_44_io_addressOut_bits;
	wire _casServers_43_io_addressIn_ready;
	wire _casServers_43_io_addressOut_valid;
	wire [63:0] _casServers_43_io_addressOut_bits;
	wire _casServers_42_io_addressIn_ready;
	wire _casServers_42_io_addressOut_valid;
	wire [63:0] _casServers_42_io_addressOut_bits;
	wire _casServers_41_io_addressIn_ready;
	wire _casServers_41_io_addressOut_valid;
	wire [63:0] _casServers_41_io_addressOut_bits;
	wire _casServers_40_io_addressIn_ready;
	wire _casServers_40_io_addressOut_valid;
	wire [63:0] _casServers_40_io_addressOut_bits;
	wire _casServers_39_io_addressIn_ready;
	wire _casServers_39_io_addressOut_valid;
	wire [63:0] _casServers_39_io_addressOut_bits;
	wire _casServers_38_io_addressIn_ready;
	wire _casServers_38_io_addressOut_valid;
	wire [63:0] _casServers_38_io_addressOut_bits;
	wire _casServers_37_io_addressIn_ready;
	wire _casServers_37_io_addressOut_valid;
	wire [63:0] _casServers_37_io_addressOut_bits;
	wire _casServers_36_io_addressIn_ready;
	wire _casServers_36_io_addressOut_valid;
	wire [63:0] _casServers_36_io_addressOut_bits;
	wire _casServers_35_io_addressIn_ready;
	wire _casServers_35_io_addressOut_valid;
	wire [63:0] _casServers_35_io_addressOut_bits;
	wire _casServers_34_io_addressIn_ready;
	wire _casServers_34_io_addressOut_valid;
	wire [63:0] _casServers_34_io_addressOut_bits;
	wire _casServers_33_io_addressIn_ready;
	wire _casServers_33_io_addressOut_valid;
	wire [63:0] _casServers_33_io_addressOut_bits;
	wire _casServers_32_io_addressIn_ready;
	wire _casServers_32_io_addressOut_valid;
	wire [63:0] _casServers_32_io_addressOut_bits;
	wire _casServers_31_io_addressIn_ready;
	wire _casServers_31_io_addressOut_valid;
	wire [63:0] _casServers_31_io_addressOut_bits;
	wire _casServers_30_io_addressIn_ready;
	wire _casServers_30_io_addressOut_valid;
	wire [63:0] _casServers_30_io_addressOut_bits;
	wire _casServers_29_io_addressIn_ready;
	wire _casServers_29_io_addressOut_valid;
	wire [63:0] _casServers_29_io_addressOut_bits;
	wire _casServers_28_io_addressIn_ready;
	wire _casServers_28_io_addressOut_valid;
	wire [63:0] _casServers_28_io_addressOut_bits;
	wire _casServers_27_io_addressIn_ready;
	wire _casServers_27_io_addressOut_valid;
	wire [63:0] _casServers_27_io_addressOut_bits;
	wire _casServers_26_io_addressIn_ready;
	wire _casServers_26_io_addressOut_valid;
	wire [63:0] _casServers_26_io_addressOut_bits;
	wire _casServers_25_io_addressIn_ready;
	wire _casServers_25_io_addressOut_valid;
	wire [63:0] _casServers_25_io_addressOut_bits;
	wire _casServers_24_io_addressIn_ready;
	wire _casServers_24_io_addressOut_valid;
	wire [63:0] _casServers_24_io_addressOut_bits;
	wire _casServers_23_io_addressIn_ready;
	wire _casServers_23_io_addressOut_valid;
	wire [63:0] _casServers_23_io_addressOut_bits;
	wire _casServers_22_io_addressIn_ready;
	wire _casServers_22_io_addressOut_valid;
	wire [63:0] _casServers_22_io_addressOut_bits;
	wire _casServers_21_io_addressIn_ready;
	wire _casServers_21_io_addressOut_valid;
	wire [63:0] _casServers_21_io_addressOut_bits;
	wire _casServers_20_io_addressIn_ready;
	wire _casServers_20_io_addressOut_valid;
	wire [63:0] _casServers_20_io_addressOut_bits;
	wire _casServers_19_io_addressIn_ready;
	wire _casServers_19_io_addressOut_valid;
	wire [63:0] _casServers_19_io_addressOut_bits;
	wire _casServers_18_io_addressIn_ready;
	wire _casServers_18_io_addressOut_valid;
	wire [63:0] _casServers_18_io_addressOut_bits;
	wire _casServers_17_io_addressIn_ready;
	wire _casServers_17_io_addressOut_valid;
	wire [63:0] _casServers_17_io_addressOut_bits;
	wire _casServers_16_io_addressIn_ready;
	wire _casServers_16_io_addressOut_valid;
	wire [63:0] _casServers_16_io_addressOut_bits;
	wire _casServers_15_io_addressIn_ready;
	wire _casServers_15_io_addressOut_valid;
	wire [63:0] _casServers_15_io_addressOut_bits;
	wire _casServers_14_io_addressIn_ready;
	wire _casServers_14_io_addressOut_valid;
	wire [63:0] _casServers_14_io_addressOut_bits;
	wire _casServers_13_io_addressIn_ready;
	wire _casServers_13_io_addressOut_valid;
	wire [63:0] _casServers_13_io_addressOut_bits;
	wire _casServers_12_io_addressIn_ready;
	wire _casServers_12_io_addressOut_valid;
	wire [63:0] _casServers_12_io_addressOut_bits;
	wire _casServers_11_io_addressIn_ready;
	wire _casServers_11_io_addressOut_valid;
	wire [63:0] _casServers_11_io_addressOut_bits;
	wire _casServers_10_io_addressIn_ready;
	wire _casServers_10_io_addressOut_valid;
	wire [63:0] _casServers_10_io_addressOut_bits;
	wire _casServers_9_io_addressIn_ready;
	wire _casServers_9_io_addressOut_valid;
	wire [63:0] _casServers_9_io_addressOut_bits;
	wire _casServers_8_io_addressIn_ready;
	wire _casServers_8_io_addressOut_valid;
	wire [63:0] _casServers_8_io_addressOut_bits;
	wire _casServers_7_io_addressIn_ready;
	wire _casServers_7_io_addressOut_valid;
	wire [63:0] _casServers_7_io_addressOut_bits;
	wire _casServers_6_io_addressIn_ready;
	wire _casServers_6_io_addressOut_valid;
	wire [63:0] _casServers_6_io_addressOut_bits;
	wire _casServers_5_io_addressIn_ready;
	wire _casServers_5_io_addressOut_valid;
	wire [63:0] _casServers_5_io_addressOut_bits;
	wire _casServers_4_io_addressIn_ready;
	wire _casServers_4_io_addressOut_valid;
	wire [63:0] _casServers_4_io_addressOut_bits;
	wire _casServers_3_io_addressIn_ready;
	wire _casServers_3_io_addressOut_valid;
	wire [63:0] _casServers_3_io_addressOut_bits;
	wire _casServers_2_io_addressIn_ready;
	wire _casServers_2_io_addressOut_valid;
	wire [63:0] _casServers_2_io_addressOut_bits;
	wire _casServers_1_io_addressIn_ready;
	wire _casServers_1_io_addressOut_valid;
	wire [63:0] _casServers_1_io_addressOut_bits;
	wire _casServers_0_io_addressIn_ready;
	wire _casServers_0_io_addressOut_valid;
	wire [63:0] _casServers_0_io_addressOut_bits;
	wire _networkUnits_63_io_addressIn_ready;
	wire _networkUnits_63_io_casAddressOut_valid;
	wire [63:0] _networkUnits_63_io_casAddressOut_bits;
	wire _networkUnits_62_io_addressIn_ready;
	wire _networkUnits_62_io_addressOut_valid;
	wire [63:0] _networkUnits_62_io_addressOut_bits;
	wire _networkUnits_62_io_casAddressOut_valid;
	wire [63:0] _networkUnits_62_io_casAddressOut_bits;
	wire _networkUnits_61_io_addressIn_ready;
	wire _networkUnits_61_io_addressOut_valid;
	wire [63:0] _networkUnits_61_io_addressOut_bits;
	wire _networkUnits_61_io_casAddressOut_valid;
	wire [63:0] _networkUnits_61_io_casAddressOut_bits;
	wire _networkUnits_60_io_addressIn_ready;
	wire _networkUnits_60_io_addressOut_valid;
	wire [63:0] _networkUnits_60_io_addressOut_bits;
	wire _networkUnits_60_io_casAddressOut_valid;
	wire [63:0] _networkUnits_60_io_casAddressOut_bits;
	wire _networkUnits_59_io_addressIn_ready;
	wire _networkUnits_59_io_addressOut_valid;
	wire [63:0] _networkUnits_59_io_addressOut_bits;
	wire _networkUnits_59_io_casAddressOut_valid;
	wire [63:0] _networkUnits_59_io_casAddressOut_bits;
	wire _networkUnits_58_io_addressIn_ready;
	wire _networkUnits_58_io_addressOut_valid;
	wire [63:0] _networkUnits_58_io_addressOut_bits;
	wire _networkUnits_58_io_casAddressOut_valid;
	wire [63:0] _networkUnits_58_io_casAddressOut_bits;
	wire _networkUnits_57_io_addressIn_ready;
	wire _networkUnits_57_io_addressOut_valid;
	wire [63:0] _networkUnits_57_io_addressOut_bits;
	wire _networkUnits_57_io_casAddressOut_valid;
	wire [63:0] _networkUnits_57_io_casAddressOut_bits;
	wire _networkUnits_56_io_addressIn_ready;
	wire _networkUnits_56_io_addressOut_valid;
	wire [63:0] _networkUnits_56_io_addressOut_bits;
	wire _networkUnits_56_io_casAddressOut_valid;
	wire [63:0] _networkUnits_56_io_casAddressOut_bits;
	wire _networkUnits_55_io_addressIn_ready;
	wire _networkUnits_55_io_addressOut_valid;
	wire [63:0] _networkUnits_55_io_addressOut_bits;
	wire _networkUnits_55_io_casAddressOut_valid;
	wire [63:0] _networkUnits_55_io_casAddressOut_bits;
	wire _networkUnits_54_io_addressIn_ready;
	wire _networkUnits_54_io_addressOut_valid;
	wire [63:0] _networkUnits_54_io_addressOut_bits;
	wire _networkUnits_54_io_casAddressOut_valid;
	wire [63:0] _networkUnits_54_io_casAddressOut_bits;
	wire _networkUnits_53_io_addressIn_ready;
	wire _networkUnits_53_io_addressOut_valid;
	wire [63:0] _networkUnits_53_io_addressOut_bits;
	wire _networkUnits_53_io_casAddressOut_valid;
	wire [63:0] _networkUnits_53_io_casAddressOut_bits;
	wire _networkUnits_52_io_addressIn_ready;
	wire _networkUnits_52_io_addressOut_valid;
	wire [63:0] _networkUnits_52_io_addressOut_bits;
	wire _networkUnits_52_io_casAddressOut_valid;
	wire [63:0] _networkUnits_52_io_casAddressOut_bits;
	wire _networkUnits_51_io_addressIn_ready;
	wire _networkUnits_51_io_addressOut_valid;
	wire [63:0] _networkUnits_51_io_addressOut_bits;
	wire _networkUnits_51_io_casAddressOut_valid;
	wire [63:0] _networkUnits_51_io_casAddressOut_bits;
	wire _networkUnits_50_io_addressIn_ready;
	wire _networkUnits_50_io_addressOut_valid;
	wire [63:0] _networkUnits_50_io_addressOut_bits;
	wire _networkUnits_50_io_casAddressOut_valid;
	wire [63:0] _networkUnits_50_io_casAddressOut_bits;
	wire _networkUnits_49_io_addressIn_ready;
	wire _networkUnits_49_io_addressOut_valid;
	wire [63:0] _networkUnits_49_io_addressOut_bits;
	wire _networkUnits_49_io_casAddressOut_valid;
	wire [63:0] _networkUnits_49_io_casAddressOut_bits;
	wire _networkUnits_48_io_addressIn_ready;
	wire _networkUnits_48_io_addressOut_valid;
	wire [63:0] _networkUnits_48_io_addressOut_bits;
	wire _networkUnits_48_io_casAddressOut_valid;
	wire [63:0] _networkUnits_48_io_casAddressOut_bits;
	wire _networkUnits_47_io_addressIn_ready;
	wire _networkUnits_47_io_addressOut_valid;
	wire [63:0] _networkUnits_47_io_addressOut_bits;
	wire _networkUnits_47_io_casAddressOut_valid;
	wire [63:0] _networkUnits_47_io_casAddressOut_bits;
	wire _networkUnits_46_io_addressIn_ready;
	wire _networkUnits_46_io_addressOut_valid;
	wire [63:0] _networkUnits_46_io_addressOut_bits;
	wire _networkUnits_46_io_casAddressOut_valid;
	wire [63:0] _networkUnits_46_io_casAddressOut_bits;
	wire _networkUnits_45_io_addressIn_ready;
	wire _networkUnits_45_io_addressOut_valid;
	wire [63:0] _networkUnits_45_io_addressOut_bits;
	wire _networkUnits_45_io_casAddressOut_valid;
	wire [63:0] _networkUnits_45_io_casAddressOut_bits;
	wire _networkUnits_44_io_addressIn_ready;
	wire _networkUnits_44_io_addressOut_valid;
	wire [63:0] _networkUnits_44_io_addressOut_bits;
	wire _networkUnits_44_io_casAddressOut_valid;
	wire [63:0] _networkUnits_44_io_casAddressOut_bits;
	wire _networkUnits_43_io_addressIn_ready;
	wire _networkUnits_43_io_addressOut_valid;
	wire [63:0] _networkUnits_43_io_addressOut_bits;
	wire _networkUnits_43_io_casAddressOut_valid;
	wire [63:0] _networkUnits_43_io_casAddressOut_bits;
	wire _networkUnits_42_io_addressIn_ready;
	wire _networkUnits_42_io_addressOut_valid;
	wire [63:0] _networkUnits_42_io_addressOut_bits;
	wire _networkUnits_42_io_casAddressOut_valid;
	wire [63:0] _networkUnits_42_io_casAddressOut_bits;
	wire _networkUnits_41_io_addressIn_ready;
	wire _networkUnits_41_io_addressOut_valid;
	wire [63:0] _networkUnits_41_io_addressOut_bits;
	wire _networkUnits_41_io_casAddressOut_valid;
	wire [63:0] _networkUnits_41_io_casAddressOut_bits;
	wire _networkUnits_40_io_addressIn_ready;
	wire _networkUnits_40_io_addressOut_valid;
	wire [63:0] _networkUnits_40_io_addressOut_bits;
	wire _networkUnits_40_io_casAddressOut_valid;
	wire [63:0] _networkUnits_40_io_casAddressOut_bits;
	wire _networkUnits_39_io_addressIn_ready;
	wire _networkUnits_39_io_addressOut_valid;
	wire [63:0] _networkUnits_39_io_addressOut_bits;
	wire _networkUnits_39_io_casAddressOut_valid;
	wire [63:0] _networkUnits_39_io_casAddressOut_bits;
	wire _networkUnits_38_io_addressIn_ready;
	wire _networkUnits_38_io_addressOut_valid;
	wire [63:0] _networkUnits_38_io_addressOut_bits;
	wire _networkUnits_38_io_casAddressOut_valid;
	wire [63:0] _networkUnits_38_io_casAddressOut_bits;
	wire _networkUnits_37_io_addressIn_ready;
	wire _networkUnits_37_io_addressOut_valid;
	wire [63:0] _networkUnits_37_io_addressOut_bits;
	wire _networkUnits_37_io_casAddressOut_valid;
	wire [63:0] _networkUnits_37_io_casAddressOut_bits;
	wire _networkUnits_36_io_addressIn_ready;
	wire _networkUnits_36_io_addressOut_valid;
	wire [63:0] _networkUnits_36_io_addressOut_bits;
	wire _networkUnits_36_io_casAddressOut_valid;
	wire [63:0] _networkUnits_36_io_casAddressOut_bits;
	wire _networkUnits_35_io_addressIn_ready;
	wire _networkUnits_35_io_addressOut_valid;
	wire [63:0] _networkUnits_35_io_addressOut_bits;
	wire _networkUnits_35_io_casAddressOut_valid;
	wire [63:0] _networkUnits_35_io_casAddressOut_bits;
	wire _networkUnits_34_io_addressIn_ready;
	wire _networkUnits_34_io_addressOut_valid;
	wire [63:0] _networkUnits_34_io_addressOut_bits;
	wire _networkUnits_34_io_casAddressOut_valid;
	wire [63:0] _networkUnits_34_io_casAddressOut_bits;
	wire _networkUnits_33_io_addressIn_ready;
	wire _networkUnits_33_io_addressOut_valid;
	wire [63:0] _networkUnits_33_io_addressOut_bits;
	wire _networkUnits_33_io_casAddressOut_valid;
	wire [63:0] _networkUnits_33_io_casAddressOut_bits;
	wire _networkUnits_32_io_addressIn_ready;
	wire _networkUnits_32_io_addressOut_valid;
	wire [63:0] _networkUnits_32_io_addressOut_bits;
	wire _networkUnits_32_io_casAddressOut_valid;
	wire [63:0] _networkUnits_32_io_casAddressOut_bits;
	wire _networkUnits_31_io_addressIn_ready;
	wire _networkUnits_31_io_addressOut_valid;
	wire [63:0] _networkUnits_31_io_addressOut_bits;
	wire _networkUnits_31_io_casAddressOut_valid;
	wire [63:0] _networkUnits_31_io_casAddressOut_bits;
	wire _networkUnits_30_io_addressIn_ready;
	wire _networkUnits_30_io_addressOut_valid;
	wire [63:0] _networkUnits_30_io_addressOut_bits;
	wire _networkUnits_30_io_casAddressOut_valid;
	wire [63:0] _networkUnits_30_io_casAddressOut_bits;
	wire _networkUnits_29_io_addressIn_ready;
	wire _networkUnits_29_io_addressOut_valid;
	wire [63:0] _networkUnits_29_io_addressOut_bits;
	wire _networkUnits_29_io_casAddressOut_valid;
	wire [63:0] _networkUnits_29_io_casAddressOut_bits;
	wire _networkUnits_28_io_addressIn_ready;
	wire _networkUnits_28_io_addressOut_valid;
	wire [63:0] _networkUnits_28_io_addressOut_bits;
	wire _networkUnits_28_io_casAddressOut_valid;
	wire [63:0] _networkUnits_28_io_casAddressOut_bits;
	wire _networkUnits_27_io_addressIn_ready;
	wire _networkUnits_27_io_addressOut_valid;
	wire [63:0] _networkUnits_27_io_addressOut_bits;
	wire _networkUnits_27_io_casAddressOut_valid;
	wire [63:0] _networkUnits_27_io_casAddressOut_bits;
	wire _networkUnits_26_io_addressIn_ready;
	wire _networkUnits_26_io_addressOut_valid;
	wire [63:0] _networkUnits_26_io_addressOut_bits;
	wire _networkUnits_26_io_casAddressOut_valid;
	wire [63:0] _networkUnits_26_io_casAddressOut_bits;
	wire _networkUnits_25_io_addressIn_ready;
	wire _networkUnits_25_io_addressOut_valid;
	wire [63:0] _networkUnits_25_io_addressOut_bits;
	wire _networkUnits_25_io_casAddressOut_valid;
	wire [63:0] _networkUnits_25_io_casAddressOut_bits;
	wire _networkUnits_24_io_addressIn_ready;
	wire _networkUnits_24_io_addressOut_valid;
	wire [63:0] _networkUnits_24_io_addressOut_bits;
	wire _networkUnits_24_io_casAddressOut_valid;
	wire [63:0] _networkUnits_24_io_casAddressOut_bits;
	wire _networkUnits_23_io_addressIn_ready;
	wire _networkUnits_23_io_addressOut_valid;
	wire [63:0] _networkUnits_23_io_addressOut_bits;
	wire _networkUnits_23_io_casAddressOut_valid;
	wire [63:0] _networkUnits_23_io_casAddressOut_bits;
	wire _networkUnits_22_io_addressIn_ready;
	wire _networkUnits_22_io_addressOut_valid;
	wire [63:0] _networkUnits_22_io_addressOut_bits;
	wire _networkUnits_22_io_casAddressOut_valid;
	wire [63:0] _networkUnits_22_io_casAddressOut_bits;
	wire _networkUnits_21_io_addressIn_ready;
	wire _networkUnits_21_io_addressOut_valid;
	wire [63:0] _networkUnits_21_io_addressOut_bits;
	wire _networkUnits_21_io_casAddressOut_valid;
	wire [63:0] _networkUnits_21_io_casAddressOut_bits;
	wire _networkUnits_20_io_addressIn_ready;
	wire _networkUnits_20_io_addressOut_valid;
	wire [63:0] _networkUnits_20_io_addressOut_bits;
	wire _networkUnits_20_io_casAddressOut_valid;
	wire [63:0] _networkUnits_20_io_casAddressOut_bits;
	wire _networkUnits_19_io_addressIn_ready;
	wire _networkUnits_19_io_addressOut_valid;
	wire [63:0] _networkUnits_19_io_addressOut_bits;
	wire _networkUnits_19_io_casAddressOut_valid;
	wire [63:0] _networkUnits_19_io_casAddressOut_bits;
	wire _networkUnits_18_io_addressIn_ready;
	wire _networkUnits_18_io_addressOut_valid;
	wire [63:0] _networkUnits_18_io_addressOut_bits;
	wire _networkUnits_18_io_casAddressOut_valid;
	wire [63:0] _networkUnits_18_io_casAddressOut_bits;
	wire _networkUnits_17_io_addressIn_ready;
	wire _networkUnits_17_io_addressOut_valid;
	wire [63:0] _networkUnits_17_io_addressOut_bits;
	wire _networkUnits_17_io_casAddressOut_valid;
	wire [63:0] _networkUnits_17_io_casAddressOut_bits;
	wire _networkUnits_16_io_addressIn_ready;
	wire _networkUnits_16_io_addressOut_valid;
	wire [63:0] _networkUnits_16_io_addressOut_bits;
	wire _networkUnits_16_io_casAddressOut_valid;
	wire [63:0] _networkUnits_16_io_casAddressOut_bits;
	wire _networkUnits_15_io_addressIn_ready;
	wire _networkUnits_15_io_addressOut_valid;
	wire [63:0] _networkUnits_15_io_addressOut_bits;
	wire _networkUnits_15_io_casAddressOut_valid;
	wire [63:0] _networkUnits_15_io_casAddressOut_bits;
	wire _networkUnits_14_io_addressIn_ready;
	wire _networkUnits_14_io_addressOut_valid;
	wire [63:0] _networkUnits_14_io_addressOut_bits;
	wire _networkUnits_14_io_casAddressOut_valid;
	wire [63:0] _networkUnits_14_io_casAddressOut_bits;
	wire _networkUnits_13_io_addressIn_ready;
	wire _networkUnits_13_io_addressOut_valid;
	wire [63:0] _networkUnits_13_io_addressOut_bits;
	wire _networkUnits_13_io_casAddressOut_valid;
	wire [63:0] _networkUnits_13_io_casAddressOut_bits;
	wire _networkUnits_12_io_addressIn_ready;
	wire _networkUnits_12_io_addressOut_valid;
	wire [63:0] _networkUnits_12_io_addressOut_bits;
	wire _networkUnits_12_io_casAddressOut_valid;
	wire [63:0] _networkUnits_12_io_casAddressOut_bits;
	wire _networkUnits_11_io_addressIn_ready;
	wire _networkUnits_11_io_addressOut_valid;
	wire [63:0] _networkUnits_11_io_addressOut_bits;
	wire _networkUnits_11_io_casAddressOut_valid;
	wire [63:0] _networkUnits_11_io_casAddressOut_bits;
	wire _networkUnits_10_io_addressIn_ready;
	wire _networkUnits_10_io_addressOut_valid;
	wire [63:0] _networkUnits_10_io_addressOut_bits;
	wire _networkUnits_10_io_casAddressOut_valid;
	wire [63:0] _networkUnits_10_io_casAddressOut_bits;
	wire _networkUnits_9_io_addressIn_ready;
	wire _networkUnits_9_io_addressOut_valid;
	wire [63:0] _networkUnits_9_io_addressOut_bits;
	wire _networkUnits_9_io_casAddressOut_valid;
	wire [63:0] _networkUnits_9_io_casAddressOut_bits;
	wire _networkUnits_8_io_addressIn_ready;
	wire _networkUnits_8_io_addressOut_valid;
	wire [63:0] _networkUnits_8_io_addressOut_bits;
	wire _networkUnits_8_io_casAddressOut_valid;
	wire [63:0] _networkUnits_8_io_casAddressOut_bits;
	wire _networkUnits_7_io_addressIn_ready;
	wire _networkUnits_7_io_addressOut_valid;
	wire [63:0] _networkUnits_7_io_addressOut_bits;
	wire _networkUnits_7_io_casAddressOut_valid;
	wire [63:0] _networkUnits_7_io_casAddressOut_bits;
	wire _networkUnits_6_io_addressIn_ready;
	wire _networkUnits_6_io_addressOut_valid;
	wire [63:0] _networkUnits_6_io_addressOut_bits;
	wire _networkUnits_6_io_casAddressOut_valid;
	wire [63:0] _networkUnits_6_io_casAddressOut_bits;
	wire _networkUnits_5_io_addressIn_ready;
	wire _networkUnits_5_io_addressOut_valid;
	wire [63:0] _networkUnits_5_io_addressOut_bits;
	wire _networkUnits_5_io_casAddressOut_valid;
	wire [63:0] _networkUnits_5_io_casAddressOut_bits;
	wire _networkUnits_4_io_addressIn_ready;
	wire _networkUnits_4_io_addressOut_valid;
	wire [63:0] _networkUnits_4_io_addressOut_bits;
	wire _networkUnits_4_io_casAddressOut_valid;
	wire [63:0] _networkUnits_4_io_casAddressOut_bits;
	wire _networkUnits_3_io_addressIn_ready;
	wire _networkUnits_3_io_addressOut_valid;
	wire [63:0] _networkUnits_3_io_addressOut_bits;
	wire _networkUnits_3_io_casAddressOut_valid;
	wire [63:0] _networkUnits_3_io_casAddressOut_bits;
	wire _networkUnits_2_io_addressIn_ready;
	wire _networkUnits_2_io_addressOut_valid;
	wire [63:0] _networkUnits_2_io_addressOut_bits;
	wire _networkUnits_2_io_casAddressOut_valid;
	wire [63:0] _networkUnits_2_io_casAddressOut_bits;
	wire _networkUnits_1_io_addressIn_ready;
	wire _networkUnits_1_io_addressOut_valid;
	wire [63:0] _networkUnits_1_io_addressOut_bits;
	wire _networkUnits_1_io_casAddressOut_valid;
	wire [63:0] _networkUnits_1_io_casAddressOut_bits;
	wire _networkUnits_0_io_addressIn_ready;
	wire _networkUnits_0_io_addressOut_valid;
	wire [63:0] _networkUnits_0_io_addressOut_bits;
	wire _networkUnits_0_io_casAddressOut_valid;
	wire [63:0] _networkUnits_0_io_casAddressOut_bits;
	wire _vcasNetworkUnits_3_io_addressIn0_ready;
	wire _vcasNetworkUnits_3_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_3_io_addressOut_bits;
	wire _vcasNetworkUnits_2_io_addressIn0_ready;
	wire _vcasNetworkUnits_2_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_2_io_addressOut_bits;
	wire _vcasNetworkUnits_1_io_addressIn0_ready;
	wire _vcasNetworkUnits_1_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_1_io_addressOut_bits;
	wire _vcasNetworkUnits_0_io_addressOut_valid;
	wire [63:0] _vcasNetworkUnits_0_io_addressOut_bits;
	AllocatorServerNetworkUnit vcasNetworkUnits_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(),
		.io_addressIn0_valid(1'h0),
		.io_addressIn0_bits(64'h0000000000000000),
		.io_addressIn1_ready(io_connVCAS_0_ready),
		.io_addressIn1_valid(io_connVCAS_0_valid),
		.io_addressIn1_bits(io_connVCAS_0_bits),
		.io_addressOut_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_0_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_0_io_addressOut_bits)
	);
	AllocatorServerNetworkUnit vcasNetworkUnits_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(_vcasNetworkUnits_1_io_addressIn0_ready),
		.io_addressIn0_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressIn0_bits(_networkUnits_15_io_addressOut_bits),
		.io_addressIn1_ready(io_connVCAS_1_ready),
		.io_addressIn1_valid(io_connVCAS_1_valid),
		.io_addressIn1_bits(io_connVCAS_1_bits),
		.io_addressOut_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_1_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_1_io_addressOut_bits)
	);
	AllocatorServerNetworkUnit vcasNetworkUnits_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(_vcasNetworkUnits_2_io_addressIn0_ready),
		.io_addressIn0_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressIn0_bits(_networkUnits_31_io_addressOut_bits),
		.io_addressIn1_ready(io_connVCAS_2_ready),
		.io_addressIn1_valid(io_connVCAS_2_valid),
		.io_addressIn1_bits(io_connVCAS_2_bits),
		.io_addressOut_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_2_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_2_io_addressOut_bits)
	);
	AllocatorServerNetworkUnit vcasNetworkUnits_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn0_ready(_vcasNetworkUnits_3_io_addressIn0_ready),
		.io_addressIn0_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressIn0_bits(_networkUnits_47_io_addressOut_bits),
		.io_addressIn1_ready(io_connVCAS_3_ready),
		.io_addressIn1_valid(io_connVCAS_3_valid),
		.io_addressIn1_bits(io_connVCAS_3_bits),
		.io_addressOut_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressOut_valid(_vcasNetworkUnits_3_io_addressOut_valid),
		.io_addressOut_bits(_vcasNetworkUnits_3_io_addressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_0_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_0_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_0_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_0_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_0_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_0_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_0_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_1_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_1_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_1_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_1_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_1_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_2_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_2_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_2_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_2_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_2_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_3_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_3_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_3_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_3_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_3_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_4_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_4_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_4_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_4_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_4_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_5_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_5_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_5_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_5_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_5_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_6_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_6_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_6_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_6_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_6_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_7_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_7_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_7_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_7_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_7_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_8_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_8_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_8_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_8_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_8_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_9_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_9_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_9_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_9_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_9_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_10_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_10_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_10_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_10_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_10_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_11_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_11_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_11_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_11_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_11_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_12_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_12_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_12_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_12_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_12_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_13_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_13_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_13_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_13_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_13_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_14_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_14_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_14_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_14_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_14_io_addressOut_bits),
		.io_addressOut_ready(_vcasNetworkUnits_1_io_addressIn0_ready),
		.io_addressOut_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_15_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_15_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_15_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_15_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_1_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_1_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_16_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_16_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_16_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_16_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_16_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_17_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_17_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_17_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_17_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_17_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_18_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_18_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_18_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_18_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_18_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_19_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_19_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_19_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_19_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_19_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_20_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_20_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_20_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_20_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_20_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_21_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_21_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_21_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_21_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_21_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_22_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_22_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_22_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_22_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_22_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_23_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_23_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_23_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_23_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_23_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_24_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_24_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_24_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_24_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_24_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_25_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_25_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_25_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_25_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_25_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_26_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_26_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_26_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_26_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_26_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_27_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_27_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_27_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_27_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_27_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_28_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_28_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_28_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_28_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_28_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_29_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_29_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_29_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_29_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_29_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_30_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_30_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_30_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_30_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_30_io_addressOut_bits),
		.io_addressOut_ready(_vcasNetworkUnits_2_io_addressIn0_ready),
		.io_addressOut_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_31_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_31_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_31_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_31_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_2_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_2_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_32_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_32_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_32_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_32_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_32_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_33_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_33_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_33_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_33_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_33_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_34_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_34_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_34_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_34_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_34_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_35_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_35_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_35_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_35_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_35_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_36_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_36_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_36_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_36_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_36_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_37_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_37_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_37_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_37_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_37_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_38_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_38_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_38_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_38_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_38_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_39_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_39_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_39_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_39_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_39_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_40_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_40_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_40_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_40_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_40_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_41_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_41_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_41_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_41_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_41_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_42_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_42_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_42_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_42_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_42_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_43_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_43_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_43_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_43_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_43_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_44_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_44_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_44_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_44_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_44_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_45_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_45_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_45_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_45_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_45_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_46_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_46_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_46_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_46_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_46_io_addressOut_bits),
		.io_addressOut_ready(_vcasNetworkUnits_3_io_addressIn0_ready),
		.io_addressOut_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_47_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_47_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_47_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_47_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressIn_valid(_vcasNetworkUnits_3_io_addressOut_valid),
		.io_addressIn_bits(_vcasNetworkUnits_3_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_48_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_48_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_48_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_48_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_48_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_49_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_49_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_49_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_49_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_49_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_50_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_50_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_50_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_50_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_50_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_51_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_51_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_51_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_51_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_51_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_52_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_52_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_52_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_52_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_52_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_53_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_53_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_53_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_53_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_53_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_54_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_54_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_54_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_54_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_54_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_55_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_55_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_55_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_55_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_55_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_56_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_56_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_56_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_56_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_56_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_57_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_57_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_57_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_57_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_57_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_58_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_58_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_58_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_58_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_58_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_59_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_59_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_59_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_59_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_59_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_60_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_60_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_60_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_60_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_60_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_61_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_61_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_61_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_61_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_61_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_62_io_addressOut_bits),
		.io_casAddressOut_ready(_casServers_62_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_62_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_62_io_casAddressOut_bits)
	);
	AllocatorNetworkUnit networkUnits_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_62_io_addressOut_bits),
		.io_addressOut_ready(1'h0),
		.io_addressOut_valid(),
		.io_addressOut_bits(),
		.io_casAddressOut_ready(_casServers_63_io_addressIn_ready),
		.io_casAddressOut_valid(_networkUnits_63_io_casAddressOut_valid),
		.io_casAddressOut_bits(_networkUnits_63_io_casAddressOut_bits)
	);
	AllocatorClient casServers_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_0_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_0_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_0_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_0_io_addressIn_ready),
		.io_addressOut_valid(_casServers_0_io_addressOut_valid),
		.io_addressOut_bits(_casServers_0_io_addressOut_bits)
	);
	AllocatorClient casServers_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_1_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_1_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_1_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_1_io_addressIn_ready),
		.io_addressOut_valid(_casServers_1_io_addressOut_valid),
		.io_addressOut_bits(_casServers_1_io_addressOut_bits)
	);
	AllocatorClient casServers_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_2_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_2_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_2_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_2_io_addressIn_ready),
		.io_addressOut_valid(_casServers_2_io_addressOut_valid),
		.io_addressOut_bits(_casServers_2_io_addressOut_bits)
	);
	AllocatorClient casServers_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_3_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_3_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_3_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_3_io_addressIn_ready),
		.io_addressOut_valid(_casServers_3_io_addressOut_valid),
		.io_addressOut_bits(_casServers_3_io_addressOut_bits)
	);
	AllocatorClient casServers_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_4_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_4_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_4_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_4_io_addressIn_ready),
		.io_addressOut_valid(_casServers_4_io_addressOut_valid),
		.io_addressOut_bits(_casServers_4_io_addressOut_bits)
	);
	AllocatorClient casServers_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_5_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_5_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_5_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_5_io_addressIn_ready),
		.io_addressOut_valid(_casServers_5_io_addressOut_valid),
		.io_addressOut_bits(_casServers_5_io_addressOut_bits)
	);
	AllocatorClient casServers_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_6_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_6_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_6_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_6_io_addressIn_ready),
		.io_addressOut_valid(_casServers_6_io_addressOut_valid),
		.io_addressOut_bits(_casServers_6_io_addressOut_bits)
	);
	AllocatorClient casServers_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_7_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_7_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_7_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_7_io_addressIn_ready),
		.io_addressOut_valid(_casServers_7_io_addressOut_valid),
		.io_addressOut_bits(_casServers_7_io_addressOut_bits)
	);
	AllocatorClient casServers_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_8_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_8_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_8_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_8_io_addressIn_ready),
		.io_addressOut_valid(_casServers_8_io_addressOut_valid),
		.io_addressOut_bits(_casServers_8_io_addressOut_bits)
	);
	AllocatorClient casServers_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_9_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_9_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_9_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_9_io_addressIn_ready),
		.io_addressOut_valid(_casServers_9_io_addressOut_valid),
		.io_addressOut_bits(_casServers_9_io_addressOut_bits)
	);
	AllocatorClient casServers_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_10_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_10_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_10_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_10_io_addressIn_ready),
		.io_addressOut_valid(_casServers_10_io_addressOut_valid),
		.io_addressOut_bits(_casServers_10_io_addressOut_bits)
	);
	AllocatorClient casServers_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_11_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_11_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_11_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_11_io_addressIn_ready),
		.io_addressOut_valid(_casServers_11_io_addressOut_valid),
		.io_addressOut_bits(_casServers_11_io_addressOut_bits)
	);
	AllocatorClient casServers_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_12_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_12_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_12_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_12_io_addressIn_ready),
		.io_addressOut_valid(_casServers_12_io_addressOut_valid),
		.io_addressOut_bits(_casServers_12_io_addressOut_bits)
	);
	AllocatorClient casServers_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_13_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_13_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_13_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_13_io_addressIn_ready),
		.io_addressOut_valid(_casServers_13_io_addressOut_valid),
		.io_addressOut_bits(_casServers_13_io_addressOut_bits)
	);
	AllocatorClient casServers_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_14_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_14_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_14_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_14_io_addressIn_ready),
		.io_addressOut_valid(_casServers_14_io_addressOut_valid),
		.io_addressOut_bits(_casServers_14_io_addressOut_bits)
	);
	AllocatorClient casServers_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_15_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_15_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_15_io_addressIn_ready),
		.io_addressOut_valid(_casServers_15_io_addressOut_valid),
		.io_addressOut_bits(_casServers_15_io_addressOut_bits)
	);
	AllocatorClient casServers_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_16_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_16_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_16_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_16_io_addressIn_ready),
		.io_addressOut_valid(_casServers_16_io_addressOut_valid),
		.io_addressOut_bits(_casServers_16_io_addressOut_bits)
	);
	AllocatorClient casServers_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_17_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_17_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_17_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_17_io_addressIn_ready),
		.io_addressOut_valid(_casServers_17_io_addressOut_valid),
		.io_addressOut_bits(_casServers_17_io_addressOut_bits)
	);
	AllocatorClient casServers_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_18_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_18_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_18_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_18_io_addressIn_ready),
		.io_addressOut_valid(_casServers_18_io_addressOut_valid),
		.io_addressOut_bits(_casServers_18_io_addressOut_bits)
	);
	AllocatorClient casServers_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_19_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_19_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_19_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_19_io_addressIn_ready),
		.io_addressOut_valid(_casServers_19_io_addressOut_valid),
		.io_addressOut_bits(_casServers_19_io_addressOut_bits)
	);
	AllocatorClient casServers_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_20_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_20_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_20_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_20_io_addressIn_ready),
		.io_addressOut_valid(_casServers_20_io_addressOut_valid),
		.io_addressOut_bits(_casServers_20_io_addressOut_bits)
	);
	AllocatorClient casServers_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_21_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_21_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_21_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_21_io_addressIn_ready),
		.io_addressOut_valid(_casServers_21_io_addressOut_valid),
		.io_addressOut_bits(_casServers_21_io_addressOut_bits)
	);
	AllocatorClient casServers_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_22_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_22_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_22_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_22_io_addressIn_ready),
		.io_addressOut_valid(_casServers_22_io_addressOut_valid),
		.io_addressOut_bits(_casServers_22_io_addressOut_bits)
	);
	AllocatorClient casServers_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_23_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_23_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_23_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_23_io_addressIn_ready),
		.io_addressOut_valid(_casServers_23_io_addressOut_valid),
		.io_addressOut_bits(_casServers_23_io_addressOut_bits)
	);
	AllocatorClient casServers_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_24_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_24_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_24_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_24_io_addressIn_ready),
		.io_addressOut_valid(_casServers_24_io_addressOut_valid),
		.io_addressOut_bits(_casServers_24_io_addressOut_bits)
	);
	AllocatorClient casServers_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_25_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_25_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_25_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_25_io_addressIn_ready),
		.io_addressOut_valid(_casServers_25_io_addressOut_valid),
		.io_addressOut_bits(_casServers_25_io_addressOut_bits)
	);
	AllocatorClient casServers_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_26_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_26_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_26_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_26_io_addressIn_ready),
		.io_addressOut_valid(_casServers_26_io_addressOut_valid),
		.io_addressOut_bits(_casServers_26_io_addressOut_bits)
	);
	AllocatorClient casServers_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_27_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_27_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_27_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_27_io_addressIn_ready),
		.io_addressOut_valid(_casServers_27_io_addressOut_valid),
		.io_addressOut_bits(_casServers_27_io_addressOut_bits)
	);
	AllocatorClient casServers_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_28_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_28_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_28_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_28_io_addressIn_ready),
		.io_addressOut_valid(_casServers_28_io_addressOut_valid),
		.io_addressOut_bits(_casServers_28_io_addressOut_bits)
	);
	AllocatorClient casServers_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_29_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_29_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_29_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_29_io_addressIn_ready),
		.io_addressOut_valid(_casServers_29_io_addressOut_valid),
		.io_addressOut_bits(_casServers_29_io_addressOut_bits)
	);
	AllocatorClient casServers_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_30_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_30_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_30_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_30_io_addressIn_ready),
		.io_addressOut_valid(_casServers_30_io_addressOut_valid),
		.io_addressOut_bits(_casServers_30_io_addressOut_bits)
	);
	AllocatorClient casServers_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_31_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_31_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_31_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_31_io_addressIn_ready),
		.io_addressOut_valid(_casServers_31_io_addressOut_valid),
		.io_addressOut_bits(_casServers_31_io_addressOut_bits)
	);
	AllocatorClient casServers_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_32_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_32_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_32_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_32_io_addressIn_ready),
		.io_addressOut_valid(_casServers_32_io_addressOut_valid),
		.io_addressOut_bits(_casServers_32_io_addressOut_bits)
	);
	AllocatorClient casServers_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_33_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_33_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_33_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_33_io_addressIn_ready),
		.io_addressOut_valid(_casServers_33_io_addressOut_valid),
		.io_addressOut_bits(_casServers_33_io_addressOut_bits)
	);
	AllocatorClient casServers_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_34_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_34_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_34_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_34_io_addressIn_ready),
		.io_addressOut_valid(_casServers_34_io_addressOut_valid),
		.io_addressOut_bits(_casServers_34_io_addressOut_bits)
	);
	AllocatorClient casServers_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_35_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_35_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_35_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_35_io_addressIn_ready),
		.io_addressOut_valid(_casServers_35_io_addressOut_valid),
		.io_addressOut_bits(_casServers_35_io_addressOut_bits)
	);
	AllocatorClient casServers_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_36_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_36_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_36_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_36_io_addressIn_ready),
		.io_addressOut_valid(_casServers_36_io_addressOut_valid),
		.io_addressOut_bits(_casServers_36_io_addressOut_bits)
	);
	AllocatorClient casServers_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_37_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_37_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_37_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_37_io_addressIn_ready),
		.io_addressOut_valid(_casServers_37_io_addressOut_valid),
		.io_addressOut_bits(_casServers_37_io_addressOut_bits)
	);
	AllocatorClient casServers_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_38_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_38_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_38_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_38_io_addressIn_ready),
		.io_addressOut_valid(_casServers_38_io_addressOut_valid),
		.io_addressOut_bits(_casServers_38_io_addressOut_bits)
	);
	AllocatorClient casServers_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_39_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_39_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_39_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_39_io_addressIn_ready),
		.io_addressOut_valid(_casServers_39_io_addressOut_valid),
		.io_addressOut_bits(_casServers_39_io_addressOut_bits)
	);
	AllocatorClient casServers_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_40_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_40_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_40_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_40_io_addressIn_ready),
		.io_addressOut_valid(_casServers_40_io_addressOut_valid),
		.io_addressOut_bits(_casServers_40_io_addressOut_bits)
	);
	AllocatorClient casServers_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_41_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_41_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_41_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_41_io_addressIn_ready),
		.io_addressOut_valid(_casServers_41_io_addressOut_valid),
		.io_addressOut_bits(_casServers_41_io_addressOut_bits)
	);
	AllocatorClient casServers_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_42_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_42_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_42_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_42_io_addressIn_ready),
		.io_addressOut_valid(_casServers_42_io_addressOut_valid),
		.io_addressOut_bits(_casServers_42_io_addressOut_bits)
	);
	AllocatorClient casServers_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_43_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_43_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_43_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_43_io_addressIn_ready),
		.io_addressOut_valid(_casServers_43_io_addressOut_valid),
		.io_addressOut_bits(_casServers_43_io_addressOut_bits)
	);
	AllocatorClient casServers_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_44_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_44_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_44_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_44_io_addressIn_ready),
		.io_addressOut_valid(_casServers_44_io_addressOut_valid),
		.io_addressOut_bits(_casServers_44_io_addressOut_bits)
	);
	AllocatorClient casServers_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_45_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_45_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_45_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_45_io_addressIn_ready),
		.io_addressOut_valid(_casServers_45_io_addressOut_valid),
		.io_addressOut_bits(_casServers_45_io_addressOut_bits)
	);
	AllocatorClient casServers_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_46_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_46_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_46_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_46_io_addressIn_ready),
		.io_addressOut_valid(_casServers_46_io_addressOut_valid),
		.io_addressOut_bits(_casServers_46_io_addressOut_bits)
	);
	AllocatorClient casServers_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_47_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_47_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_47_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_47_io_addressIn_ready),
		.io_addressOut_valid(_casServers_47_io_addressOut_valid),
		.io_addressOut_bits(_casServers_47_io_addressOut_bits)
	);
	AllocatorClient casServers_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_48_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_48_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_48_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_48_io_addressIn_ready),
		.io_addressOut_valid(_casServers_48_io_addressOut_valid),
		.io_addressOut_bits(_casServers_48_io_addressOut_bits)
	);
	AllocatorClient casServers_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_49_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_49_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_49_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_49_io_addressIn_ready),
		.io_addressOut_valid(_casServers_49_io_addressOut_valid),
		.io_addressOut_bits(_casServers_49_io_addressOut_bits)
	);
	AllocatorClient casServers_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_50_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_50_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_50_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_50_io_addressIn_ready),
		.io_addressOut_valid(_casServers_50_io_addressOut_valid),
		.io_addressOut_bits(_casServers_50_io_addressOut_bits)
	);
	AllocatorClient casServers_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_51_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_51_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_51_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_51_io_addressIn_ready),
		.io_addressOut_valid(_casServers_51_io_addressOut_valid),
		.io_addressOut_bits(_casServers_51_io_addressOut_bits)
	);
	AllocatorClient casServers_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_52_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_52_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_52_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_52_io_addressIn_ready),
		.io_addressOut_valid(_casServers_52_io_addressOut_valid),
		.io_addressOut_bits(_casServers_52_io_addressOut_bits)
	);
	AllocatorClient casServers_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_53_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_53_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_53_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_53_io_addressIn_ready),
		.io_addressOut_valid(_casServers_53_io_addressOut_valid),
		.io_addressOut_bits(_casServers_53_io_addressOut_bits)
	);
	AllocatorClient casServers_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_54_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_54_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_54_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_54_io_addressIn_ready),
		.io_addressOut_valid(_casServers_54_io_addressOut_valid),
		.io_addressOut_bits(_casServers_54_io_addressOut_bits)
	);
	AllocatorClient casServers_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_55_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_55_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_55_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_55_io_addressIn_ready),
		.io_addressOut_valid(_casServers_55_io_addressOut_valid),
		.io_addressOut_bits(_casServers_55_io_addressOut_bits)
	);
	AllocatorClient casServers_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_56_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_56_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_56_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_56_io_addressIn_ready),
		.io_addressOut_valid(_casServers_56_io_addressOut_valid),
		.io_addressOut_bits(_casServers_56_io_addressOut_bits)
	);
	AllocatorClient casServers_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_57_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_57_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_57_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_57_io_addressIn_ready),
		.io_addressOut_valid(_casServers_57_io_addressOut_valid),
		.io_addressOut_bits(_casServers_57_io_addressOut_bits)
	);
	AllocatorClient casServers_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_58_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_58_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_58_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_58_io_addressIn_ready),
		.io_addressOut_valid(_casServers_58_io_addressOut_valid),
		.io_addressOut_bits(_casServers_58_io_addressOut_bits)
	);
	AllocatorClient casServers_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_59_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_59_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_59_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_59_io_addressIn_ready),
		.io_addressOut_valid(_casServers_59_io_addressOut_valid),
		.io_addressOut_bits(_casServers_59_io_addressOut_bits)
	);
	AllocatorClient casServers_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_60_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_60_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_60_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_60_io_addressIn_ready),
		.io_addressOut_valid(_casServers_60_io_addressOut_valid),
		.io_addressOut_bits(_casServers_60_io_addressOut_bits)
	);
	AllocatorClient casServers_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_61_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_61_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_61_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_61_io_addressIn_ready),
		.io_addressOut_valid(_casServers_61_io_addressOut_valid),
		.io_addressOut_bits(_casServers_61_io_addressOut_bits)
	);
	AllocatorClient casServers_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_62_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_62_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_62_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_62_io_addressIn_ready),
		.io_addressOut_valid(_casServers_62_io_addressOut_valid),
		.io_addressOut_bits(_casServers_62_io_addressOut_bits)
	);
	AllocatorClient casServers_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_casServers_63_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_63_io_casAddressOut_valid),
		.io_addressIn_bits(_networkUnits_63_io_casAddressOut_bits),
		.io_addressOut_ready(_queues_63_io_addressIn_ready),
		.io_addressOut_valid(_casServers_63_io_addressOut_valid),
		.io_addressOut_bits(_casServers_63_io_addressOut_bits)
	);
	AllocatorBuffer queues_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_0_io_addressIn_ready),
		.io_addressIn_valid(_casServers_0_io_addressOut_valid),
		.io_addressIn_bits(_casServers_0_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_0_ready),
		.io_addressOut_valid(io_connPE_0_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_1_io_addressIn_ready),
		.io_addressIn_valid(_casServers_1_io_addressOut_valid),
		.io_addressIn_bits(_casServers_1_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_1_ready),
		.io_addressOut_valid(io_connPE_1_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_2_io_addressIn_ready),
		.io_addressIn_valid(_casServers_2_io_addressOut_valid),
		.io_addressIn_bits(_casServers_2_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_2_ready),
		.io_addressOut_valid(io_connPE_2_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_3_io_addressIn_ready),
		.io_addressIn_valid(_casServers_3_io_addressOut_valid),
		.io_addressIn_bits(_casServers_3_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_3_ready),
		.io_addressOut_valid(io_connPE_3_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_4_io_addressIn_ready),
		.io_addressIn_valid(_casServers_4_io_addressOut_valid),
		.io_addressIn_bits(_casServers_4_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_4_ready),
		.io_addressOut_valid(io_connPE_4_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_5_io_addressIn_ready),
		.io_addressIn_valid(_casServers_5_io_addressOut_valid),
		.io_addressIn_bits(_casServers_5_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_5_ready),
		.io_addressOut_valid(io_connPE_5_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_6_io_addressIn_ready),
		.io_addressIn_valid(_casServers_6_io_addressOut_valid),
		.io_addressIn_bits(_casServers_6_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_6_ready),
		.io_addressOut_valid(io_connPE_6_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_7_io_addressIn_ready),
		.io_addressIn_valid(_casServers_7_io_addressOut_valid),
		.io_addressIn_bits(_casServers_7_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_7_ready),
		.io_addressOut_valid(io_connPE_7_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_8_io_addressIn_ready),
		.io_addressIn_valid(_casServers_8_io_addressOut_valid),
		.io_addressIn_bits(_casServers_8_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_8_ready),
		.io_addressOut_valid(io_connPE_8_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_9_io_addressIn_ready),
		.io_addressIn_valid(_casServers_9_io_addressOut_valid),
		.io_addressIn_bits(_casServers_9_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_9_ready),
		.io_addressOut_valid(io_connPE_9_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_10_io_addressIn_ready),
		.io_addressIn_valid(_casServers_10_io_addressOut_valid),
		.io_addressIn_bits(_casServers_10_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_10_ready),
		.io_addressOut_valid(io_connPE_10_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_11_io_addressIn_ready),
		.io_addressIn_valid(_casServers_11_io_addressOut_valid),
		.io_addressIn_bits(_casServers_11_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_11_ready),
		.io_addressOut_valid(io_connPE_11_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_12_io_addressIn_ready),
		.io_addressIn_valid(_casServers_12_io_addressOut_valid),
		.io_addressIn_bits(_casServers_12_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_12_ready),
		.io_addressOut_valid(io_connPE_12_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_13_io_addressIn_ready),
		.io_addressIn_valid(_casServers_13_io_addressOut_valid),
		.io_addressIn_bits(_casServers_13_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_13_ready),
		.io_addressOut_valid(io_connPE_13_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_14_io_addressIn_ready),
		.io_addressIn_valid(_casServers_14_io_addressOut_valid),
		.io_addressIn_bits(_casServers_14_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_14_ready),
		.io_addressOut_valid(io_connPE_14_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_15_io_addressIn_ready),
		.io_addressIn_valid(_casServers_15_io_addressOut_valid),
		.io_addressIn_bits(_casServers_15_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_15_ready),
		.io_addressOut_valid(io_connPE_15_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_16_io_addressIn_ready),
		.io_addressIn_valid(_casServers_16_io_addressOut_valid),
		.io_addressIn_bits(_casServers_16_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_16_ready),
		.io_addressOut_valid(io_connPE_16_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_17_io_addressIn_ready),
		.io_addressIn_valid(_casServers_17_io_addressOut_valid),
		.io_addressIn_bits(_casServers_17_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_17_ready),
		.io_addressOut_valid(io_connPE_17_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_18_io_addressIn_ready),
		.io_addressIn_valid(_casServers_18_io_addressOut_valid),
		.io_addressIn_bits(_casServers_18_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_18_ready),
		.io_addressOut_valid(io_connPE_18_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_19_io_addressIn_ready),
		.io_addressIn_valid(_casServers_19_io_addressOut_valid),
		.io_addressIn_bits(_casServers_19_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_19_ready),
		.io_addressOut_valid(io_connPE_19_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_20_io_addressIn_ready),
		.io_addressIn_valid(_casServers_20_io_addressOut_valid),
		.io_addressIn_bits(_casServers_20_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_20_ready),
		.io_addressOut_valid(io_connPE_20_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_21_io_addressIn_ready),
		.io_addressIn_valid(_casServers_21_io_addressOut_valid),
		.io_addressIn_bits(_casServers_21_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_21_ready),
		.io_addressOut_valid(io_connPE_21_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_22_io_addressIn_ready),
		.io_addressIn_valid(_casServers_22_io_addressOut_valid),
		.io_addressIn_bits(_casServers_22_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_22_ready),
		.io_addressOut_valid(io_connPE_22_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_23_io_addressIn_ready),
		.io_addressIn_valid(_casServers_23_io_addressOut_valid),
		.io_addressIn_bits(_casServers_23_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_23_ready),
		.io_addressOut_valid(io_connPE_23_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_24_io_addressIn_ready),
		.io_addressIn_valid(_casServers_24_io_addressOut_valid),
		.io_addressIn_bits(_casServers_24_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_24_ready),
		.io_addressOut_valid(io_connPE_24_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_25_io_addressIn_ready),
		.io_addressIn_valid(_casServers_25_io_addressOut_valid),
		.io_addressIn_bits(_casServers_25_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_25_ready),
		.io_addressOut_valid(io_connPE_25_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_26_io_addressIn_ready),
		.io_addressIn_valid(_casServers_26_io_addressOut_valid),
		.io_addressIn_bits(_casServers_26_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_26_ready),
		.io_addressOut_valid(io_connPE_26_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_27_io_addressIn_ready),
		.io_addressIn_valid(_casServers_27_io_addressOut_valid),
		.io_addressIn_bits(_casServers_27_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_27_ready),
		.io_addressOut_valid(io_connPE_27_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_28_io_addressIn_ready),
		.io_addressIn_valid(_casServers_28_io_addressOut_valid),
		.io_addressIn_bits(_casServers_28_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_28_ready),
		.io_addressOut_valid(io_connPE_28_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_29_io_addressIn_ready),
		.io_addressIn_valid(_casServers_29_io_addressOut_valid),
		.io_addressIn_bits(_casServers_29_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_29_ready),
		.io_addressOut_valid(io_connPE_29_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_30_io_addressIn_ready),
		.io_addressIn_valid(_casServers_30_io_addressOut_valid),
		.io_addressIn_bits(_casServers_30_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_30_ready),
		.io_addressOut_valid(io_connPE_30_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_31_io_addressIn_ready),
		.io_addressIn_valid(_casServers_31_io_addressOut_valid),
		.io_addressIn_bits(_casServers_31_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_31_ready),
		.io_addressOut_valid(io_connPE_31_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_32_io_addressIn_ready),
		.io_addressIn_valid(_casServers_32_io_addressOut_valid),
		.io_addressIn_bits(_casServers_32_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_32_ready),
		.io_addressOut_valid(io_connPE_32_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_33_io_addressIn_ready),
		.io_addressIn_valid(_casServers_33_io_addressOut_valid),
		.io_addressIn_bits(_casServers_33_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_33_ready),
		.io_addressOut_valid(io_connPE_33_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_34_io_addressIn_ready),
		.io_addressIn_valid(_casServers_34_io_addressOut_valid),
		.io_addressIn_bits(_casServers_34_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_34_ready),
		.io_addressOut_valid(io_connPE_34_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_35_io_addressIn_ready),
		.io_addressIn_valid(_casServers_35_io_addressOut_valid),
		.io_addressIn_bits(_casServers_35_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_35_ready),
		.io_addressOut_valid(io_connPE_35_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_36_io_addressIn_ready),
		.io_addressIn_valid(_casServers_36_io_addressOut_valid),
		.io_addressIn_bits(_casServers_36_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_36_ready),
		.io_addressOut_valid(io_connPE_36_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_37_io_addressIn_ready),
		.io_addressIn_valid(_casServers_37_io_addressOut_valid),
		.io_addressIn_bits(_casServers_37_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_37_ready),
		.io_addressOut_valid(io_connPE_37_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_38_io_addressIn_ready),
		.io_addressIn_valid(_casServers_38_io_addressOut_valid),
		.io_addressIn_bits(_casServers_38_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_38_ready),
		.io_addressOut_valid(io_connPE_38_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_39_io_addressIn_ready),
		.io_addressIn_valid(_casServers_39_io_addressOut_valid),
		.io_addressIn_bits(_casServers_39_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_39_ready),
		.io_addressOut_valid(io_connPE_39_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_40_io_addressIn_ready),
		.io_addressIn_valid(_casServers_40_io_addressOut_valid),
		.io_addressIn_bits(_casServers_40_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_40_ready),
		.io_addressOut_valid(io_connPE_40_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_41_io_addressIn_ready),
		.io_addressIn_valid(_casServers_41_io_addressOut_valid),
		.io_addressIn_bits(_casServers_41_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_41_ready),
		.io_addressOut_valid(io_connPE_41_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_42_io_addressIn_ready),
		.io_addressIn_valid(_casServers_42_io_addressOut_valid),
		.io_addressIn_bits(_casServers_42_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_42_ready),
		.io_addressOut_valid(io_connPE_42_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_43_io_addressIn_ready),
		.io_addressIn_valid(_casServers_43_io_addressOut_valid),
		.io_addressIn_bits(_casServers_43_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_43_ready),
		.io_addressOut_valid(io_connPE_43_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_44_io_addressIn_ready),
		.io_addressIn_valid(_casServers_44_io_addressOut_valid),
		.io_addressIn_bits(_casServers_44_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_44_ready),
		.io_addressOut_valid(io_connPE_44_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_45_io_addressIn_ready),
		.io_addressIn_valid(_casServers_45_io_addressOut_valid),
		.io_addressIn_bits(_casServers_45_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_45_ready),
		.io_addressOut_valid(io_connPE_45_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_46_io_addressIn_ready),
		.io_addressIn_valid(_casServers_46_io_addressOut_valid),
		.io_addressIn_bits(_casServers_46_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_46_ready),
		.io_addressOut_valid(io_connPE_46_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_47_io_addressIn_ready),
		.io_addressIn_valid(_casServers_47_io_addressOut_valid),
		.io_addressIn_bits(_casServers_47_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_47_ready),
		.io_addressOut_valid(io_connPE_47_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_48_io_addressIn_ready),
		.io_addressIn_valid(_casServers_48_io_addressOut_valid),
		.io_addressIn_bits(_casServers_48_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_48_ready),
		.io_addressOut_valid(io_connPE_48_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_49_io_addressIn_ready),
		.io_addressIn_valid(_casServers_49_io_addressOut_valid),
		.io_addressIn_bits(_casServers_49_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_49_ready),
		.io_addressOut_valid(io_connPE_49_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_50_io_addressIn_ready),
		.io_addressIn_valid(_casServers_50_io_addressOut_valid),
		.io_addressIn_bits(_casServers_50_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_50_ready),
		.io_addressOut_valid(io_connPE_50_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_51_io_addressIn_ready),
		.io_addressIn_valid(_casServers_51_io_addressOut_valid),
		.io_addressIn_bits(_casServers_51_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_51_ready),
		.io_addressOut_valid(io_connPE_51_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_52_io_addressIn_ready),
		.io_addressIn_valid(_casServers_52_io_addressOut_valid),
		.io_addressIn_bits(_casServers_52_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_52_ready),
		.io_addressOut_valid(io_connPE_52_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_53_io_addressIn_ready),
		.io_addressIn_valid(_casServers_53_io_addressOut_valid),
		.io_addressIn_bits(_casServers_53_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_53_ready),
		.io_addressOut_valid(io_connPE_53_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_54_io_addressIn_ready),
		.io_addressIn_valid(_casServers_54_io_addressOut_valid),
		.io_addressIn_bits(_casServers_54_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_54_ready),
		.io_addressOut_valid(io_connPE_54_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_55_io_addressIn_ready),
		.io_addressIn_valid(_casServers_55_io_addressOut_valid),
		.io_addressIn_bits(_casServers_55_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_55_ready),
		.io_addressOut_valid(io_connPE_55_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_56_io_addressIn_ready),
		.io_addressIn_valid(_casServers_56_io_addressOut_valid),
		.io_addressIn_bits(_casServers_56_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_56_ready),
		.io_addressOut_valid(io_connPE_56_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_57_io_addressIn_ready),
		.io_addressIn_valid(_casServers_57_io_addressOut_valid),
		.io_addressIn_bits(_casServers_57_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_57_ready),
		.io_addressOut_valid(io_connPE_57_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_58_io_addressIn_ready),
		.io_addressIn_valid(_casServers_58_io_addressOut_valid),
		.io_addressIn_bits(_casServers_58_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_58_ready),
		.io_addressOut_valid(io_connPE_58_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_59_io_addressIn_ready),
		.io_addressIn_valid(_casServers_59_io_addressOut_valid),
		.io_addressIn_bits(_casServers_59_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_59_ready),
		.io_addressOut_valid(io_connPE_59_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_60_io_addressIn_ready),
		.io_addressIn_valid(_casServers_60_io_addressOut_valid),
		.io_addressIn_bits(_casServers_60_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_60_ready),
		.io_addressOut_valid(io_connPE_60_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_61_io_addressIn_ready),
		.io_addressIn_valid(_casServers_61_io_addressOut_valid),
		.io_addressIn_bits(_casServers_61_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_61_ready),
		.io_addressOut_valid(io_connPE_61_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_62_io_addressIn_ready),
		.io_addressIn_valid(_casServers_62_io_addressOut_valid),
		.io_addressIn_bits(_casServers_62_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_62_ready),
		.io_addressOut_valid(io_connPE_62_valid),
		.io_addressOut_bits()
	);
	AllocatorBuffer queues_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_queues_63_io_addressIn_ready),
		.io_addressIn_valid(_casServers_63_io_addressOut_valid),
		.io_addressIn_bits(_casServers_63_io_addressOut_bits),
		.io_addressOut_ready(io_connPE_63_ready),
		.io_addressOut_valid(io_connPE_63_valid),
		.io_addressOut_bits()
	);
endmodule
module AllocatorServer (
	clock,
	reset,
	io_dataOut_ready,
	io_dataOut_valid,
	io_dataOut_bits,
	io_axi_mgmt_ar_ready,
	io_axi_mgmt_ar_valid,
	io_axi_mgmt_ar_bits_addr,
	io_axi_mgmt_ar_bits_prot,
	io_axi_mgmt_r_ready,
	io_axi_mgmt_r_valid,
	io_axi_mgmt_r_bits_data,
	io_axi_mgmt_r_bits_resp,
	io_axi_mgmt_aw_ready,
	io_axi_mgmt_aw_valid,
	io_axi_mgmt_aw_bits_addr,
	io_axi_mgmt_aw_bits_prot,
	io_axi_mgmt_w_ready,
	io_axi_mgmt_w_valid,
	io_axi_mgmt_w_bits_data,
	io_axi_mgmt_w_bits_strb,
	io_axi_mgmt_b_ready,
	io_axi_mgmt_b_valid,
	io_axi_mgmt_b_bits_resp,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits
);
	input clock;
	input reset;
	input io_dataOut_ready;
	output wire io_dataOut_valid;
	output wire [63:0] io_dataOut_bits;
	output wire io_axi_mgmt_ar_ready;
	input io_axi_mgmt_ar_valid;
	input [5:0] io_axi_mgmt_ar_bits_addr;
	input [2:0] io_axi_mgmt_ar_bits_prot;
	input io_axi_mgmt_r_ready;
	output wire io_axi_mgmt_r_valid;
	output wire [63:0] io_axi_mgmt_r_bits_data;
	output wire [1:0] io_axi_mgmt_r_bits_resp;
	output wire io_axi_mgmt_aw_ready;
	input io_axi_mgmt_aw_valid;
	input [5:0] io_axi_mgmt_aw_bits_addr;
	input [2:0] io_axi_mgmt_aw_bits_prot;
	output wire io_axi_mgmt_w_ready;
	input io_axi_mgmt_w_valid;
	input [63:0] io_axi_mgmt_w_bits_data;
	input [7:0] io_axi_mgmt_w_bits_strb;
	input io_axi_mgmt_b_ready;
	output wire io_axi_mgmt_b_valid;
	output wire [1:0] io_axi_mgmt_b_bits_resp;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [63:0] io_read_data_bits;
	wire _wrRespQueue__io_enq_ready;
	wire _wrRespQueue__io_deq_valid;
	wire _wrReqData__deq_q_io_enq_ready;
	wire _wrReqData__deq_q_io_deq_valid;
	wire [63:0] _wrReqData__deq_q_io_deq_bits_data;
	wire [7:0] _wrReqData__deq_q_io_deq_bits_strb;
	wire _wrReq__deq_q_io_enq_ready;
	wire _wrReq__deq_q_io_deq_valid;
	wire [5:0] _wrReq__deq_q_io_deq_bits_addr;
	wire _rdRespQueue__io_enq_ready;
	wire _rdRespQueue__io_deq_valid;
	wire [63:0] _rdRespQueue__io_deq_bits_data;
	wire [1:0] _rdRespQueue__io_deq_bits_resp;
	wire _rdReq__deq_q_io_enq_ready;
	wire _rdReq__deq_q_io_deq_valid;
	wire [5:0] _rdReq__deq_q_io_deq_bits_addr;
	wire _s_axil__sinkBuffer_1_io_enq_ready;
	wire _s_axil__sourceBuffer_2_io_deq_valid;
	wire [63:0] _s_axil__sourceBuffer_2_io_deq_bits_data;
	wire [7:0] _s_axil__sourceBuffer_2_io_deq_bits_strb;
	wire _s_axil__sourceBuffer_1_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_1_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_1_io_deq_bits_prot;
	wire _s_axil__sinkBuffer_io_enq_ready;
	wire _s_axil__sourceBuffer_io_deq_valid;
	wire [5:0] _s_axil__sourceBuffer_io_deq_bits_addr;
	wire [2:0] _s_axil__sourceBuffer_io_deq_bits_prot;
	wire rdReq = _rdReq__deq_q_io_deq_valid & _rdRespQueue__io_enq_ready;
	wire wrReq = (_wrReq__deq_q_io_deq_valid & _wrReqData__deq_q_io_deq_valid) & _wrRespQueue__io_enq_ready;
	reg [63:0] rAddr;
	reg [63:0] rPause;
	reg [63:0] avaialbleSize;
	reg [2:0] stateReg;
	reg [63:0] continuationsRegisters_0;
	reg [63:0] continuationsRegisters_1;
	reg [63:0] continuationsRegisters_2;
	reg [63:0] continuationsRegisters_3;
	reg [63:0] continuationsRegisters_4;
	reg [63:0] continuationsRegisters_5;
	reg [63:0] continuationsRegisters_6;
	reg [63:0] continuationsRegisters_7;
	reg [63:0] continuationsRegisters_8;
	reg [63:0] continuationsRegisters_9;
	reg [63:0] continuationsRegisters_10;
	reg [63:0] continuationsRegisters_11;
	reg [63:0] continuationsRegisters_12;
	reg [63:0] continuationsRegisters_13;
	reg [63:0] continuationsRegisters_14;
	reg [63:0] continuationsRegisters_15;
	reg [3:0] burstCounter;
	wire io_read_address_valid_0 = stateReg == 3'h1;
	wire _GEN = stateReg == 3'h2;
	wire _GEN_0 = stateReg == 3'h3;
	wire [1023:0] _GEN_1 = {continuationsRegisters_15, continuationsRegisters_14, continuationsRegisters_13, continuationsRegisters_12, continuationsRegisters_11, continuationsRegisters_10, continuationsRegisters_9, continuationsRegisters_8, continuationsRegisters_7, continuationsRegisters_6, continuationsRegisters_5, continuationsRegisters_4, continuationsRegisters_3, continuationsRegisters_2, continuationsRegisters_1, continuationsRegisters_0};
	always @(posedge clock)
		if (reset) begin
			rAddr <= 64'h0000000000000000;
			rPause <= 64'h0000000000000000;
			avaialbleSize <= 64'h0000000000000000;
			stateReg <= 3'h0;
			continuationsRegisters_0 <= 64'h0000000000000000;
			continuationsRegisters_1 <= 64'h0000000000000000;
			continuationsRegisters_2 <= 64'h0000000000000000;
			continuationsRegisters_3 <= 64'h0000000000000000;
			continuationsRegisters_4 <= 64'h0000000000000000;
			continuationsRegisters_5 <= 64'h0000000000000000;
			continuationsRegisters_6 <= 64'h0000000000000000;
			continuationsRegisters_7 <= 64'h0000000000000000;
			continuationsRegisters_8 <= 64'h0000000000000000;
			continuationsRegisters_9 <= 64'h0000000000000000;
			continuationsRegisters_10 <= 64'h0000000000000000;
			continuationsRegisters_11 <= 64'h0000000000000000;
			continuationsRegisters_12 <= 64'h0000000000000000;
			continuationsRegisters_13 <= 64'h0000000000000000;
			continuationsRegisters_14 <= 64'h0000000000000000;
			continuationsRegisters_15 <= 64'h0000000000000000;
			burstCounter <= 4'hf;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_2;
			reg _GEN_3;
			reg _GEN_4;
			reg _GEN_5;
			_GEN_2 = stateReg == 3'h0;
			_GEN_3 = burstCounter == 4'h0;
			_GEN_4 = _GEN_2 | io_read_address_valid_0;
			_GEN_5 = _GEN_3 & io_read_data_valid;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h1))
				rAddr <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rAddr[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rAddr[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rAddr[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rAddr[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rAddr[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rAddr[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rAddr[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rAddr[7:0])};
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h0))
				rPause <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : rPause[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : rPause[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : rPause[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : rPause[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : rPause[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : rPause[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : rPause[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : rPause[7:0])};
			else if (~_GEN_2 | (|avaialbleSize[63:4]))
				;
			else
				rPause <= 64'hffffffffffffffff;
			if (wrReq & (_wrReq__deq_q_io_deq_bits_addr[5:3] == 3'h2))
				avaialbleSize <= {(_wrReqData__deq_q_io_deq_bits_strb[7] ? _wrReqData__deq_q_io_deq_bits_data[63:56] : avaialbleSize[63:56]), (_wrReqData__deq_q_io_deq_bits_strb[6] ? _wrReqData__deq_q_io_deq_bits_data[55:48] : avaialbleSize[55:48]), (_wrReqData__deq_q_io_deq_bits_strb[5] ? _wrReqData__deq_q_io_deq_bits_data[47:40] : avaialbleSize[47:40]), (_wrReqData__deq_q_io_deq_bits_strb[4] ? _wrReqData__deq_q_io_deq_bits_data[39:32] : avaialbleSize[39:32]), (_wrReqData__deq_q_io_deq_bits_strb[3] ? _wrReqData__deq_q_io_deq_bits_data[31:24] : avaialbleSize[31:24]), (_wrReqData__deq_q_io_deq_bits_strb[2] ? _wrReqData__deq_q_io_deq_bits_data[23:16] : avaialbleSize[23:16]), (_wrReqData__deq_q_io_deq_bits_strb[1] ? _wrReqData__deq_q_io_deq_bits_data[15:8] : avaialbleSize[15:8]), (_wrReqData__deq_q_io_deq_bits_strb[0] ? _wrReqData__deq_q_io_deq_bits_data[7:0] : avaialbleSize[7:0])};
			else if (_GEN_4 | ~_GEN)
				;
			else if (_GEN_5)
				avaialbleSize <= avaialbleSize - 64'h0000000000000001;
			else if (io_read_data_valid)
				avaialbleSize <= avaialbleSize - 64'h0000000000000001;
			if (_GEN_2)
				stateReg <= (|avaialbleSize[63:4] ? 3'h1 : 3'h4);
			else if (io_read_address_valid_0) begin
				if (io_read_address_ready) begin
					stateReg <= 3'h2;
					burstCounter <= 4'hf;
				end
			end
			else if (_GEN) begin
				if (_GEN_5) begin
					stateReg <= 3'h3;
					burstCounter <= 4'hf;
				end
				else if (io_read_data_valid)
					burstCounter <= burstCounter - 4'h1;
			end
			else begin
				if ((_GEN_0 ? _GEN_3 & io_dataOut_ready : (stateReg == 3'h4) & (rPause == 64'h0000000000000000)))
					stateReg <= 3'h0;
				if (_GEN_0 & io_dataOut_ready)
					burstCounter <= burstCounter - 4'h1;
			end
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & _GEN_3))
				;
			else
				continuationsRegisters_0 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h1)))
				;
			else
				continuationsRegisters_1 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h2)))
				;
			else
				continuationsRegisters_2 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h3)))
				;
			else
				continuationsRegisters_3 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h4)))
				;
			else
				continuationsRegisters_4 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h5)))
				;
			else
				continuationsRegisters_5 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h6)))
				;
			else
				continuationsRegisters_6 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h7)))
				;
			else
				continuationsRegisters_7 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h8)))
				;
			else
				continuationsRegisters_8 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'h9)))
				;
			else
				continuationsRegisters_9 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'ha)))
				;
			else
				continuationsRegisters_10 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'hb)))
				;
			else
				continuationsRegisters_11 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'hc)))
				;
			else
				continuationsRegisters_12 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'hd)))
				;
			else
				continuationsRegisters_13 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (burstCounter == 4'he)))
				;
			else
				continuationsRegisters_14 <= io_read_data_bits;
			if (_GEN_4 | ~((_GEN & io_read_data_valid) & (&burstCounter)))
				;
			else
				continuationsRegisters_15 <= io_read_data_bits;
		end
	Queue2_AddressChannel_2 s_axil__sourceBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_ar_ready),
		.io_enq_valid(io_axi_mgmt_ar_valid),
		.io_enq_bits_addr(io_axi_mgmt_ar_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_ar_bits_prot),
		.io_deq_ready(_rdReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot)
	);
	Queue2_ReadDataChannel s_axil__sinkBuffer(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_enq_valid(_rdRespQueue__io_deq_valid),
		.io_enq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_enq_bits_resp(_rdRespQueue__io_deq_bits_resp),
		.io_deq_ready(io_axi_mgmt_r_ready),
		.io_deq_valid(io_axi_mgmt_r_valid),
		.io_deq_bits_data(io_axi_mgmt_r_bits_data),
		.io_deq_bits_resp(io_axi_mgmt_r_bits_resp)
	);
	Queue2_AddressChannel_2 s_axil__sourceBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_aw_ready),
		.io_enq_valid(io_axi_mgmt_aw_valid),
		.io_enq_bits_addr(io_axi_mgmt_aw_bits_addr),
		.io_enq_bits_prot(io_axi_mgmt_aw_bits_prot),
		.io_deq_ready(_wrReq__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_deq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_deq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot)
	);
	Queue2_WriteDataChannel s_axil__sourceBuffer_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_axi_mgmt_w_ready),
		.io_enq_valid(io_axi_mgmt_w_valid),
		.io_enq_bits_data(io_axi_mgmt_w_bits_data),
		.io_enq_bits_strb(io_axi_mgmt_w_bits_strb),
		.io_deq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_deq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_deq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_deq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb)
	);
	Queue2_WriteResponseChannel s_axil__sinkBuffer_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_enq_valid(_wrRespQueue__io_deq_valid),
		.io_enq_bits_resp(2'h0),
		.io_deq_ready(io_axi_mgmt_b_ready),
		.io_deq_valid(io_axi_mgmt_b_valid),
		.io_deq_bits_resp(io_axi_mgmt_b_bits_resp)
	);
	Queue1_AddressChannel rdReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_io_deq_bits_prot),
		.io_deq_ready(rdReq),
		.io_deq_valid(_rdReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_rdReq__deq_q_io_deq_bits_addr)
	);
	Queue1_ReadDataChannel rdRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_rdRespQueue__io_enq_ready),
		.io_enq_valid(rdReq),
		.io_enq_bits_data((_rdReq__deq_q_io_deq_bits_addr[5:3] == 3'h2 ? avaialbleSize : (_rdReq__deq_q_io_deq_bits_addr[5:3] == 3'h1 ? rAddr : (_rdReq__deq_q_io_deq_bits_addr[5:3] == 3'h0 ? rPause : 64'hffffffffffffffff)))),
		.io_deq_ready(_s_axil__sinkBuffer_io_enq_ready),
		.io_deq_valid(_rdRespQueue__io_deq_valid),
		.io_deq_bits_data(_rdRespQueue__io_deq_bits_data),
		.io_deq_bits_resp(_rdRespQueue__io_deq_bits_resp)
	);
	Queue1_AddressChannel wrReq__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReq__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_1_io_deq_valid),
		.io_enq_bits_addr(_s_axil__sourceBuffer_1_io_deq_bits_addr),
		.io_enq_bits_prot(_s_axil__sourceBuffer_1_io_deq_bits_prot),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReq__deq_q_io_deq_valid),
		.io_deq_bits_addr(_wrReq__deq_q_io_deq_bits_addr)
	);
	Queue1_WriteDataChannel wrReqData__deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrReqData__deq_q_io_enq_ready),
		.io_enq_valid(_s_axil__sourceBuffer_2_io_deq_valid),
		.io_enq_bits_data(_s_axil__sourceBuffer_2_io_deq_bits_data),
		.io_enq_bits_strb(_s_axil__sourceBuffer_2_io_deq_bits_strb),
		.io_deq_ready(wrReq),
		.io_deq_valid(_wrReqData__deq_q_io_deq_valid),
		.io_deq_bits_data(_wrReqData__deq_q_io_deq_bits_data),
		.io_deq_bits_strb(_wrReqData__deq_q_io_deq_bits_strb)
	);
	Queue1_WriteResponseChannel wrRespQueue_(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_wrRespQueue__io_enq_ready),
		.io_enq_valid(wrReq),
		.io_deq_ready(_s_axil__sinkBuffer_1_io_enq_ready),
		.io_deq_valid(_wrRespQueue__io_deq_valid)
	);
	assign io_dataOut_valid = ~(io_read_address_valid_0 | _GEN) & _GEN_0;
	assign io_dataOut_bits = _GEN_1[burstCounter * 64+:64];
	assign io_read_address_valid = io_read_address_valid_0;
	assign io_read_address_bits = rAddr + {avaialbleSize[60:0] - 61'h0000000000000010, 3'h0};
	assign io_read_data_ready = ~io_read_address_valid_0 & _GEN;
endmodule
module RVtoAXIBridge_2 (
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data
);
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [63:0] io_read_data_bits;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire axi_r_ready;
	input axi_r_valid;
	input [63:0] axi_r_bits_data;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_r_ready = io_read_data_ready;
endmodule
module AxisDownscaler_80 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataOut_TREADY,
	io_dataOut_TVALID
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	reg writeCounter;
	reg stateReg;
	always @(posedge clock)
		if (reset) begin
			writeCounter <= 1'h0;
			stateReg <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg _GEN;
			_GEN = io_dataOut_TREADY & ~writeCounter;
			if (stateReg) begin
				if (stateReg & _GEN)
					writeCounter <= writeCounter - 1'h1;
			end
			else
				writeCounter <= ~io_dataIn_TVALID & writeCounter;
			stateReg <= ((~stateReg | _GEN) | ~(io_dataOut_TREADY & writeCounter)) & stateReg;
		end
	assign io_dataIn_TREADY = ~stateReg;
	assign io_dataOut_TVALID = stateReg;
endmodule
module AxisDataWidthConverter_144 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataOut_TREADY,
	io_dataOut_TVALID
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	AxisDownscaler_80 downScaler(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_dataIn_TREADY),
		.io_dataIn_TVALID(io_dataIn_TVALID),
		.io_dataOut_TREADY(io_dataOut_TREADY),
		.io_dataOut_TVALID(io_dataOut_TVALID)
	);
endmodule
module Allocator (
	clock,
	reset,
	io_export_closureOut_0_TREADY,
	io_export_closureOut_0_TVALID,
	io_export_closureOut_1_TREADY,
	io_export_closureOut_1_TVALID,
	io_export_closureOut_2_TREADY,
	io_export_closureOut_2_TVALID,
	io_export_closureOut_3_TREADY,
	io_export_closureOut_3_TVALID,
	io_export_closureOut_4_TREADY,
	io_export_closureOut_4_TVALID,
	io_export_closureOut_5_TREADY,
	io_export_closureOut_5_TVALID,
	io_export_closureOut_6_TREADY,
	io_export_closureOut_6_TVALID,
	io_export_closureOut_7_TREADY,
	io_export_closureOut_7_TVALID,
	io_export_closureOut_8_TREADY,
	io_export_closureOut_8_TVALID,
	io_export_closureOut_9_TREADY,
	io_export_closureOut_9_TVALID,
	io_export_closureOut_10_TREADY,
	io_export_closureOut_10_TVALID,
	io_export_closureOut_11_TREADY,
	io_export_closureOut_11_TVALID,
	io_export_closureOut_12_TREADY,
	io_export_closureOut_12_TVALID,
	io_export_closureOut_13_TREADY,
	io_export_closureOut_13_TVALID,
	io_export_closureOut_14_TREADY,
	io_export_closureOut_14_TVALID,
	io_export_closureOut_15_TREADY,
	io_export_closureOut_15_TVALID,
	io_export_closureOut_16_TREADY,
	io_export_closureOut_16_TVALID,
	io_export_closureOut_17_TREADY,
	io_export_closureOut_17_TVALID,
	io_export_closureOut_18_TREADY,
	io_export_closureOut_18_TVALID,
	io_export_closureOut_19_TREADY,
	io_export_closureOut_19_TVALID,
	io_export_closureOut_20_TREADY,
	io_export_closureOut_20_TVALID,
	io_export_closureOut_21_TREADY,
	io_export_closureOut_21_TVALID,
	io_export_closureOut_22_TREADY,
	io_export_closureOut_22_TVALID,
	io_export_closureOut_23_TREADY,
	io_export_closureOut_23_TVALID,
	io_export_closureOut_24_TREADY,
	io_export_closureOut_24_TVALID,
	io_export_closureOut_25_TREADY,
	io_export_closureOut_25_TVALID,
	io_export_closureOut_26_TREADY,
	io_export_closureOut_26_TVALID,
	io_export_closureOut_27_TREADY,
	io_export_closureOut_27_TVALID,
	io_export_closureOut_28_TREADY,
	io_export_closureOut_28_TVALID,
	io_export_closureOut_29_TREADY,
	io_export_closureOut_29_TVALID,
	io_export_closureOut_30_TREADY,
	io_export_closureOut_30_TVALID,
	io_export_closureOut_31_TREADY,
	io_export_closureOut_31_TVALID,
	io_export_closureOut_32_TREADY,
	io_export_closureOut_32_TVALID,
	io_export_closureOut_33_TREADY,
	io_export_closureOut_33_TVALID,
	io_export_closureOut_34_TREADY,
	io_export_closureOut_34_TVALID,
	io_export_closureOut_35_TREADY,
	io_export_closureOut_35_TVALID,
	io_export_closureOut_36_TREADY,
	io_export_closureOut_36_TVALID,
	io_export_closureOut_37_TREADY,
	io_export_closureOut_37_TVALID,
	io_export_closureOut_38_TREADY,
	io_export_closureOut_38_TVALID,
	io_export_closureOut_39_TREADY,
	io_export_closureOut_39_TVALID,
	io_export_closureOut_40_TREADY,
	io_export_closureOut_40_TVALID,
	io_export_closureOut_41_TREADY,
	io_export_closureOut_41_TVALID,
	io_export_closureOut_42_TREADY,
	io_export_closureOut_42_TVALID,
	io_export_closureOut_43_TREADY,
	io_export_closureOut_43_TVALID,
	io_export_closureOut_44_TREADY,
	io_export_closureOut_44_TVALID,
	io_export_closureOut_45_TREADY,
	io_export_closureOut_45_TVALID,
	io_export_closureOut_46_TREADY,
	io_export_closureOut_46_TVALID,
	io_export_closureOut_47_TREADY,
	io_export_closureOut_47_TVALID,
	io_export_closureOut_48_TREADY,
	io_export_closureOut_48_TVALID,
	io_export_closureOut_49_TREADY,
	io_export_closureOut_49_TVALID,
	io_export_closureOut_50_TREADY,
	io_export_closureOut_50_TVALID,
	io_export_closureOut_51_TREADY,
	io_export_closureOut_51_TVALID,
	io_export_closureOut_52_TREADY,
	io_export_closureOut_52_TVALID,
	io_export_closureOut_53_TREADY,
	io_export_closureOut_53_TVALID,
	io_export_closureOut_54_TREADY,
	io_export_closureOut_54_TVALID,
	io_export_closureOut_55_TREADY,
	io_export_closureOut_55_TVALID,
	io_export_closureOut_56_TREADY,
	io_export_closureOut_56_TVALID,
	io_export_closureOut_57_TREADY,
	io_export_closureOut_57_TVALID,
	io_export_closureOut_58_TREADY,
	io_export_closureOut_58_TVALID,
	io_export_closureOut_59_TREADY,
	io_export_closureOut_59_TVALID,
	io_export_closureOut_60_TREADY,
	io_export_closureOut_60_TVALID,
	io_export_closureOut_61_TREADY,
	io_export_closureOut_61_TVALID,
	io_export_closureOut_62_TREADY,
	io_export_closureOut_62_TVALID,
	io_export_closureOut_63_TREADY,
	io_export_closureOut_63_TVALID,
	io_internal_vcas_axi_full_0_ar_ready,
	io_internal_vcas_axi_full_0_ar_valid,
	io_internal_vcas_axi_full_0_ar_bits_addr,
	io_internal_vcas_axi_full_0_r_ready,
	io_internal_vcas_axi_full_0_r_valid,
	io_internal_vcas_axi_full_0_r_bits_data,
	io_internal_vcas_axi_full_1_ar_ready,
	io_internal_vcas_axi_full_1_ar_valid,
	io_internal_vcas_axi_full_1_ar_bits_addr,
	io_internal_vcas_axi_full_1_r_ready,
	io_internal_vcas_axi_full_1_r_valid,
	io_internal_vcas_axi_full_1_r_bits_data,
	io_internal_vcas_axi_full_2_ar_ready,
	io_internal_vcas_axi_full_2_ar_valid,
	io_internal_vcas_axi_full_2_ar_bits_addr,
	io_internal_vcas_axi_full_2_r_ready,
	io_internal_vcas_axi_full_2_r_valid,
	io_internal_vcas_axi_full_2_r_bits_data,
	io_internal_vcas_axi_full_3_ar_ready,
	io_internal_vcas_axi_full_3_ar_valid,
	io_internal_vcas_axi_full_3_ar_bits_addr,
	io_internal_vcas_axi_full_3_r_ready,
	io_internal_vcas_axi_full_3_r_valid,
	io_internal_vcas_axi_full_3_r_bits_data,
	io_internal_axi_mgmt_vcas_0_ar_ready,
	io_internal_axi_mgmt_vcas_0_ar_valid,
	io_internal_axi_mgmt_vcas_0_ar_bits_addr,
	io_internal_axi_mgmt_vcas_0_ar_bits_prot,
	io_internal_axi_mgmt_vcas_0_r_ready,
	io_internal_axi_mgmt_vcas_0_r_valid,
	io_internal_axi_mgmt_vcas_0_r_bits_data,
	io_internal_axi_mgmt_vcas_0_r_bits_resp,
	io_internal_axi_mgmt_vcas_0_aw_ready,
	io_internal_axi_mgmt_vcas_0_aw_valid,
	io_internal_axi_mgmt_vcas_0_aw_bits_addr,
	io_internal_axi_mgmt_vcas_0_aw_bits_prot,
	io_internal_axi_mgmt_vcas_0_w_ready,
	io_internal_axi_mgmt_vcas_0_w_valid,
	io_internal_axi_mgmt_vcas_0_w_bits_data,
	io_internal_axi_mgmt_vcas_0_w_bits_strb,
	io_internal_axi_mgmt_vcas_0_b_ready,
	io_internal_axi_mgmt_vcas_0_b_valid,
	io_internal_axi_mgmt_vcas_0_b_bits_resp,
	io_internal_axi_mgmt_vcas_1_ar_ready,
	io_internal_axi_mgmt_vcas_1_ar_valid,
	io_internal_axi_mgmt_vcas_1_ar_bits_addr,
	io_internal_axi_mgmt_vcas_1_ar_bits_prot,
	io_internal_axi_mgmt_vcas_1_r_ready,
	io_internal_axi_mgmt_vcas_1_r_valid,
	io_internal_axi_mgmt_vcas_1_r_bits_data,
	io_internal_axi_mgmt_vcas_1_r_bits_resp,
	io_internal_axi_mgmt_vcas_1_aw_ready,
	io_internal_axi_mgmt_vcas_1_aw_valid,
	io_internal_axi_mgmt_vcas_1_aw_bits_addr,
	io_internal_axi_mgmt_vcas_1_aw_bits_prot,
	io_internal_axi_mgmt_vcas_1_w_ready,
	io_internal_axi_mgmt_vcas_1_w_valid,
	io_internal_axi_mgmt_vcas_1_w_bits_data,
	io_internal_axi_mgmt_vcas_1_w_bits_strb,
	io_internal_axi_mgmt_vcas_1_b_ready,
	io_internal_axi_mgmt_vcas_1_b_valid,
	io_internal_axi_mgmt_vcas_1_b_bits_resp,
	io_internal_axi_mgmt_vcas_2_ar_ready,
	io_internal_axi_mgmt_vcas_2_ar_valid,
	io_internal_axi_mgmt_vcas_2_ar_bits_addr,
	io_internal_axi_mgmt_vcas_2_ar_bits_prot,
	io_internal_axi_mgmt_vcas_2_r_ready,
	io_internal_axi_mgmt_vcas_2_r_valid,
	io_internal_axi_mgmt_vcas_2_r_bits_data,
	io_internal_axi_mgmt_vcas_2_r_bits_resp,
	io_internal_axi_mgmt_vcas_2_aw_ready,
	io_internal_axi_mgmt_vcas_2_aw_valid,
	io_internal_axi_mgmt_vcas_2_aw_bits_addr,
	io_internal_axi_mgmt_vcas_2_aw_bits_prot,
	io_internal_axi_mgmt_vcas_2_w_ready,
	io_internal_axi_mgmt_vcas_2_w_valid,
	io_internal_axi_mgmt_vcas_2_w_bits_data,
	io_internal_axi_mgmt_vcas_2_w_bits_strb,
	io_internal_axi_mgmt_vcas_2_b_ready,
	io_internal_axi_mgmt_vcas_2_b_valid,
	io_internal_axi_mgmt_vcas_2_b_bits_resp,
	io_internal_axi_mgmt_vcas_3_ar_ready,
	io_internal_axi_mgmt_vcas_3_ar_valid,
	io_internal_axi_mgmt_vcas_3_ar_bits_addr,
	io_internal_axi_mgmt_vcas_3_ar_bits_prot,
	io_internal_axi_mgmt_vcas_3_r_ready,
	io_internal_axi_mgmt_vcas_3_r_valid,
	io_internal_axi_mgmt_vcas_3_r_bits_data,
	io_internal_axi_mgmt_vcas_3_r_bits_resp,
	io_internal_axi_mgmt_vcas_3_aw_ready,
	io_internal_axi_mgmt_vcas_3_aw_valid,
	io_internal_axi_mgmt_vcas_3_aw_bits_addr,
	io_internal_axi_mgmt_vcas_3_aw_bits_prot,
	io_internal_axi_mgmt_vcas_3_w_ready,
	io_internal_axi_mgmt_vcas_3_w_valid,
	io_internal_axi_mgmt_vcas_3_w_bits_data,
	io_internal_axi_mgmt_vcas_3_w_bits_strb,
	io_internal_axi_mgmt_vcas_3_b_ready,
	io_internal_axi_mgmt_vcas_3_b_valid,
	io_internal_axi_mgmt_vcas_3_b_bits_resp
);
	input clock;
	input reset;
	input io_export_closureOut_0_TREADY;
	output wire io_export_closureOut_0_TVALID;
	input io_export_closureOut_1_TREADY;
	output wire io_export_closureOut_1_TVALID;
	input io_export_closureOut_2_TREADY;
	output wire io_export_closureOut_2_TVALID;
	input io_export_closureOut_3_TREADY;
	output wire io_export_closureOut_3_TVALID;
	input io_export_closureOut_4_TREADY;
	output wire io_export_closureOut_4_TVALID;
	input io_export_closureOut_5_TREADY;
	output wire io_export_closureOut_5_TVALID;
	input io_export_closureOut_6_TREADY;
	output wire io_export_closureOut_6_TVALID;
	input io_export_closureOut_7_TREADY;
	output wire io_export_closureOut_7_TVALID;
	input io_export_closureOut_8_TREADY;
	output wire io_export_closureOut_8_TVALID;
	input io_export_closureOut_9_TREADY;
	output wire io_export_closureOut_9_TVALID;
	input io_export_closureOut_10_TREADY;
	output wire io_export_closureOut_10_TVALID;
	input io_export_closureOut_11_TREADY;
	output wire io_export_closureOut_11_TVALID;
	input io_export_closureOut_12_TREADY;
	output wire io_export_closureOut_12_TVALID;
	input io_export_closureOut_13_TREADY;
	output wire io_export_closureOut_13_TVALID;
	input io_export_closureOut_14_TREADY;
	output wire io_export_closureOut_14_TVALID;
	input io_export_closureOut_15_TREADY;
	output wire io_export_closureOut_15_TVALID;
	input io_export_closureOut_16_TREADY;
	output wire io_export_closureOut_16_TVALID;
	input io_export_closureOut_17_TREADY;
	output wire io_export_closureOut_17_TVALID;
	input io_export_closureOut_18_TREADY;
	output wire io_export_closureOut_18_TVALID;
	input io_export_closureOut_19_TREADY;
	output wire io_export_closureOut_19_TVALID;
	input io_export_closureOut_20_TREADY;
	output wire io_export_closureOut_20_TVALID;
	input io_export_closureOut_21_TREADY;
	output wire io_export_closureOut_21_TVALID;
	input io_export_closureOut_22_TREADY;
	output wire io_export_closureOut_22_TVALID;
	input io_export_closureOut_23_TREADY;
	output wire io_export_closureOut_23_TVALID;
	input io_export_closureOut_24_TREADY;
	output wire io_export_closureOut_24_TVALID;
	input io_export_closureOut_25_TREADY;
	output wire io_export_closureOut_25_TVALID;
	input io_export_closureOut_26_TREADY;
	output wire io_export_closureOut_26_TVALID;
	input io_export_closureOut_27_TREADY;
	output wire io_export_closureOut_27_TVALID;
	input io_export_closureOut_28_TREADY;
	output wire io_export_closureOut_28_TVALID;
	input io_export_closureOut_29_TREADY;
	output wire io_export_closureOut_29_TVALID;
	input io_export_closureOut_30_TREADY;
	output wire io_export_closureOut_30_TVALID;
	input io_export_closureOut_31_TREADY;
	output wire io_export_closureOut_31_TVALID;
	input io_export_closureOut_32_TREADY;
	output wire io_export_closureOut_32_TVALID;
	input io_export_closureOut_33_TREADY;
	output wire io_export_closureOut_33_TVALID;
	input io_export_closureOut_34_TREADY;
	output wire io_export_closureOut_34_TVALID;
	input io_export_closureOut_35_TREADY;
	output wire io_export_closureOut_35_TVALID;
	input io_export_closureOut_36_TREADY;
	output wire io_export_closureOut_36_TVALID;
	input io_export_closureOut_37_TREADY;
	output wire io_export_closureOut_37_TVALID;
	input io_export_closureOut_38_TREADY;
	output wire io_export_closureOut_38_TVALID;
	input io_export_closureOut_39_TREADY;
	output wire io_export_closureOut_39_TVALID;
	input io_export_closureOut_40_TREADY;
	output wire io_export_closureOut_40_TVALID;
	input io_export_closureOut_41_TREADY;
	output wire io_export_closureOut_41_TVALID;
	input io_export_closureOut_42_TREADY;
	output wire io_export_closureOut_42_TVALID;
	input io_export_closureOut_43_TREADY;
	output wire io_export_closureOut_43_TVALID;
	input io_export_closureOut_44_TREADY;
	output wire io_export_closureOut_44_TVALID;
	input io_export_closureOut_45_TREADY;
	output wire io_export_closureOut_45_TVALID;
	input io_export_closureOut_46_TREADY;
	output wire io_export_closureOut_46_TVALID;
	input io_export_closureOut_47_TREADY;
	output wire io_export_closureOut_47_TVALID;
	input io_export_closureOut_48_TREADY;
	output wire io_export_closureOut_48_TVALID;
	input io_export_closureOut_49_TREADY;
	output wire io_export_closureOut_49_TVALID;
	input io_export_closureOut_50_TREADY;
	output wire io_export_closureOut_50_TVALID;
	input io_export_closureOut_51_TREADY;
	output wire io_export_closureOut_51_TVALID;
	input io_export_closureOut_52_TREADY;
	output wire io_export_closureOut_52_TVALID;
	input io_export_closureOut_53_TREADY;
	output wire io_export_closureOut_53_TVALID;
	input io_export_closureOut_54_TREADY;
	output wire io_export_closureOut_54_TVALID;
	input io_export_closureOut_55_TREADY;
	output wire io_export_closureOut_55_TVALID;
	input io_export_closureOut_56_TREADY;
	output wire io_export_closureOut_56_TVALID;
	input io_export_closureOut_57_TREADY;
	output wire io_export_closureOut_57_TVALID;
	input io_export_closureOut_58_TREADY;
	output wire io_export_closureOut_58_TVALID;
	input io_export_closureOut_59_TREADY;
	output wire io_export_closureOut_59_TVALID;
	input io_export_closureOut_60_TREADY;
	output wire io_export_closureOut_60_TVALID;
	input io_export_closureOut_61_TREADY;
	output wire io_export_closureOut_61_TVALID;
	input io_export_closureOut_62_TREADY;
	output wire io_export_closureOut_62_TVALID;
	input io_export_closureOut_63_TREADY;
	output wire io_export_closureOut_63_TVALID;
	input io_internal_vcas_axi_full_0_ar_ready;
	output wire io_internal_vcas_axi_full_0_ar_valid;
	output wire [63:0] io_internal_vcas_axi_full_0_ar_bits_addr;
	output wire io_internal_vcas_axi_full_0_r_ready;
	input io_internal_vcas_axi_full_0_r_valid;
	input [63:0] io_internal_vcas_axi_full_0_r_bits_data;
	input io_internal_vcas_axi_full_1_ar_ready;
	output wire io_internal_vcas_axi_full_1_ar_valid;
	output wire [63:0] io_internal_vcas_axi_full_1_ar_bits_addr;
	output wire io_internal_vcas_axi_full_1_r_ready;
	input io_internal_vcas_axi_full_1_r_valid;
	input [63:0] io_internal_vcas_axi_full_1_r_bits_data;
	input io_internal_vcas_axi_full_2_ar_ready;
	output wire io_internal_vcas_axi_full_2_ar_valid;
	output wire [63:0] io_internal_vcas_axi_full_2_ar_bits_addr;
	output wire io_internal_vcas_axi_full_2_r_ready;
	input io_internal_vcas_axi_full_2_r_valid;
	input [63:0] io_internal_vcas_axi_full_2_r_bits_data;
	input io_internal_vcas_axi_full_3_ar_ready;
	output wire io_internal_vcas_axi_full_3_ar_valid;
	output wire [63:0] io_internal_vcas_axi_full_3_ar_bits_addr;
	output wire io_internal_vcas_axi_full_3_r_ready;
	input io_internal_vcas_axi_full_3_r_valid;
	input [63:0] io_internal_vcas_axi_full_3_r_bits_data;
	output wire io_internal_axi_mgmt_vcas_0_ar_ready;
	input io_internal_axi_mgmt_vcas_0_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_0_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_0_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_0_r_ready;
	output wire io_internal_axi_mgmt_vcas_0_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_0_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_0_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_0_aw_ready;
	input io_internal_axi_mgmt_vcas_0_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_0_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_0_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_0_w_ready;
	input io_internal_axi_mgmt_vcas_0_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_0_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_0_w_bits_strb;
	input io_internal_axi_mgmt_vcas_0_b_ready;
	output wire io_internal_axi_mgmt_vcas_0_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_0_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_1_ar_ready;
	input io_internal_axi_mgmt_vcas_1_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_1_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_1_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_1_r_ready;
	output wire io_internal_axi_mgmt_vcas_1_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_1_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_1_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_1_aw_ready;
	input io_internal_axi_mgmt_vcas_1_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_1_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_1_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_1_w_ready;
	input io_internal_axi_mgmt_vcas_1_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_1_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_1_w_bits_strb;
	input io_internal_axi_mgmt_vcas_1_b_ready;
	output wire io_internal_axi_mgmt_vcas_1_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_1_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_2_ar_ready;
	input io_internal_axi_mgmt_vcas_2_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_2_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_2_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_2_r_ready;
	output wire io_internal_axi_mgmt_vcas_2_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_2_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_2_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_2_aw_ready;
	input io_internal_axi_mgmt_vcas_2_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_2_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_2_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_2_w_ready;
	input io_internal_axi_mgmt_vcas_2_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_2_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_2_w_bits_strb;
	input io_internal_axi_mgmt_vcas_2_b_ready;
	output wire io_internal_axi_mgmt_vcas_2_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_2_b_bits_resp;
	output wire io_internal_axi_mgmt_vcas_3_ar_ready;
	input io_internal_axi_mgmt_vcas_3_ar_valid;
	input [5:0] io_internal_axi_mgmt_vcas_3_ar_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_3_ar_bits_prot;
	input io_internal_axi_mgmt_vcas_3_r_ready;
	output wire io_internal_axi_mgmt_vcas_3_r_valid;
	output wire [63:0] io_internal_axi_mgmt_vcas_3_r_bits_data;
	output wire [1:0] io_internal_axi_mgmt_vcas_3_r_bits_resp;
	output wire io_internal_axi_mgmt_vcas_3_aw_ready;
	input io_internal_axi_mgmt_vcas_3_aw_valid;
	input [5:0] io_internal_axi_mgmt_vcas_3_aw_bits_addr;
	input [2:0] io_internal_axi_mgmt_vcas_3_aw_bits_prot;
	output wire io_internal_axi_mgmt_vcas_3_w_ready;
	input io_internal_axi_mgmt_vcas_3_w_valid;
	input [63:0] io_internal_axi_mgmt_vcas_3_w_bits_data;
	input [7:0] io_internal_axi_mgmt_vcas_3_w_bits_strb;
	input io_internal_axi_mgmt_vcas_3_b_ready;
	output wire io_internal_axi_mgmt_vcas_3_b_valid;
	output wire [1:0] io_internal_axi_mgmt_vcas_3_b_bits_resp;
	wire _axis_stream_converters_out_63_io_dataIn_TREADY;
	wire _axis_stream_converters_out_62_io_dataIn_TREADY;
	wire _axis_stream_converters_out_61_io_dataIn_TREADY;
	wire _axis_stream_converters_out_60_io_dataIn_TREADY;
	wire _axis_stream_converters_out_59_io_dataIn_TREADY;
	wire _axis_stream_converters_out_58_io_dataIn_TREADY;
	wire _axis_stream_converters_out_57_io_dataIn_TREADY;
	wire _axis_stream_converters_out_56_io_dataIn_TREADY;
	wire _axis_stream_converters_out_55_io_dataIn_TREADY;
	wire _axis_stream_converters_out_54_io_dataIn_TREADY;
	wire _axis_stream_converters_out_53_io_dataIn_TREADY;
	wire _axis_stream_converters_out_52_io_dataIn_TREADY;
	wire _axis_stream_converters_out_51_io_dataIn_TREADY;
	wire _axis_stream_converters_out_50_io_dataIn_TREADY;
	wire _axis_stream_converters_out_49_io_dataIn_TREADY;
	wire _axis_stream_converters_out_48_io_dataIn_TREADY;
	wire _axis_stream_converters_out_47_io_dataIn_TREADY;
	wire _axis_stream_converters_out_46_io_dataIn_TREADY;
	wire _axis_stream_converters_out_45_io_dataIn_TREADY;
	wire _axis_stream_converters_out_44_io_dataIn_TREADY;
	wire _axis_stream_converters_out_43_io_dataIn_TREADY;
	wire _axis_stream_converters_out_42_io_dataIn_TREADY;
	wire _axis_stream_converters_out_41_io_dataIn_TREADY;
	wire _axis_stream_converters_out_40_io_dataIn_TREADY;
	wire _axis_stream_converters_out_39_io_dataIn_TREADY;
	wire _axis_stream_converters_out_38_io_dataIn_TREADY;
	wire _axis_stream_converters_out_37_io_dataIn_TREADY;
	wire _axis_stream_converters_out_36_io_dataIn_TREADY;
	wire _axis_stream_converters_out_35_io_dataIn_TREADY;
	wire _axis_stream_converters_out_34_io_dataIn_TREADY;
	wire _axis_stream_converters_out_33_io_dataIn_TREADY;
	wire _axis_stream_converters_out_32_io_dataIn_TREADY;
	wire _axis_stream_converters_out_31_io_dataIn_TREADY;
	wire _axis_stream_converters_out_30_io_dataIn_TREADY;
	wire _axis_stream_converters_out_29_io_dataIn_TREADY;
	wire _axis_stream_converters_out_28_io_dataIn_TREADY;
	wire _axis_stream_converters_out_27_io_dataIn_TREADY;
	wire _axis_stream_converters_out_26_io_dataIn_TREADY;
	wire _axis_stream_converters_out_25_io_dataIn_TREADY;
	wire _axis_stream_converters_out_24_io_dataIn_TREADY;
	wire _axis_stream_converters_out_23_io_dataIn_TREADY;
	wire _axis_stream_converters_out_22_io_dataIn_TREADY;
	wire _axis_stream_converters_out_21_io_dataIn_TREADY;
	wire _axis_stream_converters_out_20_io_dataIn_TREADY;
	wire _axis_stream_converters_out_19_io_dataIn_TREADY;
	wire _axis_stream_converters_out_18_io_dataIn_TREADY;
	wire _axis_stream_converters_out_17_io_dataIn_TREADY;
	wire _axis_stream_converters_out_16_io_dataIn_TREADY;
	wire _axis_stream_converters_out_15_io_dataIn_TREADY;
	wire _axis_stream_converters_out_14_io_dataIn_TREADY;
	wire _axis_stream_converters_out_13_io_dataIn_TREADY;
	wire _axis_stream_converters_out_12_io_dataIn_TREADY;
	wire _axis_stream_converters_out_11_io_dataIn_TREADY;
	wire _axis_stream_converters_out_10_io_dataIn_TREADY;
	wire _axis_stream_converters_out_9_io_dataIn_TREADY;
	wire _axis_stream_converters_out_8_io_dataIn_TREADY;
	wire _axis_stream_converters_out_7_io_dataIn_TREADY;
	wire _axis_stream_converters_out_6_io_dataIn_TREADY;
	wire _axis_stream_converters_out_5_io_dataIn_TREADY;
	wire _axis_stream_converters_out_4_io_dataIn_TREADY;
	wire _axis_stream_converters_out_3_io_dataIn_TREADY;
	wire _axis_stream_converters_out_2_io_dataIn_TREADY;
	wire _axis_stream_converters_out_1_io_dataIn_TREADY;
	wire _axis_stream_converters_out_0_io_dataIn_TREADY;
	wire _vcasRvmRO_3_io_read_address_ready;
	wire _vcasRvmRO_3_io_read_data_valid;
	wire [63:0] _vcasRvmRO_3_io_read_data_bits;
	wire _vcasRvmRO_2_io_read_address_ready;
	wire _vcasRvmRO_2_io_read_data_valid;
	wire [63:0] _vcasRvmRO_2_io_read_data_bits;
	wire _vcasRvmRO_1_io_read_address_ready;
	wire _vcasRvmRO_1_io_read_data_valid;
	wire [63:0] _vcasRvmRO_1_io_read_data_bits;
	wire _vcasRvmRO_0_io_read_address_ready;
	wire _vcasRvmRO_0_io_read_data_valid;
	wire [63:0] _vcasRvmRO_0_io_read_data_bits;
	wire _vcas_3_io_dataOut_valid;
	wire [63:0] _vcas_3_io_dataOut_bits;
	wire _vcas_3_io_read_address_valid;
	wire [63:0] _vcas_3_io_read_address_bits;
	wire _vcas_3_io_read_data_ready;
	wire _vcas_2_io_dataOut_valid;
	wire [63:0] _vcas_2_io_dataOut_bits;
	wire _vcas_2_io_read_address_valid;
	wire [63:0] _vcas_2_io_read_address_bits;
	wire _vcas_2_io_read_data_ready;
	wire _vcas_1_io_dataOut_valid;
	wire [63:0] _vcas_1_io_dataOut_bits;
	wire _vcas_1_io_read_address_valid;
	wire [63:0] _vcas_1_io_read_address_bits;
	wire _vcas_1_io_read_data_ready;
	wire _vcas_0_io_dataOut_valid;
	wire [63:0] _vcas_0_io_dataOut_bits;
	wire _vcas_0_io_read_address_valid;
	wire [63:0] _vcas_0_io_read_address_bits;
	wire _vcas_0_io_read_data_ready;
	wire _continuationNetwork_io_connVCAS_0_ready;
	wire _continuationNetwork_io_connVCAS_1_ready;
	wire _continuationNetwork_io_connVCAS_2_ready;
	wire _continuationNetwork_io_connVCAS_3_ready;
	wire _continuationNetwork_io_connPE_0_valid;
	wire _continuationNetwork_io_connPE_1_valid;
	wire _continuationNetwork_io_connPE_2_valid;
	wire _continuationNetwork_io_connPE_3_valid;
	wire _continuationNetwork_io_connPE_4_valid;
	wire _continuationNetwork_io_connPE_5_valid;
	wire _continuationNetwork_io_connPE_6_valid;
	wire _continuationNetwork_io_connPE_7_valid;
	wire _continuationNetwork_io_connPE_8_valid;
	wire _continuationNetwork_io_connPE_9_valid;
	wire _continuationNetwork_io_connPE_10_valid;
	wire _continuationNetwork_io_connPE_11_valid;
	wire _continuationNetwork_io_connPE_12_valid;
	wire _continuationNetwork_io_connPE_13_valid;
	wire _continuationNetwork_io_connPE_14_valid;
	wire _continuationNetwork_io_connPE_15_valid;
	wire _continuationNetwork_io_connPE_16_valid;
	wire _continuationNetwork_io_connPE_17_valid;
	wire _continuationNetwork_io_connPE_18_valid;
	wire _continuationNetwork_io_connPE_19_valid;
	wire _continuationNetwork_io_connPE_20_valid;
	wire _continuationNetwork_io_connPE_21_valid;
	wire _continuationNetwork_io_connPE_22_valid;
	wire _continuationNetwork_io_connPE_23_valid;
	wire _continuationNetwork_io_connPE_24_valid;
	wire _continuationNetwork_io_connPE_25_valid;
	wire _continuationNetwork_io_connPE_26_valid;
	wire _continuationNetwork_io_connPE_27_valid;
	wire _continuationNetwork_io_connPE_28_valid;
	wire _continuationNetwork_io_connPE_29_valid;
	wire _continuationNetwork_io_connPE_30_valid;
	wire _continuationNetwork_io_connPE_31_valid;
	wire _continuationNetwork_io_connPE_32_valid;
	wire _continuationNetwork_io_connPE_33_valid;
	wire _continuationNetwork_io_connPE_34_valid;
	wire _continuationNetwork_io_connPE_35_valid;
	wire _continuationNetwork_io_connPE_36_valid;
	wire _continuationNetwork_io_connPE_37_valid;
	wire _continuationNetwork_io_connPE_38_valid;
	wire _continuationNetwork_io_connPE_39_valid;
	wire _continuationNetwork_io_connPE_40_valid;
	wire _continuationNetwork_io_connPE_41_valid;
	wire _continuationNetwork_io_connPE_42_valid;
	wire _continuationNetwork_io_connPE_43_valid;
	wire _continuationNetwork_io_connPE_44_valid;
	wire _continuationNetwork_io_connPE_45_valid;
	wire _continuationNetwork_io_connPE_46_valid;
	wire _continuationNetwork_io_connPE_47_valid;
	wire _continuationNetwork_io_connPE_48_valid;
	wire _continuationNetwork_io_connPE_49_valid;
	wire _continuationNetwork_io_connPE_50_valid;
	wire _continuationNetwork_io_connPE_51_valid;
	wire _continuationNetwork_io_connPE_52_valid;
	wire _continuationNetwork_io_connPE_53_valid;
	wire _continuationNetwork_io_connPE_54_valid;
	wire _continuationNetwork_io_connPE_55_valid;
	wire _continuationNetwork_io_connPE_56_valid;
	wire _continuationNetwork_io_connPE_57_valid;
	wire _continuationNetwork_io_connPE_58_valid;
	wire _continuationNetwork_io_connPE_59_valid;
	wire _continuationNetwork_io_connPE_60_valid;
	wire _continuationNetwork_io_connPE_61_valid;
	wire _continuationNetwork_io_connPE_62_valid;
	wire _continuationNetwork_io_connPE_63_valid;
	AllocatorNetwork continuationNetwork(
		.clock(clock),
		.reset(reset),
		.io_connVCAS_0_ready(_continuationNetwork_io_connVCAS_0_ready),
		.io_connVCAS_0_valid(_vcas_0_io_dataOut_valid),
		.io_connVCAS_0_bits(_vcas_0_io_dataOut_bits),
		.io_connVCAS_1_ready(_continuationNetwork_io_connVCAS_1_ready),
		.io_connVCAS_1_valid(_vcas_1_io_dataOut_valid),
		.io_connVCAS_1_bits(_vcas_1_io_dataOut_bits),
		.io_connVCAS_2_ready(_continuationNetwork_io_connVCAS_2_ready),
		.io_connVCAS_2_valid(_vcas_2_io_dataOut_valid),
		.io_connVCAS_2_bits(_vcas_2_io_dataOut_bits),
		.io_connVCAS_3_ready(_continuationNetwork_io_connVCAS_3_ready),
		.io_connVCAS_3_valid(_vcas_3_io_dataOut_valid),
		.io_connVCAS_3_bits(_vcas_3_io_dataOut_bits),
		.io_connPE_0_ready(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_connPE_0_valid(_continuationNetwork_io_connPE_0_valid),
		.io_connPE_1_ready(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_connPE_1_valid(_continuationNetwork_io_connPE_1_valid),
		.io_connPE_2_ready(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_connPE_2_valid(_continuationNetwork_io_connPE_2_valid),
		.io_connPE_3_ready(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_connPE_3_valid(_continuationNetwork_io_connPE_3_valid),
		.io_connPE_4_ready(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_connPE_4_valid(_continuationNetwork_io_connPE_4_valid),
		.io_connPE_5_ready(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_connPE_5_valid(_continuationNetwork_io_connPE_5_valid),
		.io_connPE_6_ready(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_connPE_6_valid(_continuationNetwork_io_connPE_6_valid),
		.io_connPE_7_ready(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_connPE_7_valid(_continuationNetwork_io_connPE_7_valid),
		.io_connPE_8_ready(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_connPE_8_valid(_continuationNetwork_io_connPE_8_valid),
		.io_connPE_9_ready(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_connPE_9_valid(_continuationNetwork_io_connPE_9_valid),
		.io_connPE_10_ready(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_connPE_10_valid(_continuationNetwork_io_connPE_10_valid),
		.io_connPE_11_ready(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_connPE_11_valid(_continuationNetwork_io_connPE_11_valid),
		.io_connPE_12_ready(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_connPE_12_valid(_continuationNetwork_io_connPE_12_valid),
		.io_connPE_13_ready(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_connPE_13_valid(_continuationNetwork_io_connPE_13_valid),
		.io_connPE_14_ready(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_connPE_14_valid(_continuationNetwork_io_connPE_14_valid),
		.io_connPE_15_ready(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_connPE_15_valid(_continuationNetwork_io_connPE_15_valid),
		.io_connPE_16_ready(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_connPE_16_valid(_continuationNetwork_io_connPE_16_valid),
		.io_connPE_17_ready(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_connPE_17_valid(_continuationNetwork_io_connPE_17_valid),
		.io_connPE_18_ready(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_connPE_18_valid(_continuationNetwork_io_connPE_18_valid),
		.io_connPE_19_ready(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_connPE_19_valid(_continuationNetwork_io_connPE_19_valid),
		.io_connPE_20_ready(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_connPE_20_valid(_continuationNetwork_io_connPE_20_valid),
		.io_connPE_21_ready(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_connPE_21_valid(_continuationNetwork_io_connPE_21_valid),
		.io_connPE_22_ready(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_connPE_22_valid(_continuationNetwork_io_connPE_22_valid),
		.io_connPE_23_ready(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_connPE_23_valid(_continuationNetwork_io_connPE_23_valid),
		.io_connPE_24_ready(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_connPE_24_valid(_continuationNetwork_io_connPE_24_valid),
		.io_connPE_25_ready(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_connPE_25_valid(_continuationNetwork_io_connPE_25_valid),
		.io_connPE_26_ready(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_connPE_26_valid(_continuationNetwork_io_connPE_26_valid),
		.io_connPE_27_ready(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_connPE_27_valid(_continuationNetwork_io_connPE_27_valid),
		.io_connPE_28_ready(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_connPE_28_valid(_continuationNetwork_io_connPE_28_valid),
		.io_connPE_29_ready(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_connPE_29_valid(_continuationNetwork_io_connPE_29_valid),
		.io_connPE_30_ready(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_connPE_30_valid(_continuationNetwork_io_connPE_30_valid),
		.io_connPE_31_ready(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_connPE_31_valid(_continuationNetwork_io_connPE_31_valid),
		.io_connPE_32_ready(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_connPE_32_valid(_continuationNetwork_io_connPE_32_valid),
		.io_connPE_33_ready(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_connPE_33_valid(_continuationNetwork_io_connPE_33_valid),
		.io_connPE_34_ready(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_connPE_34_valid(_continuationNetwork_io_connPE_34_valid),
		.io_connPE_35_ready(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_connPE_35_valid(_continuationNetwork_io_connPE_35_valid),
		.io_connPE_36_ready(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_connPE_36_valid(_continuationNetwork_io_connPE_36_valid),
		.io_connPE_37_ready(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_connPE_37_valid(_continuationNetwork_io_connPE_37_valid),
		.io_connPE_38_ready(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_connPE_38_valid(_continuationNetwork_io_connPE_38_valid),
		.io_connPE_39_ready(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_connPE_39_valid(_continuationNetwork_io_connPE_39_valid),
		.io_connPE_40_ready(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_connPE_40_valid(_continuationNetwork_io_connPE_40_valid),
		.io_connPE_41_ready(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_connPE_41_valid(_continuationNetwork_io_connPE_41_valid),
		.io_connPE_42_ready(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_connPE_42_valid(_continuationNetwork_io_connPE_42_valid),
		.io_connPE_43_ready(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_connPE_43_valid(_continuationNetwork_io_connPE_43_valid),
		.io_connPE_44_ready(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_connPE_44_valid(_continuationNetwork_io_connPE_44_valid),
		.io_connPE_45_ready(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_connPE_45_valid(_continuationNetwork_io_connPE_45_valid),
		.io_connPE_46_ready(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_connPE_46_valid(_continuationNetwork_io_connPE_46_valid),
		.io_connPE_47_ready(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_connPE_47_valid(_continuationNetwork_io_connPE_47_valid),
		.io_connPE_48_ready(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_connPE_48_valid(_continuationNetwork_io_connPE_48_valid),
		.io_connPE_49_ready(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_connPE_49_valid(_continuationNetwork_io_connPE_49_valid),
		.io_connPE_50_ready(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_connPE_50_valid(_continuationNetwork_io_connPE_50_valid),
		.io_connPE_51_ready(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_connPE_51_valid(_continuationNetwork_io_connPE_51_valid),
		.io_connPE_52_ready(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_connPE_52_valid(_continuationNetwork_io_connPE_52_valid),
		.io_connPE_53_ready(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_connPE_53_valid(_continuationNetwork_io_connPE_53_valid),
		.io_connPE_54_ready(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_connPE_54_valid(_continuationNetwork_io_connPE_54_valid),
		.io_connPE_55_ready(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_connPE_55_valid(_continuationNetwork_io_connPE_55_valid),
		.io_connPE_56_ready(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_connPE_56_valid(_continuationNetwork_io_connPE_56_valid),
		.io_connPE_57_ready(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_connPE_57_valid(_continuationNetwork_io_connPE_57_valid),
		.io_connPE_58_ready(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_connPE_58_valid(_continuationNetwork_io_connPE_58_valid),
		.io_connPE_59_ready(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_connPE_59_valid(_continuationNetwork_io_connPE_59_valid),
		.io_connPE_60_ready(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_connPE_60_valid(_continuationNetwork_io_connPE_60_valid),
		.io_connPE_61_ready(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_connPE_61_valid(_continuationNetwork_io_connPE_61_valid),
		.io_connPE_62_ready(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_connPE_62_valid(_continuationNetwork_io_connPE_62_valid),
		.io_connPE_63_ready(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_connPE_63_valid(_continuationNetwork_io_connPE_63_valid)
	);
	AllocatorServer vcas_0(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_0_ready),
		.io_dataOut_valid(_vcas_0_io_dataOut_valid),
		.io_dataOut_bits(_vcas_0_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_0_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_0_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_0_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_0_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_0_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_0_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_0_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_0_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_0_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_0_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_0_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_0_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_0_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_0_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_0_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_0_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_0_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_0_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_0_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_0_io_read_address_ready),
		.io_read_address_valid(_vcas_0_io_read_address_valid),
		.io_read_address_bits(_vcas_0_io_read_address_bits),
		.io_read_data_ready(_vcas_0_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_0_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_0_io_read_data_bits)
	);
	AllocatorServer vcas_1(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_1_ready),
		.io_dataOut_valid(_vcas_1_io_dataOut_valid),
		.io_dataOut_bits(_vcas_1_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_1_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_1_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_1_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_1_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_1_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_1_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_1_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_1_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_1_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_1_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_1_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_1_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_1_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_1_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_1_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_1_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_1_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_1_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_1_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_1_io_read_address_ready),
		.io_read_address_valid(_vcas_1_io_read_address_valid),
		.io_read_address_bits(_vcas_1_io_read_address_bits),
		.io_read_data_ready(_vcas_1_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_1_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_1_io_read_data_bits)
	);
	AllocatorServer vcas_2(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_2_ready),
		.io_dataOut_valid(_vcas_2_io_dataOut_valid),
		.io_dataOut_bits(_vcas_2_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_2_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_2_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_2_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_2_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_2_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_2_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_2_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_2_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_2_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_2_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_2_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_2_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_2_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_2_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_2_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_2_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_2_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_2_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_2_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_2_io_read_address_ready),
		.io_read_address_valid(_vcas_2_io_read_address_valid),
		.io_read_address_bits(_vcas_2_io_read_address_bits),
		.io_read_data_ready(_vcas_2_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_2_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_2_io_read_data_bits)
	);
	AllocatorServer vcas_3(
		.clock(clock),
		.reset(reset),
		.io_dataOut_ready(_continuationNetwork_io_connVCAS_3_ready),
		.io_dataOut_valid(_vcas_3_io_dataOut_valid),
		.io_dataOut_bits(_vcas_3_io_dataOut_bits),
		.io_axi_mgmt_ar_ready(io_internal_axi_mgmt_vcas_3_ar_ready),
		.io_axi_mgmt_ar_valid(io_internal_axi_mgmt_vcas_3_ar_valid),
		.io_axi_mgmt_ar_bits_addr(io_internal_axi_mgmt_vcas_3_ar_bits_addr),
		.io_axi_mgmt_ar_bits_prot(io_internal_axi_mgmt_vcas_3_ar_bits_prot),
		.io_axi_mgmt_r_ready(io_internal_axi_mgmt_vcas_3_r_ready),
		.io_axi_mgmt_r_valid(io_internal_axi_mgmt_vcas_3_r_valid),
		.io_axi_mgmt_r_bits_data(io_internal_axi_mgmt_vcas_3_r_bits_data),
		.io_axi_mgmt_r_bits_resp(io_internal_axi_mgmt_vcas_3_r_bits_resp),
		.io_axi_mgmt_aw_ready(io_internal_axi_mgmt_vcas_3_aw_ready),
		.io_axi_mgmt_aw_valid(io_internal_axi_mgmt_vcas_3_aw_valid),
		.io_axi_mgmt_aw_bits_addr(io_internal_axi_mgmt_vcas_3_aw_bits_addr),
		.io_axi_mgmt_aw_bits_prot(io_internal_axi_mgmt_vcas_3_aw_bits_prot),
		.io_axi_mgmt_w_ready(io_internal_axi_mgmt_vcas_3_w_ready),
		.io_axi_mgmt_w_valid(io_internal_axi_mgmt_vcas_3_w_valid),
		.io_axi_mgmt_w_bits_data(io_internal_axi_mgmt_vcas_3_w_bits_data),
		.io_axi_mgmt_w_bits_strb(io_internal_axi_mgmt_vcas_3_w_bits_strb),
		.io_axi_mgmt_b_ready(io_internal_axi_mgmt_vcas_3_b_ready),
		.io_axi_mgmt_b_valid(io_internal_axi_mgmt_vcas_3_b_valid),
		.io_axi_mgmt_b_bits_resp(io_internal_axi_mgmt_vcas_3_b_bits_resp),
		.io_read_address_ready(_vcasRvmRO_3_io_read_address_ready),
		.io_read_address_valid(_vcas_3_io_read_address_valid),
		.io_read_address_bits(_vcas_3_io_read_address_bits),
		.io_read_data_ready(_vcas_3_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_3_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_3_io_read_data_bits)
	);
	RVtoAXIBridge_2 vcasRvmRO_0(
		.io_read_address_ready(_vcasRvmRO_0_io_read_address_ready),
		.io_read_address_valid(_vcas_0_io_read_address_valid),
		.io_read_address_bits(_vcas_0_io_read_address_bits),
		.io_read_data_ready(_vcas_0_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_0_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_0_io_read_data_bits),
		.axi_ar_ready(io_internal_vcas_axi_full_0_ar_ready),
		.axi_ar_valid(io_internal_vcas_axi_full_0_ar_valid),
		.axi_ar_bits_addr(io_internal_vcas_axi_full_0_ar_bits_addr),
		.axi_r_ready(io_internal_vcas_axi_full_0_r_ready),
		.axi_r_valid(io_internal_vcas_axi_full_0_r_valid),
		.axi_r_bits_data(io_internal_vcas_axi_full_0_r_bits_data)
	);
	RVtoAXIBridge_2 vcasRvmRO_1(
		.io_read_address_ready(_vcasRvmRO_1_io_read_address_ready),
		.io_read_address_valid(_vcas_1_io_read_address_valid),
		.io_read_address_bits(_vcas_1_io_read_address_bits),
		.io_read_data_ready(_vcas_1_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_1_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_1_io_read_data_bits),
		.axi_ar_ready(io_internal_vcas_axi_full_1_ar_ready),
		.axi_ar_valid(io_internal_vcas_axi_full_1_ar_valid),
		.axi_ar_bits_addr(io_internal_vcas_axi_full_1_ar_bits_addr),
		.axi_r_ready(io_internal_vcas_axi_full_1_r_ready),
		.axi_r_valid(io_internal_vcas_axi_full_1_r_valid),
		.axi_r_bits_data(io_internal_vcas_axi_full_1_r_bits_data)
	);
	RVtoAXIBridge_2 vcasRvmRO_2(
		.io_read_address_ready(_vcasRvmRO_2_io_read_address_ready),
		.io_read_address_valid(_vcas_2_io_read_address_valid),
		.io_read_address_bits(_vcas_2_io_read_address_bits),
		.io_read_data_ready(_vcas_2_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_2_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_2_io_read_data_bits),
		.axi_ar_ready(io_internal_vcas_axi_full_2_ar_ready),
		.axi_ar_valid(io_internal_vcas_axi_full_2_ar_valid),
		.axi_ar_bits_addr(io_internal_vcas_axi_full_2_ar_bits_addr),
		.axi_r_ready(io_internal_vcas_axi_full_2_r_ready),
		.axi_r_valid(io_internal_vcas_axi_full_2_r_valid),
		.axi_r_bits_data(io_internal_vcas_axi_full_2_r_bits_data)
	);
	RVtoAXIBridge_2 vcasRvmRO_3(
		.io_read_address_ready(_vcasRvmRO_3_io_read_address_ready),
		.io_read_address_valid(_vcas_3_io_read_address_valid),
		.io_read_address_bits(_vcas_3_io_read_address_bits),
		.io_read_data_ready(_vcas_3_io_read_data_ready),
		.io_read_data_valid(_vcasRvmRO_3_io_read_data_valid),
		.io_read_data_bits(_vcasRvmRO_3_io_read_data_bits),
		.axi_ar_ready(io_internal_vcas_axi_full_3_ar_ready),
		.axi_ar_valid(io_internal_vcas_axi_full_3_ar_valid),
		.axi_ar_bits_addr(io_internal_vcas_axi_full_3_ar_bits_addr),
		.axi_r_ready(io_internal_vcas_axi_full_3_r_ready),
		.axi_r_valid(io_internal_vcas_axi_full_3_r_valid),
		.axi_r_bits_data(io_internal_vcas_axi_full_3_r_bits_data)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_0(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_0_valid),
		.io_dataOut_TREADY(io_export_closureOut_0_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_0_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_1(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_1_valid),
		.io_dataOut_TREADY(io_export_closureOut_1_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_1_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_2(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_2_valid),
		.io_dataOut_TREADY(io_export_closureOut_2_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_2_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_3(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_3_valid),
		.io_dataOut_TREADY(io_export_closureOut_3_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_3_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_4(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_4_valid),
		.io_dataOut_TREADY(io_export_closureOut_4_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_4_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_5(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_5_valid),
		.io_dataOut_TREADY(io_export_closureOut_5_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_5_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_6(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_6_valid),
		.io_dataOut_TREADY(io_export_closureOut_6_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_6_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_7(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_7_valid),
		.io_dataOut_TREADY(io_export_closureOut_7_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_7_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_8(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_8_valid),
		.io_dataOut_TREADY(io_export_closureOut_8_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_8_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_9(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_9_valid),
		.io_dataOut_TREADY(io_export_closureOut_9_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_9_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_10(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_10_valid),
		.io_dataOut_TREADY(io_export_closureOut_10_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_10_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_11(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_11_valid),
		.io_dataOut_TREADY(io_export_closureOut_11_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_11_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_12(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_12_valid),
		.io_dataOut_TREADY(io_export_closureOut_12_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_12_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_13(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_13_valid),
		.io_dataOut_TREADY(io_export_closureOut_13_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_13_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_14(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_14_valid),
		.io_dataOut_TREADY(io_export_closureOut_14_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_14_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_15(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_15_valid),
		.io_dataOut_TREADY(io_export_closureOut_15_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_15_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_16(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_16_valid),
		.io_dataOut_TREADY(io_export_closureOut_16_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_16_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_17(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_17_valid),
		.io_dataOut_TREADY(io_export_closureOut_17_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_17_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_18(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_18_valid),
		.io_dataOut_TREADY(io_export_closureOut_18_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_18_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_19(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_19_valid),
		.io_dataOut_TREADY(io_export_closureOut_19_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_19_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_20(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_20_valid),
		.io_dataOut_TREADY(io_export_closureOut_20_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_20_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_21(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_21_valid),
		.io_dataOut_TREADY(io_export_closureOut_21_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_21_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_22(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_22_valid),
		.io_dataOut_TREADY(io_export_closureOut_22_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_22_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_23(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_23_valid),
		.io_dataOut_TREADY(io_export_closureOut_23_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_23_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_24(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_24_valid),
		.io_dataOut_TREADY(io_export_closureOut_24_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_24_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_25(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_25_valid),
		.io_dataOut_TREADY(io_export_closureOut_25_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_25_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_26(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_26_valid),
		.io_dataOut_TREADY(io_export_closureOut_26_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_26_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_27(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_27_valid),
		.io_dataOut_TREADY(io_export_closureOut_27_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_27_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_28(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_28_valid),
		.io_dataOut_TREADY(io_export_closureOut_28_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_28_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_29(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_29_valid),
		.io_dataOut_TREADY(io_export_closureOut_29_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_29_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_30(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_30_valid),
		.io_dataOut_TREADY(io_export_closureOut_30_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_30_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_31(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_31_valid),
		.io_dataOut_TREADY(io_export_closureOut_31_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_31_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_32(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_32_valid),
		.io_dataOut_TREADY(io_export_closureOut_32_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_32_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_33(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_33_valid),
		.io_dataOut_TREADY(io_export_closureOut_33_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_33_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_34(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_34_valid),
		.io_dataOut_TREADY(io_export_closureOut_34_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_34_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_35(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_35_valid),
		.io_dataOut_TREADY(io_export_closureOut_35_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_35_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_36(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_36_valid),
		.io_dataOut_TREADY(io_export_closureOut_36_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_36_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_37(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_37_valid),
		.io_dataOut_TREADY(io_export_closureOut_37_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_37_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_38(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_38_valid),
		.io_dataOut_TREADY(io_export_closureOut_38_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_38_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_39(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_39_valid),
		.io_dataOut_TREADY(io_export_closureOut_39_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_39_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_40(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_40_valid),
		.io_dataOut_TREADY(io_export_closureOut_40_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_40_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_41(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_41_valid),
		.io_dataOut_TREADY(io_export_closureOut_41_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_41_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_42(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_42_valid),
		.io_dataOut_TREADY(io_export_closureOut_42_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_42_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_43(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_43_valid),
		.io_dataOut_TREADY(io_export_closureOut_43_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_43_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_44(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_44_valid),
		.io_dataOut_TREADY(io_export_closureOut_44_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_44_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_45(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_45_valid),
		.io_dataOut_TREADY(io_export_closureOut_45_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_45_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_46(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_46_valid),
		.io_dataOut_TREADY(io_export_closureOut_46_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_46_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_47(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_47_valid),
		.io_dataOut_TREADY(io_export_closureOut_47_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_47_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_48(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_48_valid),
		.io_dataOut_TREADY(io_export_closureOut_48_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_48_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_49(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_49_valid),
		.io_dataOut_TREADY(io_export_closureOut_49_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_49_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_50(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_50_valid),
		.io_dataOut_TREADY(io_export_closureOut_50_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_50_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_51(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_51_valid),
		.io_dataOut_TREADY(io_export_closureOut_51_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_51_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_52(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_52_valid),
		.io_dataOut_TREADY(io_export_closureOut_52_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_52_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_53(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_53_valid),
		.io_dataOut_TREADY(io_export_closureOut_53_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_53_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_54(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_54_valid),
		.io_dataOut_TREADY(io_export_closureOut_54_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_54_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_55(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_55_valid),
		.io_dataOut_TREADY(io_export_closureOut_55_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_55_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_56(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_56_valid),
		.io_dataOut_TREADY(io_export_closureOut_56_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_56_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_57(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_57_valid),
		.io_dataOut_TREADY(io_export_closureOut_57_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_57_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_58(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_58_valid),
		.io_dataOut_TREADY(io_export_closureOut_58_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_58_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_59(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_59_valid),
		.io_dataOut_TREADY(io_export_closureOut_59_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_59_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_60(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_60_valid),
		.io_dataOut_TREADY(io_export_closureOut_60_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_60_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_61(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_61_valid),
		.io_dataOut_TREADY(io_export_closureOut_61_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_61_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_62(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_62_valid),
		.io_dataOut_TREADY(io_export_closureOut_62_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_62_TVALID)
	);
	AxisDataWidthConverter_144 axis_stream_converters_out_63(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_out_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(_continuationNetwork_io_connPE_63_valid),
		.io_dataOut_TREADY(io_export_closureOut_63_TREADY),
		.io_dataOut_TVALID(io_export_closureOut_63_TVALID)
	);
endmodule
module ArgumentNotifierNetworkUnit (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_peAddress_ready,
	io_peAddress_valid,
	io_peAddress_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	output wire io_peAddress_ready;
	input io_peAddress_valid;
	input [63:0] io_peAddress_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg stateReg;
	reg [63:0] addressReg;
	reg priorityReg;
	wire _GEN = io_addressIn_valid & io_peAddress_valid;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 1'h0;
			addressReg <= 64'h0000000000000000;
			priorityReg <= 1'h1;
		end
		else begin
			if (stateReg)
				stateReg <= stateReg & ~io_addressOut_ready;
			else begin
				stateReg <= (io_addressIn_valid | io_peAddress_valid) | stateReg;
				if (_GEN)
					addressReg <= (priorityReg ? io_peAddress_bits : io_addressIn_bits);
				else if (io_peAddress_valid)
					addressReg <= io_peAddress_bits;
				else if (io_addressIn_valid)
					addressReg <= io_addressIn_bits;
			end
			priorityReg <= (~stateReg & _GEN) ^ priorityReg;
		end
	assign io_addressIn_ready = ~stateReg & (_GEN ? ~priorityReg : ~io_peAddress_valid & io_addressIn_valid);
	assign io_peAddress_ready = ~stateReg & (_GEN ? priorityReg : io_peAddress_valid);
	assign io_addressOut_valid = stateReg;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h0 ? 2'h2 : 2'h1);
			end
			else if (_GEN_0 | ~(_GEN_1 & io_vasAddressOut_ready))
				;
			else
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_1 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h1 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_2 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h2 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_3 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h3 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_4 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h4 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_5 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h5 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_6 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h6 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_7 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h7 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_8 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h8 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_9 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'h9 ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_10 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'ha ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_11 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'hb ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_12 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'hc ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_13 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'hd ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_14 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (io_addressIn_bits[7:4] == 4'he ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierServerNetworkUnit_15 (
	clock,
	reset,
	io_addressIn_ready,
	io_addressIn_valid,
	io_addressIn_bits,
	io_vasAddressOut_ready,
	io_vasAddressOut_valid,
	io_vasAddressOut_bits,
	io_addressOut_ready,
	io_addressOut_valid,
	io_addressOut_bits
);
	input clock;
	input reset;
	output wire io_addressIn_ready;
	input io_addressIn_valid;
	input [63:0] io_addressIn_bits;
	input io_vasAddressOut_ready;
	output wire io_vasAddressOut_valid;
	output wire [63:0] io_vasAddressOut_bits;
	input io_addressOut_ready;
	output wire io_addressOut_valid;
	output wire [63:0] io_addressOut_bits;
	reg [1:0] stateReg;
	reg [63:0] addressReg;
	wire _GEN = stateReg == 2'h0;
	wire _GEN_0 = stateReg == 2'h1;
	wire _GEN_1 = stateReg == 2'h2;
	always @(posedge clock)
		if (reset) begin
			stateReg <= 2'h0;
			addressReg <= 64'h0000000000000000;
		end
		else begin
			if (_GEN) begin
				if (io_addressIn_valid)
					stateReg <= (&io_addressIn_bits[7:4] ? 2'h2 : 2'h1);
			end
			else if ((_GEN_0 ? io_addressOut_ready : _GEN_1 & io_vasAddressOut_ready))
				stateReg <= 2'h0;
			if (_GEN & io_addressIn_valid)
				addressReg <= io_addressIn_bits;
		end
	assign io_addressIn_ready = _GEN;
	assign io_vasAddressOut_valid = ~(_GEN | _GEN_0) & _GEN_1;
	assign io_vasAddressOut_bits = addressReg;
	assign io_addressOut_valid = ~_GEN & _GEN_0;
	assign io_addressOut_bits = addressReg;
endmodule
module ArgumentNotifierNetwork (
	clock,
	reset,
	io_connVAS_0_ready,
	io_connVAS_0_valid,
	io_connVAS_0_bits,
	io_connVAS_1_ready,
	io_connVAS_1_valid,
	io_connVAS_1_bits,
	io_connVAS_2_ready,
	io_connVAS_2_valid,
	io_connVAS_2_bits,
	io_connVAS_3_ready,
	io_connVAS_3_valid,
	io_connVAS_3_bits,
	io_connVAS_4_ready,
	io_connVAS_4_valid,
	io_connVAS_4_bits,
	io_connVAS_5_ready,
	io_connVAS_5_valid,
	io_connVAS_5_bits,
	io_connVAS_6_ready,
	io_connVAS_6_valid,
	io_connVAS_6_bits,
	io_connVAS_7_ready,
	io_connVAS_7_valid,
	io_connVAS_7_bits,
	io_connVAS_8_ready,
	io_connVAS_8_valid,
	io_connVAS_8_bits,
	io_connVAS_9_ready,
	io_connVAS_9_valid,
	io_connVAS_9_bits,
	io_connVAS_10_ready,
	io_connVAS_10_valid,
	io_connVAS_10_bits,
	io_connVAS_11_ready,
	io_connVAS_11_valid,
	io_connVAS_11_bits,
	io_connVAS_12_ready,
	io_connVAS_12_valid,
	io_connVAS_12_bits,
	io_connVAS_13_ready,
	io_connVAS_13_valid,
	io_connVAS_13_bits,
	io_connVAS_14_ready,
	io_connVAS_14_valid,
	io_connVAS_14_bits,
	io_connVAS_15_ready,
	io_connVAS_15_valid,
	io_connVAS_15_bits,
	io_connPE_0_ready,
	io_connPE_0_valid,
	io_connPE_0_bits,
	io_connPE_1_ready,
	io_connPE_1_valid,
	io_connPE_1_bits,
	io_connPE_2_ready,
	io_connPE_2_valid,
	io_connPE_2_bits,
	io_connPE_3_ready,
	io_connPE_3_valid,
	io_connPE_3_bits,
	io_connPE_4_ready,
	io_connPE_4_valid,
	io_connPE_4_bits,
	io_connPE_5_ready,
	io_connPE_5_valid,
	io_connPE_5_bits,
	io_connPE_6_ready,
	io_connPE_6_valid,
	io_connPE_6_bits,
	io_connPE_7_ready,
	io_connPE_7_valid,
	io_connPE_7_bits,
	io_connPE_8_ready,
	io_connPE_8_valid,
	io_connPE_8_bits,
	io_connPE_9_ready,
	io_connPE_9_valid,
	io_connPE_9_bits,
	io_connPE_10_ready,
	io_connPE_10_valid,
	io_connPE_10_bits,
	io_connPE_11_ready,
	io_connPE_11_valid,
	io_connPE_11_bits,
	io_connPE_12_ready,
	io_connPE_12_valid,
	io_connPE_12_bits,
	io_connPE_13_ready,
	io_connPE_13_valid,
	io_connPE_13_bits,
	io_connPE_14_ready,
	io_connPE_14_valid,
	io_connPE_14_bits,
	io_connPE_15_ready,
	io_connPE_15_valid,
	io_connPE_15_bits,
	io_connPE_16_ready,
	io_connPE_16_valid,
	io_connPE_16_bits,
	io_connPE_17_ready,
	io_connPE_17_valid,
	io_connPE_17_bits,
	io_connPE_18_ready,
	io_connPE_18_valid,
	io_connPE_18_bits,
	io_connPE_19_ready,
	io_connPE_19_valid,
	io_connPE_19_bits,
	io_connPE_20_ready,
	io_connPE_20_valid,
	io_connPE_20_bits,
	io_connPE_21_ready,
	io_connPE_21_valid,
	io_connPE_21_bits,
	io_connPE_22_ready,
	io_connPE_22_valid,
	io_connPE_22_bits,
	io_connPE_23_ready,
	io_connPE_23_valid,
	io_connPE_23_bits,
	io_connPE_24_ready,
	io_connPE_24_valid,
	io_connPE_24_bits,
	io_connPE_25_ready,
	io_connPE_25_valid,
	io_connPE_25_bits,
	io_connPE_26_ready,
	io_connPE_26_valid,
	io_connPE_26_bits,
	io_connPE_27_ready,
	io_connPE_27_valid,
	io_connPE_27_bits,
	io_connPE_28_ready,
	io_connPE_28_valid,
	io_connPE_28_bits,
	io_connPE_29_ready,
	io_connPE_29_valid,
	io_connPE_29_bits,
	io_connPE_30_ready,
	io_connPE_30_valid,
	io_connPE_30_bits,
	io_connPE_31_ready,
	io_connPE_31_valid,
	io_connPE_31_bits,
	io_connPE_32_ready,
	io_connPE_32_valid,
	io_connPE_32_bits,
	io_connPE_33_ready,
	io_connPE_33_valid,
	io_connPE_33_bits,
	io_connPE_34_ready,
	io_connPE_34_valid,
	io_connPE_34_bits,
	io_connPE_35_ready,
	io_connPE_35_valid,
	io_connPE_35_bits,
	io_connPE_36_ready,
	io_connPE_36_valid,
	io_connPE_36_bits,
	io_connPE_37_ready,
	io_connPE_37_valid,
	io_connPE_37_bits,
	io_connPE_38_ready,
	io_connPE_38_valid,
	io_connPE_38_bits,
	io_connPE_39_ready,
	io_connPE_39_valid,
	io_connPE_39_bits,
	io_connPE_40_ready,
	io_connPE_40_valid,
	io_connPE_40_bits,
	io_connPE_41_ready,
	io_connPE_41_valid,
	io_connPE_41_bits,
	io_connPE_42_ready,
	io_connPE_42_valid,
	io_connPE_42_bits,
	io_connPE_43_ready,
	io_connPE_43_valid,
	io_connPE_43_bits,
	io_connPE_44_ready,
	io_connPE_44_valid,
	io_connPE_44_bits,
	io_connPE_45_ready,
	io_connPE_45_valid,
	io_connPE_45_bits,
	io_connPE_46_ready,
	io_connPE_46_valid,
	io_connPE_46_bits,
	io_connPE_47_ready,
	io_connPE_47_valid,
	io_connPE_47_bits,
	io_connPE_48_ready,
	io_connPE_48_valid,
	io_connPE_48_bits,
	io_connPE_49_ready,
	io_connPE_49_valid,
	io_connPE_49_bits,
	io_connPE_50_ready,
	io_connPE_50_valid,
	io_connPE_50_bits,
	io_connPE_51_ready,
	io_connPE_51_valid,
	io_connPE_51_bits,
	io_connPE_52_ready,
	io_connPE_52_valid,
	io_connPE_52_bits,
	io_connPE_53_ready,
	io_connPE_53_valid,
	io_connPE_53_bits,
	io_connPE_54_ready,
	io_connPE_54_valid,
	io_connPE_54_bits,
	io_connPE_55_ready,
	io_connPE_55_valid,
	io_connPE_55_bits,
	io_connPE_56_ready,
	io_connPE_56_valid,
	io_connPE_56_bits,
	io_connPE_57_ready,
	io_connPE_57_valid,
	io_connPE_57_bits,
	io_connPE_58_ready,
	io_connPE_58_valid,
	io_connPE_58_bits,
	io_connPE_59_ready,
	io_connPE_59_valid,
	io_connPE_59_bits,
	io_connPE_60_ready,
	io_connPE_60_valid,
	io_connPE_60_bits,
	io_connPE_61_ready,
	io_connPE_61_valid,
	io_connPE_61_bits,
	io_connPE_62_ready,
	io_connPE_62_valid,
	io_connPE_62_bits,
	io_connPE_63_ready,
	io_connPE_63_valid,
	io_connPE_63_bits,
	io_connPE_64_ready,
	io_connPE_64_valid,
	io_connPE_64_bits,
	io_connPE_65_ready,
	io_connPE_65_valid,
	io_connPE_65_bits,
	io_connPE_66_ready,
	io_connPE_66_valid,
	io_connPE_66_bits,
	io_connPE_67_ready,
	io_connPE_67_valid,
	io_connPE_67_bits,
	io_connPE_68_ready,
	io_connPE_68_valid,
	io_connPE_68_bits,
	io_connPE_69_ready,
	io_connPE_69_valid,
	io_connPE_69_bits,
	io_connPE_70_ready,
	io_connPE_70_valid,
	io_connPE_70_bits,
	io_connPE_71_ready,
	io_connPE_71_valid,
	io_connPE_71_bits,
	io_connPE_72_ready,
	io_connPE_72_valid,
	io_connPE_72_bits,
	io_connPE_73_ready,
	io_connPE_73_valid,
	io_connPE_73_bits,
	io_connPE_74_ready,
	io_connPE_74_valid,
	io_connPE_74_bits,
	io_connPE_75_ready,
	io_connPE_75_valid,
	io_connPE_75_bits,
	io_connPE_76_ready,
	io_connPE_76_valid,
	io_connPE_76_bits,
	io_connPE_77_ready,
	io_connPE_77_valid,
	io_connPE_77_bits,
	io_connPE_78_ready,
	io_connPE_78_valid,
	io_connPE_78_bits,
	io_connPE_79_ready,
	io_connPE_79_valid,
	io_connPE_79_bits
);
	input clock;
	input reset;
	input io_connVAS_0_ready;
	output wire io_connVAS_0_valid;
	output wire [63:0] io_connVAS_0_bits;
	input io_connVAS_1_ready;
	output wire io_connVAS_1_valid;
	output wire [63:0] io_connVAS_1_bits;
	input io_connVAS_2_ready;
	output wire io_connVAS_2_valid;
	output wire [63:0] io_connVAS_2_bits;
	input io_connVAS_3_ready;
	output wire io_connVAS_3_valid;
	output wire [63:0] io_connVAS_3_bits;
	input io_connVAS_4_ready;
	output wire io_connVAS_4_valid;
	output wire [63:0] io_connVAS_4_bits;
	input io_connVAS_5_ready;
	output wire io_connVAS_5_valid;
	output wire [63:0] io_connVAS_5_bits;
	input io_connVAS_6_ready;
	output wire io_connVAS_6_valid;
	output wire [63:0] io_connVAS_6_bits;
	input io_connVAS_7_ready;
	output wire io_connVAS_7_valid;
	output wire [63:0] io_connVAS_7_bits;
	input io_connVAS_8_ready;
	output wire io_connVAS_8_valid;
	output wire [63:0] io_connVAS_8_bits;
	input io_connVAS_9_ready;
	output wire io_connVAS_9_valid;
	output wire [63:0] io_connVAS_9_bits;
	input io_connVAS_10_ready;
	output wire io_connVAS_10_valid;
	output wire [63:0] io_connVAS_10_bits;
	input io_connVAS_11_ready;
	output wire io_connVAS_11_valid;
	output wire [63:0] io_connVAS_11_bits;
	input io_connVAS_12_ready;
	output wire io_connVAS_12_valid;
	output wire [63:0] io_connVAS_12_bits;
	input io_connVAS_13_ready;
	output wire io_connVAS_13_valid;
	output wire [63:0] io_connVAS_13_bits;
	input io_connVAS_14_ready;
	output wire io_connVAS_14_valid;
	output wire [63:0] io_connVAS_14_bits;
	input io_connVAS_15_ready;
	output wire io_connVAS_15_valid;
	output wire [63:0] io_connVAS_15_bits;
	output wire io_connPE_0_ready;
	input io_connPE_0_valid;
	input [63:0] io_connPE_0_bits;
	output wire io_connPE_1_ready;
	input io_connPE_1_valid;
	input [63:0] io_connPE_1_bits;
	output wire io_connPE_2_ready;
	input io_connPE_2_valid;
	input [63:0] io_connPE_2_bits;
	output wire io_connPE_3_ready;
	input io_connPE_3_valid;
	input [63:0] io_connPE_3_bits;
	output wire io_connPE_4_ready;
	input io_connPE_4_valid;
	input [63:0] io_connPE_4_bits;
	output wire io_connPE_5_ready;
	input io_connPE_5_valid;
	input [63:0] io_connPE_5_bits;
	output wire io_connPE_6_ready;
	input io_connPE_6_valid;
	input [63:0] io_connPE_6_bits;
	output wire io_connPE_7_ready;
	input io_connPE_7_valid;
	input [63:0] io_connPE_7_bits;
	output wire io_connPE_8_ready;
	input io_connPE_8_valid;
	input [63:0] io_connPE_8_bits;
	output wire io_connPE_9_ready;
	input io_connPE_9_valid;
	input [63:0] io_connPE_9_bits;
	output wire io_connPE_10_ready;
	input io_connPE_10_valid;
	input [63:0] io_connPE_10_bits;
	output wire io_connPE_11_ready;
	input io_connPE_11_valid;
	input [63:0] io_connPE_11_bits;
	output wire io_connPE_12_ready;
	input io_connPE_12_valid;
	input [63:0] io_connPE_12_bits;
	output wire io_connPE_13_ready;
	input io_connPE_13_valid;
	input [63:0] io_connPE_13_bits;
	output wire io_connPE_14_ready;
	input io_connPE_14_valid;
	input [63:0] io_connPE_14_bits;
	output wire io_connPE_15_ready;
	input io_connPE_15_valid;
	input [63:0] io_connPE_15_bits;
	output wire io_connPE_16_ready;
	input io_connPE_16_valid;
	input [63:0] io_connPE_16_bits;
	output wire io_connPE_17_ready;
	input io_connPE_17_valid;
	input [63:0] io_connPE_17_bits;
	output wire io_connPE_18_ready;
	input io_connPE_18_valid;
	input [63:0] io_connPE_18_bits;
	output wire io_connPE_19_ready;
	input io_connPE_19_valid;
	input [63:0] io_connPE_19_bits;
	output wire io_connPE_20_ready;
	input io_connPE_20_valid;
	input [63:0] io_connPE_20_bits;
	output wire io_connPE_21_ready;
	input io_connPE_21_valid;
	input [63:0] io_connPE_21_bits;
	output wire io_connPE_22_ready;
	input io_connPE_22_valid;
	input [63:0] io_connPE_22_bits;
	output wire io_connPE_23_ready;
	input io_connPE_23_valid;
	input [63:0] io_connPE_23_bits;
	output wire io_connPE_24_ready;
	input io_connPE_24_valid;
	input [63:0] io_connPE_24_bits;
	output wire io_connPE_25_ready;
	input io_connPE_25_valid;
	input [63:0] io_connPE_25_bits;
	output wire io_connPE_26_ready;
	input io_connPE_26_valid;
	input [63:0] io_connPE_26_bits;
	output wire io_connPE_27_ready;
	input io_connPE_27_valid;
	input [63:0] io_connPE_27_bits;
	output wire io_connPE_28_ready;
	input io_connPE_28_valid;
	input [63:0] io_connPE_28_bits;
	output wire io_connPE_29_ready;
	input io_connPE_29_valid;
	input [63:0] io_connPE_29_bits;
	output wire io_connPE_30_ready;
	input io_connPE_30_valid;
	input [63:0] io_connPE_30_bits;
	output wire io_connPE_31_ready;
	input io_connPE_31_valid;
	input [63:0] io_connPE_31_bits;
	output wire io_connPE_32_ready;
	input io_connPE_32_valid;
	input [63:0] io_connPE_32_bits;
	output wire io_connPE_33_ready;
	input io_connPE_33_valid;
	input [63:0] io_connPE_33_bits;
	output wire io_connPE_34_ready;
	input io_connPE_34_valid;
	input [63:0] io_connPE_34_bits;
	output wire io_connPE_35_ready;
	input io_connPE_35_valid;
	input [63:0] io_connPE_35_bits;
	output wire io_connPE_36_ready;
	input io_connPE_36_valid;
	input [63:0] io_connPE_36_bits;
	output wire io_connPE_37_ready;
	input io_connPE_37_valid;
	input [63:0] io_connPE_37_bits;
	output wire io_connPE_38_ready;
	input io_connPE_38_valid;
	input [63:0] io_connPE_38_bits;
	output wire io_connPE_39_ready;
	input io_connPE_39_valid;
	input [63:0] io_connPE_39_bits;
	output wire io_connPE_40_ready;
	input io_connPE_40_valid;
	input [63:0] io_connPE_40_bits;
	output wire io_connPE_41_ready;
	input io_connPE_41_valid;
	input [63:0] io_connPE_41_bits;
	output wire io_connPE_42_ready;
	input io_connPE_42_valid;
	input [63:0] io_connPE_42_bits;
	output wire io_connPE_43_ready;
	input io_connPE_43_valid;
	input [63:0] io_connPE_43_bits;
	output wire io_connPE_44_ready;
	input io_connPE_44_valid;
	input [63:0] io_connPE_44_bits;
	output wire io_connPE_45_ready;
	input io_connPE_45_valid;
	input [63:0] io_connPE_45_bits;
	output wire io_connPE_46_ready;
	input io_connPE_46_valid;
	input [63:0] io_connPE_46_bits;
	output wire io_connPE_47_ready;
	input io_connPE_47_valid;
	input [63:0] io_connPE_47_bits;
	output wire io_connPE_48_ready;
	input io_connPE_48_valid;
	input [63:0] io_connPE_48_bits;
	output wire io_connPE_49_ready;
	input io_connPE_49_valid;
	input [63:0] io_connPE_49_bits;
	output wire io_connPE_50_ready;
	input io_connPE_50_valid;
	input [63:0] io_connPE_50_bits;
	output wire io_connPE_51_ready;
	input io_connPE_51_valid;
	input [63:0] io_connPE_51_bits;
	output wire io_connPE_52_ready;
	input io_connPE_52_valid;
	input [63:0] io_connPE_52_bits;
	output wire io_connPE_53_ready;
	input io_connPE_53_valid;
	input [63:0] io_connPE_53_bits;
	output wire io_connPE_54_ready;
	input io_connPE_54_valid;
	input [63:0] io_connPE_54_bits;
	output wire io_connPE_55_ready;
	input io_connPE_55_valid;
	input [63:0] io_connPE_55_bits;
	output wire io_connPE_56_ready;
	input io_connPE_56_valid;
	input [63:0] io_connPE_56_bits;
	output wire io_connPE_57_ready;
	input io_connPE_57_valid;
	input [63:0] io_connPE_57_bits;
	output wire io_connPE_58_ready;
	input io_connPE_58_valid;
	input [63:0] io_connPE_58_bits;
	output wire io_connPE_59_ready;
	input io_connPE_59_valid;
	input [63:0] io_connPE_59_bits;
	output wire io_connPE_60_ready;
	input io_connPE_60_valid;
	input [63:0] io_connPE_60_bits;
	output wire io_connPE_61_ready;
	input io_connPE_61_valid;
	input [63:0] io_connPE_61_bits;
	output wire io_connPE_62_ready;
	input io_connPE_62_valid;
	input [63:0] io_connPE_62_bits;
	output wire io_connPE_63_ready;
	input io_connPE_63_valid;
	input [63:0] io_connPE_63_bits;
	output wire io_connPE_64_ready;
	input io_connPE_64_valid;
	input [63:0] io_connPE_64_bits;
	output wire io_connPE_65_ready;
	input io_connPE_65_valid;
	input [63:0] io_connPE_65_bits;
	output wire io_connPE_66_ready;
	input io_connPE_66_valid;
	input [63:0] io_connPE_66_bits;
	output wire io_connPE_67_ready;
	input io_connPE_67_valid;
	input [63:0] io_connPE_67_bits;
	output wire io_connPE_68_ready;
	input io_connPE_68_valid;
	input [63:0] io_connPE_68_bits;
	output wire io_connPE_69_ready;
	input io_connPE_69_valid;
	input [63:0] io_connPE_69_bits;
	output wire io_connPE_70_ready;
	input io_connPE_70_valid;
	input [63:0] io_connPE_70_bits;
	output wire io_connPE_71_ready;
	input io_connPE_71_valid;
	input [63:0] io_connPE_71_bits;
	output wire io_connPE_72_ready;
	input io_connPE_72_valid;
	input [63:0] io_connPE_72_bits;
	output wire io_connPE_73_ready;
	input io_connPE_73_valid;
	input [63:0] io_connPE_73_bits;
	output wire io_connPE_74_ready;
	input io_connPE_74_valid;
	input [63:0] io_connPE_74_bits;
	output wire io_connPE_75_ready;
	input io_connPE_75_valid;
	input [63:0] io_connPE_75_bits;
	output wire io_connPE_76_ready;
	input io_connPE_76_valid;
	input [63:0] io_connPE_76_bits;
	output wire io_connPE_77_ready;
	input io_connPE_77_valid;
	input [63:0] io_connPE_77_bits;
	output wire io_connPE_78_ready;
	input io_connPE_78_valid;
	input [63:0] io_connPE_78_bits;
	output wire io_connPE_79_ready;
	input io_connPE_79_valid;
	input [63:0] io_connPE_79_bits;
	wire _queues_79_io_addressOut_valid;
	wire [63:0] _queues_79_io_addressOut_bits;
	wire _queues_78_io_addressOut_valid;
	wire [63:0] _queues_78_io_addressOut_bits;
	wire _queues_77_io_addressOut_valid;
	wire [63:0] _queues_77_io_addressOut_bits;
	wire _queues_76_io_addressOut_valid;
	wire [63:0] _queues_76_io_addressOut_bits;
	wire _queues_75_io_addressOut_valid;
	wire [63:0] _queues_75_io_addressOut_bits;
	wire _queues_74_io_addressOut_valid;
	wire [63:0] _queues_74_io_addressOut_bits;
	wire _queues_73_io_addressOut_valid;
	wire [63:0] _queues_73_io_addressOut_bits;
	wire _queues_72_io_addressOut_valid;
	wire [63:0] _queues_72_io_addressOut_bits;
	wire _queues_71_io_addressOut_valid;
	wire [63:0] _queues_71_io_addressOut_bits;
	wire _queues_70_io_addressOut_valid;
	wire [63:0] _queues_70_io_addressOut_bits;
	wire _queues_69_io_addressOut_valid;
	wire [63:0] _queues_69_io_addressOut_bits;
	wire _queues_68_io_addressOut_valid;
	wire [63:0] _queues_68_io_addressOut_bits;
	wire _queues_67_io_addressOut_valid;
	wire [63:0] _queues_67_io_addressOut_bits;
	wire _queues_66_io_addressOut_valid;
	wire [63:0] _queues_66_io_addressOut_bits;
	wire _queues_65_io_addressOut_valid;
	wire [63:0] _queues_65_io_addressOut_bits;
	wire _queues_64_io_addressOut_valid;
	wire [63:0] _queues_64_io_addressOut_bits;
	wire _queues_63_io_addressOut_valid;
	wire [63:0] _queues_63_io_addressOut_bits;
	wire _queues_62_io_addressOut_valid;
	wire [63:0] _queues_62_io_addressOut_bits;
	wire _queues_61_io_addressOut_valid;
	wire [63:0] _queues_61_io_addressOut_bits;
	wire _queues_60_io_addressOut_valid;
	wire [63:0] _queues_60_io_addressOut_bits;
	wire _queues_59_io_addressOut_valid;
	wire [63:0] _queues_59_io_addressOut_bits;
	wire _queues_58_io_addressOut_valid;
	wire [63:0] _queues_58_io_addressOut_bits;
	wire _queues_57_io_addressOut_valid;
	wire [63:0] _queues_57_io_addressOut_bits;
	wire _queues_56_io_addressOut_valid;
	wire [63:0] _queues_56_io_addressOut_bits;
	wire _queues_55_io_addressOut_valid;
	wire [63:0] _queues_55_io_addressOut_bits;
	wire _queues_54_io_addressOut_valid;
	wire [63:0] _queues_54_io_addressOut_bits;
	wire _queues_53_io_addressOut_valid;
	wire [63:0] _queues_53_io_addressOut_bits;
	wire _queues_52_io_addressOut_valid;
	wire [63:0] _queues_52_io_addressOut_bits;
	wire _queues_51_io_addressOut_valid;
	wire [63:0] _queues_51_io_addressOut_bits;
	wire _queues_50_io_addressOut_valid;
	wire [63:0] _queues_50_io_addressOut_bits;
	wire _queues_49_io_addressOut_valid;
	wire [63:0] _queues_49_io_addressOut_bits;
	wire _queues_48_io_addressOut_valid;
	wire [63:0] _queues_48_io_addressOut_bits;
	wire _queues_47_io_addressOut_valid;
	wire [63:0] _queues_47_io_addressOut_bits;
	wire _queues_46_io_addressOut_valid;
	wire [63:0] _queues_46_io_addressOut_bits;
	wire _queues_45_io_addressOut_valid;
	wire [63:0] _queues_45_io_addressOut_bits;
	wire _queues_44_io_addressOut_valid;
	wire [63:0] _queues_44_io_addressOut_bits;
	wire _queues_43_io_addressOut_valid;
	wire [63:0] _queues_43_io_addressOut_bits;
	wire _queues_42_io_addressOut_valid;
	wire [63:0] _queues_42_io_addressOut_bits;
	wire _queues_41_io_addressOut_valid;
	wire [63:0] _queues_41_io_addressOut_bits;
	wire _queues_40_io_addressOut_valid;
	wire [63:0] _queues_40_io_addressOut_bits;
	wire _queues_39_io_addressOut_valid;
	wire [63:0] _queues_39_io_addressOut_bits;
	wire _queues_38_io_addressOut_valid;
	wire [63:0] _queues_38_io_addressOut_bits;
	wire _queues_37_io_addressOut_valid;
	wire [63:0] _queues_37_io_addressOut_bits;
	wire _queues_36_io_addressOut_valid;
	wire [63:0] _queues_36_io_addressOut_bits;
	wire _queues_35_io_addressOut_valid;
	wire [63:0] _queues_35_io_addressOut_bits;
	wire _queues_34_io_addressOut_valid;
	wire [63:0] _queues_34_io_addressOut_bits;
	wire _queues_33_io_addressOut_valid;
	wire [63:0] _queues_33_io_addressOut_bits;
	wire _queues_32_io_addressOut_valid;
	wire [63:0] _queues_32_io_addressOut_bits;
	wire _queues_31_io_addressOut_valid;
	wire [63:0] _queues_31_io_addressOut_bits;
	wire _queues_30_io_addressOut_valid;
	wire [63:0] _queues_30_io_addressOut_bits;
	wire _queues_29_io_addressOut_valid;
	wire [63:0] _queues_29_io_addressOut_bits;
	wire _queues_28_io_addressOut_valid;
	wire [63:0] _queues_28_io_addressOut_bits;
	wire _queues_27_io_addressOut_valid;
	wire [63:0] _queues_27_io_addressOut_bits;
	wire _queues_26_io_addressOut_valid;
	wire [63:0] _queues_26_io_addressOut_bits;
	wire _queues_25_io_addressOut_valid;
	wire [63:0] _queues_25_io_addressOut_bits;
	wire _queues_24_io_addressOut_valid;
	wire [63:0] _queues_24_io_addressOut_bits;
	wire _queues_23_io_addressOut_valid;
	wire [63:0] _queues_23_io_addressOut_bits;
	wire _queues_22_io_addressOut_valid;
	wire [63:0] _queues_22_io_addressOut_bits;
	wire _queues_21_io_addressOut_valid;
	wire [63:0] _queues_21_io_addressOut_bits;
	wire _queues_20_io_addressOut_valid;
	wire [63:0] _queues_20_io_addressOut_bits;
	wire _queues_19_io_addressOut_valid;
	wire [63:0] _queues_19_io_addressOut_bits;
	wire _queues_18_io_addressOut_valid;
	wire [63:0] _queues_18_io_addressOut_bits;
	wire _queues_17_io_addressOut_valid;
	wire [63:0] _queues_17_io_addressOut_bits;
	wire _queues_16_io_addressOut_valid;
	wire [63:0] _queues_16_io_addressOut_bits;
	wire _queues_15_io_addressOut_valid;
	wire [63:0] _queues_15_io_addressOut_bits;
	wire _queues_14_io_addressOut_valid;
	wire [63:0] _queues_14_io_addressOut_bits;
	wire _queues_13_io_addressOut_valid;
	wire [63:0] _queues_13_io_addressOut_bits;
	wire _queues_12_io_addressOut_valid;
	wire [63:0] _queues_12_io_addressOut_bits;
	wire _queues_11_io_addressOut_valid;
	wire [63:0] _queues_11_io_addressOut_bits;
	wire _queues_10_io_addressOut_valid;
	wire [63:0] _queues_10_io_addressOut_bits;
	wire _queues_9_io_addressOut_valid;
	wire [63:0] _queues_9_io_addressOut_bits;
	wire _queues_8_io_addressOut_valid;
	wire [63:0] _queues_8_io_addressOut_bits;
	wire _queues_7_io_addressOut_valid;
	wire [63:0] _queues_7_io_addressOut_bits;
	wire _queues_6_io_addressOut_valid;
	wire [63:0] _queues_6_io_addressOut_bits;
	wire _queues_5_io_addressOut_valid;
	wire [63:0] _queues_5_io_addressOut_bits;
	wire _queues_4_io_addressOut_valid;
	wire [63:0] _queues_4_io_addressOut_bits;
	wire _queues_3_io_addressOut_valid;
	wire [63:0] _queues_3_io_addressOut_bits;
	wire _queues_2_io_addressOut_valid;
	wire [63:0] _queues_2_io_addressOut_bits;
	wire _queues_1_io_addressOut_valid;
	wire [63:0] _queues_1_io_addressOut_bits;
	wire _queues_0_io_addressOut_valid;
	wire [63:0] _queues_0_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_15_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_15_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_15_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_14_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_14_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_14_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_13_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_13_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_13_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_12_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_12_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_12_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_11_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_11_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_11_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_10_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_10_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_10_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_9_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_9_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_9_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_8_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_8_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_8_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_7_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_7_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_7_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_6_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_6_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_6_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_5_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_5_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_5_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_4_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_4_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_4_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_3_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_3_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_3_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_2_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_2_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_2_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_1_io_addressIn_ready;
	wire _ArgumentNotifierServerNetworkUnit_1_io_addressOut_valid;
	wire [63:0] _ArgumentNotifierServerNetworkUnit_1_io_addressOut_bits;
	wire _ArgumentNotifierServerNetworkUnit_io_addressIn_ready;
	wire _networkUnits_79_io_peAddress_ready;
	wire _networkUnits_79_io_addressOut_valid;
	wire [63:0] _networkUnits_79_io_addressOut_bits;
	wire _networkUnits_78_io_addressIn_ready;
	wire _networkUnits_78_io_peAddress_ready;
	wire _networkUnits_78_io_addressOut_valid;
	wire [63:0] _networkUnits_78_io_addressOut_bits;
	wire _networkUnits_77_io_addressIn_ready;
	wire _networkUnits_77_io_peAddress_ready;
	wire _networkUnits_77_io_addressOut_valid;
	wire [63:0] _networkUnits_77_io_addressOut_bits;
	wire _networkUnits_76_io_addressIn_ready;
	wire _networkUnits_76_io_peAddress_ready;
	wire _networkUnits_76_io_addressOut_valid;
	wire [63:0] _networkUnits_76_io_addressOut_bits;
	wire _networkUnits_75_io_addressIn_ready;
	wire _networkUnits_75_io_peAddress_ready;
	wire _networkUnits_75_io_addressOut_valid;
	wire [63:0] _networkUnits_75_io_addressOut_bits;
	wire _networkUnits_74_io_addressIn_ready;
	wire _networkUnits_74_io_peAddress_ready;
	wire _networkUnits_74_io_addressOut_valid;
	wire [63:0] _networkUnits_74_io_addressOut_bits;
	wire _networkUnits_73_io_addressIn_ready;
	wire _networkUnits_73_io_peAddress_ready;
	wire _networkUnits_73_io_addressOut_valid;
	wire [63:0] _networkUnits_73_io_addressOut_bits;
	wire _networkUnits_72_io_addressIn_ready;
	wire _networkUnits_72_io_peAddress_ready;
	wire _networkUnits_72_io_addressOut_valid;
	wire [63:0] _networkUnits_72_io_addressOut_bits;
	wire _networkUnits_71_io_addressIn_ready;
	wire _networkUnits_71_io_peAddress_ready;
	wire _networkUnits_71_io_addressOut_valid;
	wire [63:0] _networkUnits_71_io_addressOut_bits;
	wire _networkUnits_70_io_addressIn_ready;
	wire _networkUnits_70_io_peAddress_ready;
	wire _networkUnits_70_io_addressOut_valid;
	wire [63:0] _networkUnits_70_io_addressOut_bits;
	wire _networkUnits_69_io_addressIn_ready;
	wire _networkUnits_69_io_peAddress_ready;
	wire _networkUnits_69_io_addressOut_valid;
	wire [63:0] _networkUnits_69_io_addressOut_bits;
	wire _networkUnits_68_io_addressIn_ready;
	wire _networkUnits_68_io_peAddress_ready;
	wire _networkUnits_68_io_addressOut_valid;
	wire [63:0] _networkUnits_68_io_addressOut_bits;
	wire _networkUnits_67_io_addressIn_ready;
	wire _networkUnits_67_io_peAddress_ready;
	wire _networkUnits_67_io_addressOut_valid;
	wire [63:0] _networkUnits_67_io_addressOut_bits;
	wire _networkUnits_66_io_addressIn_ready;
	wire _networkUnits_66_io_peAddress_ready;
	wire _networkUnits_66_io_addressOut_valid;
	wire [63:0] _networkUnits_66_io_addressOut_bits;
	wire _networkUnits_65_io_addressIn_ready;
	wire _networkUnits_65_io_peAddress_ready;
	wire _networkUnits_65_io_addressOut_valid;
	wire [63:0] _networkUnits_65_io_addressOut_bits;
	wire _networkUnits_64_io_addressIn_ready;
	wire _networkUnits_64_io_peAddress_ready;
	wire _networkUnits_64_io_addressOut_valid;
	wire [63:0] _networkUnits_64_io_addressOut_bits;
	wire _networkUnits_63_io_addressIn_ready;
	wire _networkUnits_63_io_peAddress_ready;
	wire _networkUnits_63_io_addressOut_valid;
	wire [63:0] _networkUnits_63_io_addressOut_bits;
	wire _networkUnits_62_io_addressIn_ready;
	wire _networkUnits_62_io_peAddress_ready;
	wire _networkUnits_62_io_addressOut_valid;
	wire [63:0] _networkUnits_62_io_addressOut_bits;
	wire _networkUnits_61_io_addressIn_ready;
	wire _networkUnits_61_io_peAddress_ready;
	wire _networkUnits_61_io_addressOut_valid;
	wire [63:0] _networkUnits_61_io_addressOut_bits;
	wire _networkUnits_60_io_addressIn_ready;
	wire _networkUnits_60_io_peAddress_ready;
	wire _networkUnits_60_io_addressOut_valid;
	wire [63:0] _networkUnits_60_io_addressOut_bits;
	wire _networkUnits_59_io_addressIn_ready;
	wire _networkUnits_59_io_peAddress_ready;
	wire _networkUnits_59_io_addressOut_valid;
	wire [63:0] _networkUnits_59_io_addressOut_bits;
	wire _networkUnits_58_io_addressIn_ready;
	wire _networkUnits_58_io_peAddress_ready;
	wire _networkUnits_58_io_addressOut_valid;
	wire [63:0] _networkUnits_58_io_addressOut_bits;
	wire _networkUnits_57_io_addressIn_ready;
	wire _networkUnits_57_io_peAddress_ready;
	wire _networkUnits_57_io_addressOut_valid;
	wire [63:0] _networkUnits_57_io_addressOut_bits;
	wire _networkUnits_56_io_addressIn_ready;
	wire _networkUnits_56_io_peAddress_ready;
	wire _networkUnits_56_io_addressOut_valid;
	wire [63:0] _networkUnits_56_io_addressOut_bits;
	wire _networkUnits_55_io_addressIn_ready;
	wire _networkUnits_55_io_peAddress_ready;
	wire _networkUnits_55_io_addressOut_valid;
	wire [63:0] _networkUnits_55_io_addressOut_bits;
	wire _networkUnits_54_io_addressIn_ready;
	wire _networkUnits_54_io_peAddress_ready;
	wire _networkUnits_54_io_addressOut_valid;
	wire [63:0] _networkUnits_54_io_addressOut_bits;
	wire _networkUnits_53_io_addressIn_ready;
	wire _networkUnits_53_io_peAddress_ready;
	wire _networkUnits_53_io_addressOut_valid;
	wire [63:0] _networkUnits_53_io_addressOut_bits;
	wire _networkUnits_52_io_addressIn_ready;
	wire _networkUnits_52_io_peAddress_ready;
	wire _networkUnits_52_io_addressOut_valid;
	wire [63:0] _networkUnits_52_io_addressOut_bits;
	wire _networkUnits_51_io_addressIn_ready;
	wire _networkUnits_51_io_peAddress_ready;
	wire _networkUnits_51_io_addressOut_valid;
	wire [63:0] _networkUnits_51_io_addressOut_bits;
	wire _networkUnits_50_io_addressIn_ready;
	wire _networkUnits_50_io_peAddress_ready;
	wire _networkUnits_50_io_addressOut_valid;
	wire [63:0] _networkUnits_50_io_addressOut_bits;
	wire _networkUnits_49_io_addressIn_ready;
	wire _networkUnits_49_io_peAddress_ready;
	wire _networkUnits_49_io_addressOut_valid;
	wire [63:0] _networkUnits_49_io_addressOut_bits;
	wire _networkUnits_48_io_addressIn_ready;
	wire _networkUnits_48_io_peAddress_ready;
	wire _networkUnits_48_io_addressOut_valid;
	wire [63:0] _networkUnits_48_io_addressOut_bits;
	wire _networkUnits_47_io_addressIn_ready;
	wire _networkUnits_47_io_peAddress_ready;
	wire _networkUnits_47_io_addressOut_valid;
	wire [63:0] _networkUnits_47_io_addressOut_bits;
	wire _networkUnits_46_io_addressIn_ready;
	wire _networkUnits_46_io_peAddress_ready;
	wire _networkUnits_46_io_addressOut_valid;
	wire [63:0] _networkUnits_46_io_addressOut_bits;
	wire _networkUnits_45_io_addressIn_ready;
	wire _networkUnits_45_io_peAddress_ready;
	wire _networkUnits_45_io_addressOut_valid;
	wire [63:0] _networkUnits_45_io_addressOut_bits;
	wire _networkUnits_44_io_addressIn_ready;
	wire _networkUnits_44_io_peAddress_ready;
	wire _networkUnits_44_io_addressOut_valid;
	wire [63:0] _networkUnits_44_io_addressOut_bits;
	wire _networkUnits_43_io_addressIn_ready;
	wire _networkUnits_43_io_peAddress_ready;
	wire _networkUnits_43_io_addressOut_valid;
	wire [63:0] _networkUnits_43_io_addressOut_bits;
	wire _networkUnits_42_io_addressIn_ready;
	wire _networkUnits_42_io_peAddress_ready;
	wire _networkUnits_42_io_addressOut_valid;
	wire [63:0] _networkUnits_42_io_addressOut_bits;
	wire _networkUnits_41_io_addressIn_ready;
	wire _networkUnits_41_io_peAddress_ready;
	wire _networkUnits_41_io_addressOut_valid;
	wire [63:0] _networkUnits_41_io_addressOut_bits;
	wire _networkUnits_40_io_addressIn_ready;
	wire _networkUnits_40_io_peAddress_ready;
	wire _networkUnits_40_io_addressOut_valid;
	wire [63:0] _networkUnits_40_io_addressOut_bits;
	wire _networkUnits_39_io_addressIn_ready;
	wire _networkUnits_39_io_peAddress_ready;
	wire _networkUnits_39_io_addressOut_valid;
	wire [63:0] _networkUnits_39_io_addressOut_bits;
	wire _networkUnits_38_io_addressIn_ready;
	wire _networkUnits_38_io_peAddress_ready;
	wire _networkUnits_38_io_addressOut_valid;
	wire [63:0] _networkUnits_38_io_addressOut_bits;
	wire _networkUnits_37_io_addressIn_ready;
	wire _networkUnits_37_io_peAddress_ready;
	wire _networkUnits_37_io_addressOut_valid;
	wire [63:0] _networkUnits_37_io_addressOut_bits;
	wire _networkUnits_36_io_addressIn_ready;
	wire _networkUnits_36_io_peAddress_ready;
	wire _networkUnits_36_io_addressOut_valid;
	wire [63:0] _networkUnits_36_io_addressOut_bits;
	wire _networkUnits_35_io_addressIn_ready;
	wire _networkUnits_35_io_peAddress_ready;
	wire _networkUnits_35_io_addressOut_valid;
	wire [63:0] _networkUnits_35_io_addressOut_bits;
	wire _networkUnits_34_io_addressIn_ready;
	wire _networkUnits_34_io_peAddress_ready;
	wire _networkUnits_34_io_addressOut_valid;
	wire [63:0] _networkUnits_34_io_addressOut_bits;
	wire _networkUnits_33_io_addressIn_ready;
	wire _networkUnits_33_io_peAddress_ready;
	wire _networkUnits_33_io_addressOut_valid;
	wire [63:0] _networkUnits_33_io_addressOut_bits;
	wire _networkUnits_32_io_addressIn_ready;
	wire _networkUnits_32_io_peAddress_ready;
	wire _networkUnits_32_io_addressOut_valid;
	wire [63:0] _networkUnits_32_io_addressOut_bits;
	wire _networkUnits_31_io_addressIn_ready;
	wire _networkUnits_31_io_peAddress_ready;
	wire _networkUnits_31_io_addressOut_valid;
	wire [63:0] _networkUnits_31_io_addressOut_bits;
	wire _networkUnits_30_io_addressIn_ready;
	wire _networkUnits_30_io_peAddress_ready;
	wire _networkUnits_30_io_addressOut_valid;
	wire [63:0] _networkUnits_30_io_addressOut_bits;
	wire _networkUnits_29_io_addressIn_ready;
	wire _networkUnits_29_io_peAddress_ready;
	wire _networkUnits_29_io_addressOut_valid;
	wire [63:0] _networkUnits_29_io_addressOut_bits;
	wire _networkUnits_28_io_addressIn_ready;
	wire _networkUnits_28_io_peAddress_ready;
	wire _networkUnits_28_io_addressOut_valid;
	wire [63:0] _networkUnits_28_io_addressOut_bits;
	wire _networkUnits_27_io_addressIn_ready;
	wire _networkUnits_27_io_peAddress_ready;
	wire _networkUnits_27_io_addressOut_valid;
	wire [63:0] _networkUnits_27_io_addressOut_bits;
	wire _networkUnits_26_io_addressIn_ready;
	wire _networkUnits_26_io_peAddress_ready;
	wire _networkUnits_26_io_addressOut_valid;
	wire [63:0] _networkUnits_26_io_addressOut_bits;
	wire _networkUnits_25_io_addressIn_ready;
	wire _networkUnits_25_io_peAddress_ready;
	wire _networkUnits_25_io_addressOut_valid;
	wire [63:0] _networkUnits_25_io_addressOut_bits;
	wire _networkUnits_24_io_addressIn_ready;
	wire _networkUnits_24_io_peAddress_ready;
	wire _networkUnits_24_io_addressOut_valid;
	wire [63:0] _networkUnits_24_io_addressOut_bits;
	wire _networkUnits_23_io_addressIn_ready;
	wire _networkUnits_23_io_peAddress_ready;
	wire _networkUnits_23_io_addressOut_valid;
	wire [63:0] _networkUnits_23_io_addressOut_bits;
	wire _networkUnits_22_io_addressIn_ready;
	wire _networkUnits_22_io_peAddress_ready;
	wire _networkUnits_22_io_addressOut_valid;
	wire [63:0] _networkUnits_22_io_addressOut_bits;
	wire _networkUnits_21_io_addressIn_ready;
	wire _networkUnits_21_io_peAddress_ready;
	wire _networkUnits_21_io_addressOut_valid;
	wire [63:0] _networkUnits_21_io_addressOut_bits;
	wire _networkUnits_20_io_addressIn_ready;
	wire _networkUnits_20_io_peAddress_ready;
	wire _networkUnits_20_io_addressOut_valid;
	wire [63:0] _networkUnits_20_io_addressOut_bits;
	wire _networkUnits_19_io_addressIn_ready;
	wire _networkUnits_19_io_peAddress_ready;
	wire _networkUnits_19_io_addressOut_valid;
	wire [63:0] _networkUnits_19_io_addressOut_bits;
	wire _networkUnits_18_io_addressIn_ready;
	wire _networkUnits_18_io_peAddress_ready;
	wire _networkUnits_18_io_addressOut_valid;
	wire [63:0] _networkUnits_18_io_addressOut_bits;
	wire _networkUnits_17_io_addressIn_ready;
	wire _networkUnits_17_io_peAddress_ready;
	wire _networkUnits_17_io_addressOut_valid;
	wire [63:0] _networkUnits_17_io_addressOut_bits;
	wire _networkUnits_16_io_addressIn_ready;
	wire _networkUnits_16_io_peAddress_ready;
	wire _networkUnits_16_io_addressOut_valid;
	wire [63:0] _networkUnits_16_io_addressOut_bits;
	wire _networkUnits_15_io_addressIn_ready;
	wire _networkUnits_15_io_peAddress_ready;
	wire _networkUnits_15_io_addressOut_valid;
	wire [63:0] _networkUnits_15_io_addressOut_bits;
	wire _networkUnits_14_io_addressIn_ready;
	wire _networkUnits_14_io_peAddress_ready;
	wire _networkUnits_14_io_addressOut_valid;
	wire [63:0] _networkUnits_14_io_addressOut_bits;
	wire _networkUnits_13_io_addressIn_ready;
	wire _networkUnits_13_io_peAddress_ready;
	wire _networkUnits_13_io_addressOut_valid;
	wire [63:0] _networkUnits_13_io_addressOut_bits;
	wire _networkUnits_12_io_addressIn_ready;
	wire _networkUnits_12_io_peAddress_ready;
	wire _networkUnits_12_io_addressOut_valid;
	wire [63:0] _networkUnits_12_io_addressOut_bits;
	wire _networkUnits_11_io_addressIn_ready;
	wire _networkUnits_11_io_peAddress_ready;
	wire _networkUnits_11_io_addressOut_valid;
	wire [63:0] _networkUnits_11_io_addressOut_bits;
	wire _networkUnits_10_io_addressIn_ready;
	wire _networkUnits_10_io_peAddress_ready;
	wire _networkUnits_10_io_addressOut_valid;
	wire [63:0] _networkUnits_10_io_addressOut_bits;
	wire _networkUnits_9_io_addressIn_ready;
	wire _networkUnits_9_io_peAddress_ready;
	wire _networkUnits_9_io_addressOut_valid;
	wire [63:0] _networkUnits_9_io_addressOut_bits;
	wire _networkUnits_8_io_addressIn_ready;
	wire _networkUnits_8_io_peAddress_ready;
	wire _networkUnits_8_io_addressOut_valid;
	wire [63:0] _networkUnits_8_io_addressOut_bits;
	wire _networkUnits_7_io_addressIn_ready;
	wire _networkUnits_7_io_peAddress_ready;
	wire _networkUnits_7_io_addressOut_valid;
	wire [63:0] _networkUnits_7_io_addressOut_bits;
	wire _networkUnits_6_io_addressIn_ready;
	wire _networkUnits_6_io_peAddress_ready;
	wire _networkUnits_6_io_addressOut_valid;
	wire [63:0] _networkUnits_6_io_addressOut_bits;
	wire _networkUnits_5_io_addressIn_ready;
	wire _networkUnits_5_io_peAddress_ready;
	wire _networkUnits_5_io_addressOut_valid;
	wire [63:0] _networkUnits_5_io_addressOut_bits;
	wire _networkUnits_4_io_addressIn_ready;
	wire _networkUnits_4_io_peAddress_ready;
	wire _networkUnits_4_io_addressOut_valid;
	wire [63:0] _networkUnits_4_io_addressOut_bits;
	wire _networkUnits_3_io_addressIn_ready;
	wire _networkUnits_3_io_peAddress_ready;
	wire _networkUnits_3_io_addressOut_valid;
	wire [63:0] _networkUnits_3_io_addressOut_bits;
	wire _networkUnits_2_io_addressIn_ready;
	wire _networkUnits_2_io_peAddress_ready;
	wire _networkUnits_2_io_addressOut_valid;
	wire [63:0] _networkUnits_2_io_addressOut_bits;
	wire _networkUnits_1_io_addressIn_ready;
	wire _networkUnits_1_io_peAddress_ready;
	wire _networkUnits_1_io_addressOut_valid;
	wire [63:0] _networkUnits_1_io_addressOut_bits;
	wire _networkUnits_0_io_addressIn_ready;
	wire _networkUnits_0_io_peAddress_ready;
	wire _networkUnits_0_io_addressOut_valid;
	wire [63:0] _networkUnits_0_io_addressOut_bits;
	ArgumentNotifierNetworkUnit networkUnits_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_1_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_0_io_peAddress_ready),
		.io_peAddress_valid(_queues_0_io_addressOut_valid),
		.io_peAddress_bits(_queues_0_io_addressOut_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_15_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_0_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_2_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_1_io_peAddress_ready),
		.io_peAddress_valid(_queues_1_io_addressOut_valid),
		.io_peAddress_bits(_queues_1_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_0_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_1_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_1_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_3_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_2_io_peAddress_ready),
		.io_peAddress_valid(_queues_2_io_addressOut_valid),
		.io_peAddress_bits(_queues_2_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_1_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_2_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_2_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_4_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_3_io_peAddress_ready),
		.io_peAddress_valid(_queues_3_io_addressOut_valid),
		.io_peAddress_bits(_queues_3_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_2_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_3_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_3_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_5_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_4_io_peAddress_ready),
		.io_peAddress_valid(_queues_4_io_addressOut_valid),
		.io_peAddress_bits(_queues_4_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_3_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_4_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_4_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_6_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_5_io_peAddress_ready),
		.io_peAddress_valid(_queues_5_io_addressOut_valid),
		.io_peAddress_bits(_queues_5_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_4_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_5_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_5_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_7_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_6_io_peAddress_ready),
		.io_peAddress_valid(_queues_6_io_addressOut_valid),
		.io_peAddress_bits(_queues_6_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_5_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_6_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_6_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_8_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_7_io_peAddress_ready),
		.io_peAddress_valid(_queues_7_io_addressOut_valid),
		.io_peAddress_bits(_queues_7_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_6_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_7_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_7_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_9_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_8_io_peAddress_ready),
		.io_peAddress_valid(_queues_8_io_addressOut_valid),
		.io_peAddress_bits(_queues_8_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_7_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_8_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_8_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_10_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_9_io_peAddress_ready),
		.io_peAddress_valid(_queues_9_io_addressOut_valid),
		.io_peAddress_bits(_queues_9_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_8_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_9_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_9_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_11_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_10_io_peAddress_ready),
		.io_peAddress_valid(_queues_10_io_addressOut_valid),
		.io_peAddress_bits(_queues_10_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_9_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_10_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_10_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_12_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_11_io_peAddress_ready),
		.io_peAddress_valid(_queues_11_io_addressOut_valid),
		.io_peAddress_bits(_queues_11_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_10_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_11_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_11_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_13_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_12_io_peAddress_ready),
		.io_peAddress_valid(_queues_12_io_addressOut_valid),
		.io_peAddress_bits(_queues_12_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_11_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_12_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_12_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_14_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_13_io_peAddress_ready),
		.io_peAddress_valid(_queues_13_io_addressOut_valid),
		.io_peAddress_bits(_queues_13_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_12_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_13_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_13_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_15_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_14_io_peAddress_ready),
		.io_peAddress_valid(_queues_14_io_addressOut_valid),
		.io_peAddress_bits(_queues_14_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_13_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_14_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_14_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_16_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_15_io_peAddress_ready),
		.io_peAddress_valid(_queues_15_io_addressOut_valid),
		.io_peAddress_bits(_queues_15_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_14_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_15_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_15_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_17_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_16_io_peAddress_ready),
		.io_peAddress_valid(_queues_16_io_addressOut_valid),
		.io_peAddress_bits(_queues_16_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_15_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_16_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_16_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_18_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_17_io_peAddress_ready),
		.io_peAddress_valid(_queues_17_io_addressOut_valid),
		.io_peAddress_bits(_queues_17_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_16_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_17_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_17_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_19_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_18_io_peAddress_ready),
		.io_peAddress_valid(_queues_18_io_addressOut_valid),
		.io_peAddress_bits(_queues_18_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_17_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_18_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_18_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_20_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_19_io_peAddress_ready),
		.io_peAddress_valid(_queues_19_io_addressOut_valid),
		.io_peAddress_bits(_queues_19_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_18_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_19_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_19_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_21_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_20_io_peAddress_ready),
		.io_peAddress_valid(_queues_20_io_addressOut_valid),
		.io_peAddress_bits(_queues_20_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_19_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_20_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_20_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_22_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_21_io_peAddress_ready),
		.io_peAddress_valid(_queues_21_io_addressOut_valid),
		.io_peAddress_bits(_queues_21_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_20_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_21_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_21_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_23_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_22_io_peAddress_ready),
		.io_peAddress_valid(_queues_22_io_addressOut_valid),
		.io_peAddress_bits(_queues_22_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_21_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_22_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_22_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_24_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_23_io_peAddress_ready),
		.io_peAddress_valid(_queues_23_io_addressOut_valid),
		.io_peAddress_bits(_queues_23_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_22_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_23_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_23_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_25_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_24_io_peAddress_ready),
		.io_peAddress_valid(_queues_24_io_addressOut_valid),
		.io_peAddress_bits(_queues_24_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_23_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_24_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_24_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_26_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_25_io_peAddress_ready),
		.io_peAddress_valid(_queues_25_io_addressOut_valid),
		.io_peAddress_bits(_queues_25_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_24_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_25_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_25_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_27_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_26_io_peAddress_ready),
		.io_peAddress_valid(_queues_26_io_addressOut_valid),
		.io_peAddress_bits(_queues_26_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_25_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_26_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_26_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_28_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_27_io_peAddress_ready),
		.io_peAddress_valid(_queues_27_io_addressOut_valid),
		.io_peAddress_bits(_queues_27_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_26_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_27_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_27_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_29_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_28_io_peAddress_ready),
		.io_peAddress_valid(_queues_28_io_addressOut_valid),
		.io_peAddress_bits(_queues_28_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_27_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_28_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_28_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_30_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_29_io_peAddress_ready),
		.io_peAddress_valid(_queues_29_io_addressOut_valid),
		.io_peAddress_bits(_queues_29_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_28_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_29_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_29_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_31_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_30_io_peAddress_ready),
		.io_peAddress_valid(_queues_30_io_addressOut_valid),
		.io_peAddress_bits(_queues_30_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_29_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_30_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_30_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_32_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_31_io_peAddress_ready),
		.io_peAddress_valid(_queues_31_io_addressOut_valid),
		.io_peAddress_bits(_queues_31_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_30_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_31_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_31_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_33_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_32_io_peAddress_ready),
		.io_peAddress_valid(_queues_32_io_addressOut_valid),
		.io_peAddress_bits(_queues_32_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_31_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_32_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_32_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_34_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_33_io_peAddress_ready),
		.io_peAddress_valid(_queues_33_io_addressOut_valid),
		.io_peAddress_bits(_queues_33_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_32_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_33_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_33_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_35_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_34_io_peAddress_ready),
		.io_peAddress_valid(_queues_34_io_addressOut_valid),
		.io_peAddress_bits(_queues_34_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_33_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_34_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_34_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_36_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_35_io_peAddress_ready),
		.io_peAddress_valid(_queues_35_io_addressOut_valid),
		.io_peAddress_bits(_queues_35_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_34_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_35_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_35_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_37_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_36_io_peAddress_ready),
		.io_peAddress_valid(_queues_36_io_addressOut_valid),
		.io_peAddress_bits(_queues_36_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_35_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_36_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_36_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_38_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_37_io_peAddress_ready),
		.io_peAddress_valid(_queues_37_io_addressOut_valid),
		.io_peAddress_bits(_queues_37_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_36_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_37_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_37_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_39_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_38_io_peAddress_ready),
		.io_peAddress_valid(_queues_38_io_addressOut_valid),
		.io_peAddress_bits(_queues_38_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_37_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_38_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_38_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_40_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_39_io_peAddress_ready),
		.io_peAddress_valid(_queues_39_io_addressOut_valid),
		.io_peAddress_bits(_queues_39_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_38_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_39_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_39_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_41_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_40_io_peAddress_ready),
		.io_peAddress_valid(_queues_40_io_addressOut_valid),
		.io_peAddress_bits(_queues_40_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_39_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_40_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_40_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_42_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_41_io_peAddress_ready),
		.io_peAddress_valid(_queues_41_io_addressOut_valid),
		.io_peAddress_bits(_queues_41_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_40_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_41_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_41_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_43_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_42_io_peAddress_ready),
		.io_peAddress_valid(_queues_42_io_addressOut_valid),
		.io_peAddress_bits(_queues_42_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_41_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_42_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_42_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_44_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_43_io_peAddress_ready),
		.io_peAddress_valid(_queues_43_io_addressOut_valid),
		.io_peAddress_bits(_queues_43_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_42_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_43_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_43_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_45_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_44_io_peAddress_ready),
		.io_peAddress_valid(_queues_44_io_addressOut_valid),
		.io_peAddress_bits(_queues_44_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_43_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_44_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_44_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_46_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_45_io_peAddress_ready),
		.io_peAddress_valid(_queues_45_io_addressOut_valid),
		.io_peAddress_bits(_queues_45_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_44_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_45_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_45_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_47_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_46_io_peAddress_ready),
		.io_peAddress_valid(_queues_46_io_addressOut_valid),
		.io_peAddress_bits(_queues_46_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_45_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_46_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_46_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_48_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_47_io_peAddress_ready),
		.io_peAddress_valid(_queues_47_io_addressOut_valid),
		.io_peAddress_bits(_queues_47_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_46_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_47_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_47_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_49_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_48_io_peAddress_ready),
		.io_peAddress_valid(_queues_48_io_addressOut_valid),
		.io_peAddress_bits(_queues_48_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_47_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_48_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_48_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_50_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_49_io_peAddress_ready),
		.io_peAddress_valid(_queues_49_io_addressOut_valid),
		.io_peAddress_bits(_queues_49_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_48_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_49_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_49_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_51_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_50_io_peAddress_ready),
		.io_peAddress_valid(_queues_50_io_addressOut_valid),
		.io_peAddress_bits(_queues_50_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_49_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_50_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_50_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_52_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_51_io_peAddress_ready),
		.io_peAddress_valid(_queues_51_io_addressOut_valid),
		.io_peAddress_bits(_queues_51_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_50_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_51_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_51_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_53_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_52_io_peAddress_ready),
		.io_peAddress_valid(_queues_52_io_addressOut_valid),
		.io_peAddress_bits(_queues_52_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_51_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_52_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_52_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_54_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_53_io_peAddress_ready),
		.io_peAddress_valid(_queues_53_io_addressOut_valid),
		.io_peAddress_bits(_queues_53_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_52_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_53_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_53_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_55_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_54_io_peAddress_ready),
		.io_peAddress_valid(_queues_54_io_addressOut_valid),
		.io_peAddress_bits(_queues_54_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_53_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_54_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_54_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_56_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_55_io_peAddress_ready),
		.io_peAddress_valid(_queues_55_io_addressOut_valid),
		.io_peAddress_bits(_queues_55_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_54_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_55_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_55_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_57_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_56_io_peAddress_ready),
		.io_peAddress_valid(_queues_56_io_addressOut_valid),
		.io_peAddress_bits(_queues_56_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_55_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_56_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_56_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_58_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_57_io_peAddress_ready),
		.io_peAddress_valid(_queues_57_io_addressOut_valid),
		.io_peAddress_bits(_queues_57_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_56_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_57_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_57_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_59_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_58_io_peAddress_ready),
		.io_peAddress_valid(_queues_58_io_addressOut_valid),
		.io_peAddress_bits(_queues_58_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_57_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_58_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_58_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_60_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_59_io_peAddress_ready),
		.io_peAddress_valid(_queues_59_io_addressOut_valid),
		.io_peAddress_bits(_queues_59_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_58_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_59_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_59_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_61_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_60_io_peAddress_ready),
		.io_peAddress_valid(_queues_60_io_addressOut_valid),
		.io_peAddress_bits(_queues_60_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_59_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_60_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_60_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_62_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_61_io_peAddress_ready),
		.io_peAddress_valid(_queues_61_io_addressOut_valid),
		.io_peAddress_bits(_queues_61_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_60_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_61_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_61_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_63_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_63_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_62_io_peAddress_ready),
		.io_peAddress_valid(_queues_62_io_addressOut_valid),
		.io_peAddress_bits(_queues_62_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_61_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_62_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_62_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_64_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_64_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_63_io_peAddress_ready),
		.io_peAddress_valid(_queues_63_io_addressOut_valid),
		.io_peAddress_bits(_queues_63_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_62_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_63_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_63_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_64(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_64_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_65_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_65_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_64_io_peAddress_ready),
		.io_peAddress_valid(_queues_64_io_addressOut_valid),
		.io_peAddress_bits(_queues_64_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_63_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_64_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_64_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_65(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_65_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_66_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_66_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_65_io_peAddress_ready),
		.io_peAddress_valid(_queues_65_io_addressOut_valid),
		.io_peAddress_bits(_queues_65_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_64_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_65_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_65_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_66(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_66_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_67_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_67_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_66_io_peAddress_ready),
		.io_peAddress_valid(_queues_66_io_addressOut_valid),
		.io_peAddress_bits(_queues_66_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_65_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_66_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_66_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_67(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_67_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_68_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_68_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_67_io_peAddress_ready),
		.io_peAddress_valid(_queues_67_io_addressOut_valid),
		.io_peAddress_bits(_queues_67_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_66_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_67_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_67_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_68(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_68_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_69_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_69_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_68_io_peAddress_ready),
		.io_peAddress_valid(_queues_68_io_addressOut_valid),
		.io_peAddress_bits(_queues_68_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_67_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_68_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_68_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_69(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_69_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_70_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_70_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_69_io_peAddress_ready),
		.io_peAddress_valid(_queues_69_io_addressOut_valid),
		.io_peAddress_bits(_queues_69_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_68_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_69_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_69_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_70(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_70_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_71_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_71_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_70_io_peAddress_ready),
		.io_peAddress_valid(_queues_70_io_addressOut_valid),
		.io_peAddress_bits(_queues_70_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_69_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_70_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_70_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_71(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_71_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_72_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_72_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_71_io_peAddress_ready),
		.io_peAddress_valid(_queues_71_io_addressOut_valid),
		.io_peAddress_bits(_queues_71_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_70_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_71_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_71_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_72(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_72_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_73_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_73_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_72_io_peAddress_ready),
		.io_peAddress_valid(_queues_72_io_addressOut_valid),
		.io_peAddress_bits(_queues_72_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_71_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_72_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_72_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_73(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_73_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_74_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_74_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_73_io_peAddress_ready),
		.io_peAddress_valid(_queues_73_io_addressOut_valid),
		.io_peAddress_bits(_queues_73_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_72_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_73_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_73_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_74(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_74_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_75_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_75_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_74_io_peAddress_ready),
		.io_peAddress_valid(_queues_74_io_addressOut_valid),
		.io_peAddress_bits(_queues_74_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_73_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_74_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_74_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_75(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_75_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_76_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_76_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_75_io_peAddress_ready),
		.io_peAddress_valid(_queues_75_io_addressOut_valid),
		.io_peAddress_bits(_queues_75_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_74_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_75_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_75_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_76(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_76_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_77_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_77_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_76_io_peAddress_ready),
		.io_peAddress_valid(_queues_76_io_addressOut_valid),
		.io_peAddress_bits(_queues_76_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_75_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_76_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_76_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_77(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_77_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_78_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_78_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_77_io_peAddress_ready),
		.io_peAddress_valid(_queues_77_io_addressOut_valid),
		.io_peAddress_bits(_queues_77_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_76_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_77_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_77_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_78(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_networkUnits_78_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_79_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_79_io_addressOut_bits),
		.io_peAddress_ready(_networkUnits_78_io_peAddress_ready),
		.io_peAddress_valid(_queues_78_io_addressOut_valid),
		.io_peAddress_bits(_queues_78_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_77_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_78_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_78_io_addressOut_bits)
	);
	ArgumentNotifierNetworkUnit networkUnits_79(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(),
		.io_addressIn_valid(1'h0),
		.io_addressIn_bits(64'h0000000000000000),
		.io_peAddress_ready(_networkUnits_79_io_peAddress_ready),
		.io_peAddress_valid(_queues_79_io_addressOut_valid),
		.io_peAddress_bits(_queues_79_io_addressOut_bits),
		.io_addressOut_ready(_networkUnits_78_io_addressIn_ready),
		.io_addressOut_valid(_networkUnits_79_io_addressOut_valid),
		.io_addressOut_bits(_networkUnits_79_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit ArgumentNotifierServerNetworkUnit(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_0_ready),
		.io_vasAddressOut_valid(io_connVAS_0_valid),
		.io_vasAddressOut_bits(io_connVAS_0_bits)
	);
	ArgumentNotifierServerNetworkUnit_1 ArgumentNotifierServerNetworkUnit_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_1_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_1_ready),
		.io_vasAddressOut_valid(io_connVAS_1_valid),
		.io_vasAddressOut_bits(io_connVAS_1_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_1_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_2 ArgumentNotifierServerNetworkUnit_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_2_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_2_ready),
		.io_vasAddressOut_valid(io_connVAS_2_valid),
		.io_vasAddressOut_bits(io_connVAS_2_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_1_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_2_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_3 ArgumentNotifierServerNetworkUnit_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_3_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_3_ready),
		.io_vasAddressOut_valid(io_connVAS_3_valid),
		.io_vasAddressOut_bits(io_connVAS_3_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_2_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_3_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_4 ArgumentNotifierServerNetworkUnit_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_4_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_4_ready),
		.io_vasAddressOut_valid(io_connVAS_4_valid),
		.io_vasAddressOut_bits(io_connVAS_4_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_3_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_4_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_5 ArgumentNotifierServerNetworkUnit_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_5_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_5_ready),
		.io_vasAddressOut_valid(io_connVAS_5_valid),
		.io_vasAddressOut_bits(io_connVAS_5_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_4_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_5_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_6 ArgumentNotifierServerNetworkUnit_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_6_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_6_ready),
		.io_vasAddressOut_valid(io_connVAS_6_valid),
		.io_vasAddressOut_bits(io_connVAS_6_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_5_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_6_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_7 ArgumentNotifierServerNetworkUnit_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_7_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_7_ready),
		.io_vasAddressOut_valid(io_connVAS_7_valid),
		.io_vasAddressOut_bits(io_connVAS_7_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_6_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_7_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_8 ArgumentNotifierServerNetworkUnit_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_8_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_8_ready),
		.io_vasAddressOut_valid(io_connVAS_8_valid),
		.io_vasAddressOut_bits(io_connVAS_8_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_7_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_8_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_9 ArgumentNotifierServerNetworkUnit_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_9_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_9_ready),
		.io_vasAddressOut_valid(io_connVAS_9_valid),
		.io_vasAddressOut_bits(io_connVAS_9_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_8_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_9_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_10 ArgumentNotifierServerNetworkUnit_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_10_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_10_ready),
		.io_vasAddressOut_valid(io_connVAS_10_valid),
		.io_vasAddressOut_bits(io_connVAS_10_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_9_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_10_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_11 ArgumentNotifierServerNetworkUnit_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_11_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_11_ready),
		.io_vasAddressOut_valid(io_connVAS_11_valid),
		.io_vasAddressOut_bits(io_connVAS_11_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_10_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_11_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_12 ArgumentNotifierServerNetworkUnit_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_12_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_12_ready),
		.io_vasAddressOut_valid(io_connVAS_12_valid),
		.io_vasAddressOut_bits(io_connVAS_12_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_11_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_12_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_13 ArgumentNotifierServerNetworkUnit_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_13_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_13_ready),
		.io_vasAddressOut_valid(io_connVAS_13_valid),
		.io_vasAddressOut_bits(io_connVAS_13_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_12_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_13_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_14 ArgumentNotifierServerNetworkUnit_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_14_io_addressIn_ready),
		.io_addressIn_valid(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_valid),
		.io_addressIn_bits(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_14_ready),
		.io_vasAddressOut_valid(io_connVAS_14_valid),
		.io_vasAddressOut_bits(io_connVAS_14_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_13_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_14_io_addressOut_bits)
	);
	ArgumentNotifierServerNetworkUnit_15 ArgumentNotifierServerNetworkUnit_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(_ArgumentNotifierServerNetworkUnit_15_io_addressIn_ready),
		.io_addressIn_valid(_networkUnits_0_io_addressOut_valid),
		.io_addressIn_bits(_networkUnits_0_io_addressOut_bits),
		.io_vasAddressOut_ready(io_connVAS_15_ready),
		.io_vasAddressOut_valid(io_connVAS_15_valid),
		.io_vasAddressOut_bits(io_connVAS_15_bits),
		.io_addressOut_ready(_ArgumentNotifierServerNetworkUnit_14_io_addressIn_ready),
		.io_addressOut_valid(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_valid),
		.io_addressOut_bits(_ArgumentNotifierServerNetworkUnit_15_io_addressOut_bits)
	);
	AllocatorBuffer queues_0(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_0_ready),
		.io_addressIn_valid(io_connPE_0_valid),
		.io_addressIn_bits(io_connPE_0_bits),
		.io_addressOut_ready(_networkUnits_0_io_peAddress_ready),
		.io_addressOut_valid(_queues_0_io_addressOut_valid),
		.io_addressOut_bits(_queues_0_io_addressOut_bits)
	);
	AllocatorBuffer queues_1(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_1_ready),
		.io_addressIn_valid(io_connPE_1_valid),
		.io_addressIn_bits(io_connPE_1_bits),
		.io_addressOut_ready(_networkUnits_1_io_peAddress_ready),
		.io_addressOut_valid(_queues_1_io_addressOut_valid),
		.io_addressOut_bits(_queues_1_io_addressOut_bits)
	);
	AllocatorBuffer queues_2(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_2_ready),
		.io_addressIn_valid(io_connPE_2_valid),
		.io_addressIn_bits(io_connPE_2_bits),
		.io_addressOut_ready(_networkUnits_2_io_peAddress_ready),
		.io_addressOut_valid(_queues_2_io_addressOut_valid),
		.io_addressOut_bits(_queues_2_io_addressOut_bits)
	);
	AllocatorBuffer queues_3(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_3_ready),
		.io_addressIn_valid(io_connPE_3_valid),
		.io_addressIn_bits(io_connPE_3_bits),
		.io_addressOut_ready(_networkUnits_3_io_peAddress_ready),
		.io_addressOut_valid(_queues_3_io_addressOut_valid),
		.io_addressOut_bits(_queues_3_io_addressOut_bits)
	);
	AllocatorBuffer queues_4(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_4_ready),
		.io_addressIn_valid(io_connPE_4_valid),
		.io_addressIn_bits(io_connPE_4_bits),
		.io_addressOut_ready(_networkUnits_4_io_peAddress_ready),
		.io_addressOut_valid(_queues_4_io_addressOut_valid),
		.io_addressOut_bits(_queues_4_io_addressOut_bits)
	);
	AllocatorBuffer queues_5(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_5_ready),
		.io_addressIn_valid(io_connPE_5_valid),
		.io_addressIn_bits(io_connPE_5_bits),
		.io_addressOut_ready(_networkUnits_5_io_peAddress_ready),
		.io_addressOut_valid(_queues_5_io_addressOut_valid),
		.io_addressOut_bits(_queues_5_io_addressOut_bits)
	);
	AllocatorBuffer queues_6(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_6_ready),
		.io_addressIn_valid(io_connPE_6_valid),
		.io_addressIn_bits(io_connPE_6_bits),
		.io_addressOut_ready(_networkUnits_6_io_peAddress_ready),
		.io_addressOut_valid(_queues_6_io_addressOut_valid),
		.io_addressOut_bits(_queues_6_io_addressOut_bits)
	);
	AllocatorBuffer queues_7(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_7_ready),
		.io_addressIn_valid(io_connPE_7_valid),
		.io_addressIn_bits(io_connPE_7_bits),
		.io_addressOut_ready(_networkUnits_7_io_peAddress_ready),
		.io_addressOut_valid(_queues_7_io_addressOut_valid),
		.io_addressOut_bits(_queues_7_io_addressOut_bits)
	);
	AllocatorBuffer queues_8(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_8_ready),
		.io_addressIn_valid(io_connPE_8_valid),
		.io_addressIn_bits(io_connPE_8_bits),
		.io_addressOut_ready(_networkUnits_8_io_peAddress_ready),
		.io_addressOut_valid(_queues_8_io_addressOut_valid),
		.io_addressOut_bits(_queues_8_io_addressOut_bits)
	);
	AllocatorBuffer queues_9(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_9_ready),
		.io_addressIn_valid(io_connPE_9_valid),
		.io_addressIn_bits(io_connPE_9_bits),
		.io_addressOut_ready(_networkUnits_9_io_peAddress_ready),
		.io_addressOut_valid(_queues_9_io_addressOut_valid),
		.io_addressOut_bits(_queues_9_io_addressOut_bits)
	);
	AllocatorBuffer queues_10(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_10_ready),
		.io_addressIn_valid(io_connPE_10_valid),
		.io_addressIn_bits(io_connPE_10_bits),
		.io_addressOut_ready(_networkUnits_10_io_peAddress_ready),
		.io_addressOut_valid(_queues_10_io_addressOut_valid),
		.io_addressOut_bits(_queues_10_io_addressOut_bits)
	);
	AllocatorBuffer queues_11(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_11_ready),
		.io_addressIn_valid(io_connPE_11_valid),
		.io_addressIn_bits(io_connPE_11_bits),
		.io_addressOut_ready(_networkUnits_11_io_peAddress_ready),
		.io_addressOut_valid(_queues_11_io_addressOut_valid),
		.io_addressOut_bits(_queues_11_io_addressOut_bits)
	);
	AllocatorBuffer queues_12(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_12_ready),
		.io_addressIn_valid(io_connPE_12_valid),
		.io_addressIn_bits(io_connPE_12_bits),
		.io_addressOut_ready(_networkUnits_12_io_peAddress_ready),
		.io_addressOut_valid(_queues_12_io_addressOut_valid),
		.io_addressOut_bits(_queues_12_io_addressOut_bits)
	);
	AllocatorBuffer queues_13(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_13_ready),
		.io_addressIn_valid(io_connPE_13_valid),
		.io_addressIn_bits(io_connPE_13_bits),
		.io_addressOut_ready(_networkUnits_13_io_peAddress_ready),
		.io_addressOut_valid(_queues_13_io_addressOut_valid),
		.io_addressOut_bits(_queues_13_io_addressOut_bits)
	);
	AllocatorBuffer queues_14(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_14_ready),
		.io_addressIn_valid(io_connPE_14_valid),
		.io_addressIn_bits(io_connPE_14_bits),
		.io_addressOut_ready(_networkUnits_14_io_peAddress_ready),
		.io_addressOut_valid(_queues_14_io_addressOut_valid),
		.io_addressOut_bits(_queues_14_io_addressOut_bits)
	);
	AllocatorBuffer queues_15(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_15_ready),
		.io_addressIn_valid(io_connPE_15_valid),
		.io_addressIn_bits(io_connPE_15_bits),
		.io_addressOut_ready(_networkUnits_15_io_peAddress_ready),
		.io_addressOut_valid(_queues_15_io_addressOut_valid),
		.io_addressOut_bits(_queues_15_io_addressOut_bits)
	);
	AllocatorBuffer queues_16(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_16_ready),
		.io_addressIn_valid(io_connPE_16_valid),
		.io_addressIn_bits(io_connPE_16_bits),
		.io_addressOut_ready(_networkUnits_16_io_peAddress_ready),
		.io_addressOut_valid(_queues_16_io_addressOut_valid),
		.io_addressOut_bits(_queues_16_io_addressOut_bits)
	);
	AllocatorBuffer queues_17(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_17_ready),
		.io_addressIn_valid(io_connPE_17_valid),
		.io_addressIn_bits(io_connPE_17_bits),
		.io_addressOut_ready(_networkUnits_17_io_peAddress_ready),
		.io_addressOut_valid(_queues_17_io_addressOut_valid),
		.io_addressOut_bits(_queues_17_io_addressOut_bits)
	);
	AllocatorBuffer queues_18(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_18_ready),
		.io_addressIn_valid(io_connPE_18_valid),
		.io_addressIn_bits(io_connPE_18_bits),
		.io_addressOut_ready(_networkUnits_18_io_peAddress_ready),
		.io_addressOut_valid(_queues_18_io_addressOut_valid),
		.io_addressOut_bits(_queues_18_io_addressOut_bits)
	);
	AllocatorBuffer queues_19(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_19_ready),
		.io_addressIn_valid(io_connPE_19_valid),
		.io_addressIn_bits(io_connPE_19_bits),
		.io_addressOut_ready(_networkUnits_19_io_peAddress_ready),
		.io_addressOut_valid(_queues_19_io_addressOut_valid),
		.io_addressOut_bits(_queues_19_io_addressOut_bits)
	);
	AllocatorBuffer queues_20(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_20_ready),
		.io_addressIn_valid(io_connPE_20_valid),
		.io_addressIn_bits(io_connPE_20_bits),
		.io_addressOut_ready(_networkUnits_20_io_peAddress_ready),
		.io_addressOut_valid(_queues_20_io_addressOut_valid),
		.io_addressOut_bits(_queues_20_io_addressOut_bits)
	);
	AllocatorBuffer queues_21(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_21_ready),
		.io_addressIn_valid(io_connPE_21_valid),
		.io_addressIn_bits(io_connPE_21_bits),
		.io_addressOut_ready(_networkUnits_21_io_peAddress_ready),
		.io_addressOut_valid(_queues_21_io_addressOut_valid),
		.io_addressOut_bits(_queues_21_io_addressOut_bits)
	);
	AllocatorBuffer queues_22(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_22_ready),
		.io_addressIn_valid(io_connPE_22_valid),
		.io_addressIn_bits(io_connPE_22_bits),
		.io_addressOut_ready(_networkUnits_22_io_peAddress_ready),
		.io_addressOut_valid(_queues_22_io_addressOut_valid),
		.io_addressOut_bits(_queues_22_io_addressOut_bits)
	);
	AllocatorBuffer queues_23(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_23_ready),
		.io_addressIn_valid(io_connPE_23_valid),
		.io_addressIn_bits(io_connPE_23_bits),
		.io_addressOut_ready(_networkUnits_23_io_peAddress_ready),
		.io_addressOut_valid(_queues_23_io_addressOut_valid),
		.io_addressOut_bits(_queues_23_io_addressOut_bits)
	);
	AllocatorBuffer queues_24(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_24_ready),
		.io_addressIn_valid(io_connPE_24_valid),
		.io_addressIn_bits(io_connPE_24_bits),
		.io_addressOut_ready(_networkUnits_24_io_peAddress_ready),
		.io_addressOut_valid(_queues_24_io_addressOut_valid),
		.io_addressOut_bits(_queues_24_io_addressOut_bits)
	);
	AllocatorBuffer queues_25(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_25_ready),
		.io_addressIn_valid(io_connPE_25_valid),
		.io_addressIn_bits(io_connPE_25_bits),
		.io_addressOut_ready(_networkUnits_25_io_peAddress_ready),
		.io_addressOut_valid(_queues_25_io_addressOut_valid),
		.io_addressOut_bits(_queues_25_io_addressOut_bits)
	);
	AllocatorBuffer queues_26(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_26_ready),
		.io_addressIn_valid(io_connPE_26_valid),
		.io_addressIn_bits(io_connPE_26_bits),
		.io_addressOut_ready(_networkUnits_26_io_peAddress_ready),
		.io_addressOut_valid(_queues_26_io_addressOut_valid),
		.io_addressOut_bits(_queues_26_io_addressOut_bits)
	);
	AllocatorBuffer queues_27(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_27_ready),
		.io_addressIn_valid(io_connPE_27_valid),
		.io_addressIn_bits(io_connPE_27_bits),
		.io_addressOut_ready(_networkUnits_27_io_peAddress_ready),
		.io_addressOut_valid(_queues_27_io_addressOut_valid),
		.io_addressOut_bits(_queues_27_io_addressOut_bits)
	);
	AllocatorBuffer queues_28(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_28_ready),
		.io_addressIn_valid(io_connPE_28_valid),
		.io_addressIn_bits(io_connPE_28_bits),
		.io_addressOut_ready(_networkUnits_28_io_peAddress_ready),
		.io_addressOut_valid(_queues_28_io_addressOut_valid),
		.io_addressOut_bits(_queues_28_io_addressOut_bits)
	);
	AllocatorBuffer queues_29(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_29_ready),
		.io_addressIn_valid(io_connPE_29_valid),
		.io_addressIn_bits(io_connPE_29_bits),
		.io_addressOut_ready(_networkUnits_29_io_peAddress_ready),
		.io_addressOut_valid(_queues_29_io_addressOut_valid),
		.io_addressOut_bits(_queues_29_io_addressOut_bits)
	);
	AllocatorBuffer queues_30(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_30_ready),
		.io_addressIn_valid(io_connPE_30_valid),
		.io_addressIn_bits(io_connPE_30_bits),
		.io_addressOut_ready(_networkUnits_30_io_peAddress_ready),
		.io_addressOut_valid(_queues_30_io_addressOut_valid),
		.io_addressOut_bits(_queues_30_io_addressOut_bits)
	);
	AllocatorBuffer queues_31(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_31_ready),
		.io_addressIn_valid(io_connPE_31_valid),
		.io_addressIn_bits(io_connPE_31_bits),
		.io_addressOut_ready(_networkUnits_31_io_peAddress_ready),
		.io_addressOut_valid(_queues_31_io_addressOut_valid),
		.io_addressOut_bits(_queues_31_io_addressOut_bits)
	);
	AllocatorBuffer queues_32(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_32_ready),
		.io_addressIn_valid(io_connPE_32_valid),
		.io_addressIn_bits(io_connPE_32_bits),
		.io_addressOut_ready(_networkUnits_32_io_peAddress_ready),
		.io_addressOut_valid(_queues_32_io_addressOut_valid),
		.io_addressOut_bits(_queues_32_io_addressOut_bits)
	);
	AllocatorBuffer queues_33(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_33_ready),
		.io_addressIn_valid(io_connPE_33_valid),
		.io_addressIn_bits(io_connPE_33_bits),
		.io_addressOut_ready(_networkUnits_33_io_peAddress_ready),
		.io_addressOut_valid(_queues_33_io_addressOut_valid),
		.io_addressOut_bits(_queues_33_io_addressOut_bits)
	);
	AllocatorBuffer queues_34(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_34_ready),
		.io_addressIn_valid(io_connPE_34_valid),
		.io_addressIn_bits(io_connPE_34_bits),
		.io_addressOut_ready(_networkUnits_34_io_peAddress_ready),
		.io_addressOut_valid(_queues_34_io_addressOut_valid),
		.io_addressOut_bits(_queues_34_io_addressOut_bits)
	);
	AllocatorBuffer queues_35(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_35_ready),
		.io_addressIn_valid(io_connPE_35_valid),
		.io_addressIn_bits(io_connPE_35_bits),
		.io_addressOut_ready(_networkUnits_35_io_peAddress_ready),
		.io_addressOut_valid(_queues_35_io_addressOut_valid),
		.io_addressOut_bits(_queues_35_io_addressOut_bits)
	);
	AllocatorBuffer queues_36(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_36_ready),
		.io_addressIn_valid(io_connPE_36_valid),
		.io_addressIn_bits(io_connPE_36_bits),
		.io_addressOut_ready(_networkUnits_36_io_peAddress_ready),
		.io_addressOut_valid(_queues_36_io_addressOut_valid),
		.io_addressOut_bits(_queues_36_io_addressOut_bits)
	);
	AllocatorBuffer queues_37(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_37_ready),
		.io_addressIn_valid(io_connPE_37_valid),
		.io_addressIn_bits(io_connPE_37_bits),
		.io_addressOut_ready(_networkUnits_37_io_peAddress_ready),
		.io_addressOut_valid(_queues_37_io_addressOut_valid),
		.io_addressOut_bits(_queues_37_io_addressOut_bits)
	);
	AllocatorBuffer queues_38(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_38_ready),
		.io_addressIn_valid(io_connPE_38_valid),
		.io_addressIn_bits(io_connPE_38_bits),
		.io_addressOut_ready(_networkUnits_38_io_peAddress_ready),
		.io_addressOut_valid(_queues_38_io_addressOut_valid),
		.io_addressOut_bits(_queues_38_io_addressOut_bits)
	);
	AllocatorBuffer queues_39(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_39_ready),
		.io_addressIn_valid(io_connPE_39_valid),
		.io_addressIn_bits(io_connPE_39_bits),
		.io_addressOut_ready(_networkUnits_39_io_peAddress_ready),
		.io_addressOut_valid(_queues_39_io_addressOut_valid),
		.io_addressOut_bits(_queues_39_io_addressOut_bits)
	);
	AllocatorBuffer queues_40(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_40_ready),
		.io_addressIn_valid(io_connPE_40_valid),
		.io_addressIn_bits(io_connPE_40_bits),
		.io_addressOut_ready(_networkUnits_40_io_peAddress_ready),
		.io_addressOut_valid(_queues_40_io_addressOut_valid),
		.io_addressOut_bits(_queues_40_io_addressOut_bits)
	);
	AllocatorBuffer queues_41(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_41_ready),
		.io_addressIn_valid(io_connPE_41_valid),
		.io_addressIn_bits(io_connPE_41_bits),
		.io_addressOut_ready(_networkUnits_41_io_peAddress_ready),
		.io_addressOut_valid(_queues_41_io_addressOut_valid),
		.io_addressOut_bits(_queues_41_io_addressOut_bits)
	);
	AllocatorBuffer queues_42(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_42_ready),
		.io_addressIn_valid(io_connPE_42_valid),
		.io_addressIn_bits(io_connPE_42_bits),
		.io_addressOut_ready(_networkUnits_42_io_peAddress_ready),
		.io_addressOut_valid(_queues_42_io_addressOut_valid),
		.io_addressOut_bits(_queues_42_io_addressOut_bits)
	);
	AllocatorBuffer queues_43(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_43_ready),
		.io_addressIn_valid(io_connPE_43_valid),
		.io_addressIn_bits(io_connPE_43_bits),
		.io_addressOut_ready(_networkUnits_43_io_peAddress_ready),
		.io_addressOut_valid(_queues_43_io_addressOut_valid),
		.io_addressOut_bits(_queues_43_io_addressOut_bits)
	);
	AllocatorBuffer queues_44(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_44_ready),
		.io_addressIn_valid(io_connPE_44_valid),
		.io_addressIn_bits(io_connPE_44_bits),
		.io_addressOut_ready(_networkUnits_44_io_peAddress_ready),
		.io_addressOut_valid(_queues_44_io_addressOut_valid),
		.io_addressOut_bits(_queues_44_io_addressOut_bits)
	);
	AllocatorBuffer queues_45(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_45_ready),
		.io_addressIn_valid(io_connPE_45_valid),
		.io_addressIn_bits(io_connPE_45_bits),
		.io_addressOut_ready(_networkUnits_45_io_peAddress_ready),
		.io_addressOut_valid(_queues_45_io_addressOut_valid),
		.io_addressOut_bits(_queues_45_io_addressOut_bits)
	);
	AllocatorBuffer queues_46(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_46_ready),
		.io_addressIn_valid(io_connPE_46_valid),
		.io_addressIn_bits(io_connPE_46_bits),
		.io_addressOut_ready(_networkUnits_46_io_peAddress_ready),
		.io_addressOut_valid(_queues_46_io_addressOut_valid),
		.io_addressOut_bits(_queues_46_io_addressOut_bits)
	);
	AllocatorBuffer queues_47(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_47_ready),
		.io_addressIn_valid(io_connPE_47_valid),
		.io_addressIn_bits(io_connPE_47_bits),
		.io_addressOut_ready(_networkUnits_47_io_peAddress_ready),
		.io_addressOut_valid(_queues_47_io_addressOut_valid),
		.io_addressOut_bits(_queues_47_io_addressOut_bits)
	);
	AllocatorBuffer queues_48(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_48_ready),
		.io_addressIn_valid(io_connPE_48_valid),
		.io_addressIn_bits(io_connPE_48_bits),
		.io_addressOut_ready(_networkUnits_48_io_peAddress_ready),
		.io_addressOut_valid(_queues_48_io_addressOut_valid),
		.io_addressOut_bits(_queues_48_io_addressOut_bits)
	);
	AllocatorBuffer queues_49(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_49_ready),
		.io_addressIn_valid(io_connPE_49_valid),
		.io_addressIn_bits(io_connPE_49_bits),
		.io_addressOut_ready(_networkUnits_49_io_peAddress_ready),
		.io_addressOut_valid(_queues_49_io_addressOut_valid),
		.io_addressOut_bits(_queues_49_io_addressOut_bits)
	);
	AllocatorBuffer queues_50(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_50_ready),
		.io_addressIn_valid(io_connPE_50_valid),
		.io_addressIn_bits(io_connPE_50_bits),
		.io_addressOut_ready(_networkUnits_50_io_peAddress_ready),
		.io_addressOut_valid(_queues_50_io_addressOut_valid),
		.io_addressOut_bits(_queues_50_io_addressOut_bits)
	);
	AllocatorBuffer queues_51(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_51_ready),
		.io_addressIn_valid(io_connPE_51_valid),
		.io_addressIn_bits(io_connPE_51_bits),
		.io_addressOut_ready(_networkUnits_51_io_peAddress_ready),
		.io_addressOut_valid(_queues_51_io_addressOut_valid),
		.io_addressOut_bits(_queues_51_io_addressOut_bits)
	);
	AllocatorBuffer queues_52(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_52_ready),
		.io_addressIn_valid(io_connPE_52_valid),
		.io_addressIn_bits(io_connPE_52_bits),
		.io_addressOut_ready(_networkUnits_52_io_peAddress_ready),
		.io_addressOut_valid(_queues_52_io_addressOut_valid),
		.io_addressOut_bits(_queues_52_io_addressOut_bits)
	);
	AllocatorBuffer queues_53(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_53_ready),
		.io_addressIn_valid(io_connPE_53_valid),
		.io_addressIn_bits(io_connPE_53_bits),
		.io_addressOut_ready(_networkUnits_53_io_peAddress_ready),
		.io_addressOut_valid(_queues_53_io_addressOut_valid),
		.io_addressOut_bits(_queues_53_io_addressOut_bits)
	);
	AllocatorBuffer queues_54(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_54_ready),
		.io_addressIn_valid(io_connPE_54_valid),
		.io_addressIn_bits(io_connPE_54_bits),
		.io_addressOut_ready(_networkUnits_54_io_peAddress_ready),
		.io_addressOut_valid(_queues_54_io_addressOut_valid),
		.io_addressOut_bits(_queues_54_io_addressOut_bits)
	);
	AllocatorBuffer queues_55(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_55_ready),
		.io_addressIn_valid(io_connPE_55_valid),
		.io_addressIn_bits(io_connPE_55_bits),
		.io_addressOut_ready(_networkUnits_55_io_peAddress_ready),
		.io_addressOut_valid(_queues_55_io_addressOut_valid),
		.io_addressOut_bits(_queues_55_io_addressOut_bits)
	);
	AllocatorBuffer queues_56(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_56_ready),
		.io_addressIn_valid(io_connPE_56_valid),
		.io_addressIn_bits(io_connPE_56_bits),
		.io_addressOut_ready(_networkUnits_56_io_peAddress_ready),
		.io_addressOut_valid(_queues_56_io_addressOut_valid),
		.io_addressOut_bits(_queues_56_io_addressOut_bits)
	);
	AllocatorBuffer queues_57(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_57_ready),
		.io_addressIn_valid(io_connPE_57_valid),
		.io_addressIn_bits(io_connPE_57_bits),
		.io_addressOut_ready(_networkUnits_57_io_peAddress_ready),
		.io_addressOut_valid(_queues_57_io_addressOut_valid),
		.io_addressOut_bits(_queues_57_io_addressOut_bits)
	);
	AllocatorBuffer queues_58(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_58_ready),
		.io_addressIn_valid(io_connPE_58_valid),
		.io_addressIn_bits(io_connPE_58_bits),
		.io_addressOut_ready(_networkUnits_58_io_peAddress_ready),
		.io_addressOut_valid(_queues_58_io_addressOut_valid),
		.io_addressOut_bits(_queues_58_io_addressOut_bits)
	);
	AllocatorBuffer queues_59(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_59_ready),
		.io_addressIn_valid(io_connPE_59_valid),
		.io_addressIn_bits(io_connPE_59_bits),
		.io_addressOut_ready(_networkUnits_59_io_peAddress_ready),
		.io_addressOut_valid(_queues_59_io_addressOut_valid),
		.io_addressOut_bits(_queues_59_io_addressOut_bits)
	);
	AllocatorBuffer queues_60(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_60_ready),
		.io_addressIn_valid(io_connPE_60_valid),
		.io_addressIn_bits(io_connPE_60_bits),
		.io_addressOut_ready(_networkUnits_60_io_peAddress_ready),
		.io_addressOut_valid(_queues_60_io_addressOut_valid),
		.io_addressOut_bits(_queues_60_io_addressOut_bits)
	);
	AllocatorBuffer queues_61(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_61_ready),
		.io_addressIn_valid(io_connPE_61_valid),
		.io_addressIn_bits(io_connPE_61_bits),
		.io_addressOut_ready(_networkUnits_61_io_peAddress_ready),
		.io_addressOut_valid(_queues_61_io_addressOut_valid),
		.io_addressOut_bits(_queues_61_io_addressOut_bits)
	);
	AllocatorBuffer queues_62(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_62_ready),
		.io_addressIn_valid(io_connPE_62_valid),
		.io_addressIn_bits(io_connPE_62_bits),
		.io_addressOut_ready(_networkUnits_62_io_peAddress_ready),
		.io_addressOut_valid(_queues_62_io_addressOut_valid),
		.io_addressOut_bits(_queues_62_io_addressOut_bits)
	);
	AllocatorBuffer queues_63(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_63_ready),
		.io_addressIn_valid(io_connPE_63_valid),
		.io_addressIn_bits(io_connPE_63_bits),
		.io_addressOut_ready(_networkUnits_63_io_peAddress_ready),
		.io_addressOut_valid(_queues_63_io_addressOut_valid),
		.io_addressOut_bits(_queues_63_io_addressOut_bits)
	);
	AllocatorBuffer queues_64(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_64_ready),
		.io_addressIn_valid(io_connPE_64_valid),
		.io_addressIn_bits(io_connPE_64_bits),
		.io_addressOut_ready(_networkUnits_64_io_peAddress_ready),
		.io_addressOut_valid(_queues_64_io_addressOut_valid),
		.io_addressOut_bits(_queues_64_io_addressOut_bits)
	);
	AllocatorBuffer queues_65(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_65_ready),
		.io_addressIn_valid(io_connPE_65_valid),
		.io_addressIn_bits(io_connPE_65_bits),
		.io_addressOut_ready(_networkUnits_65_io_peAddress_ready),
		.io_addressOut_valid(_queues_65_io_addressOut_valid),
		.io_addressOut_bits(_queues_65_io_addressOut_bits)
	);
	AllocatorBuffer queues_66(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_66_ready),
		.io_addressIn_valid(io_connPE_66_valid),
		.io_addressIn_bits(io_connPE_66_bits),
		.io_addressOut_ready(_networkUnits_66_io_peAddress_ready),
		.io_addressOut_valid(_queues_66_io_addressOut_valid),
		.io_addressOut_bits(_queues_66_io_addressOut_bits)
	);
	AllocatorBuffer queues_67(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_67_ready),
		.io_addressIn_valid(io_connPE_67_valid),
		.io_addressIn_bits(io_connPE_67_bits),
		.io_addressOut_ready(_networkUnits_67_io_peAddress_ready),
		.io_addressOut_valid(_queues_67_io_addressOut_valid),
		.io_addressOut_bits(_queues_67_io_addressOut_bits)
	);
	AllocatorBuffer queues_68(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_68_ready),
		.io_addressIn_valid(io_connPE_68_valid),
		.io_addressIn_bits(io_connPE_68_bits),
		.io_addressOut_ready(_networkUnits_68_io_peAddress_ready),
		.io_addressOut_valid(_queues_68_io_addressOut_valid),
		.io_addressOut_bits(_queues_68_io_addressOut_bits)
	);
	AllocatorBuffer queues_69(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_69_ready),
		.io_addressIn_valid(io_connPE_69_valid),
		.io_addressIn_bits(io_connPE_69_bits),
		.io_addressOut_ready(_networkUnits_69_io_peAddress_ready),
		.io_addressOut_valid(_queues_69_io_addressOut_valid),
		.io_addressOut_bits(_queues_69_io_addressOut_bits)
	);
	AllocatorBuffer queues_70(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_70_ready),
		.io_addressIn_valid(io_connPE_70_valid),
		.io_addressIn_bits(io_connPE_70_bits),
		.io_addressOut_ready(_networkUnits_70_io_peAddress_ready),
		.io_addressOut_valid(_queues_70_io_addressOut_valid),
		.io_addressOut_bits(_queues_70_io_addressOut_bits)
	);
	AllocatorBuffer queues_71(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_71_ready),
		.io_addressIn_valid(io_connPE_71_valid),
		.io_addressIn_bits(io_connPE_71_bits),
		.io_addressOut_ready(_networkUnits_71_io_peAddress_ready),
		.io_addressOut_valid(_queues_71_io_addressOut_valid),
		.io_addressOut_bits(_queues_71_io_addressOut_bits)
	);
	AllocatorBuffer queues_72(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_72_ready),
		.io_addressIn_valid(io_connPE_72_valid),
		.io_addressIn_bits(io_connPE_72_bits),
		.io_addressOut_ready(_networkUnits_72_io_peAddress_ready),
		.io_addressOut_valid(_queues_72_io_addressOut_valid),
		.io_addressOut_bits(_queues_72_io_addressOut_bits)
	);
	AllocatorBuffer queues_73(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_73_ready),
		.io_addressIn_valid(io_connPE_73_valid),
		.io_addressIn_bits(io_connPE_73_bits),
		.io_addressOut_ready(_networkUnits_73_io_peAddress_ready),
		.io_addressOut_valid(_queues_73_io_addressOut_valid),
		.io_addressOut_bits(_queues_73_io_addressOut_bits)
	);
	AllocatorBuffer queues_74(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_74_ready),
		.io_addressIn_valid(io_connPE_74_valid),
		.io_addressIn_bits(io_connPE_74_bits),
		.io_addressOut_ready(_networkUnits_74_io_peAddress_ready),
		.io_addressOut_valid(_queues_74_io_addressOut_valid),
		.io_addressOut_bits(_queues_74_io_addressOut_bits)
	);
	AllocatorBuffer queues_75(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_75_ready),
		.io_addressIn_valid(io_connPE_75_valid),
		.io_addressIn_bits(io_connPE_75_bits),
		.io_addressOut_ready(_networkUnits_75_io_peAddress_ready),
		.io_addressOut_valid(_queues_75_io_addressOut_valid),
		.io_addressOut_bits(_queues_75_io_addressOut_bits)
	);
	AllocatorBuffer queues_76(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_76_ready),
		.io_addressIn_valid(io_connPE_76_valid),
		.io_addressIn_bits(io_connPE_76_bits),
		.io_addressOut_ready(_networkUnits_76_io_peAddress_ready),
		.io_addressOut_valid(_queues_76_io_addressOut_valid),
		.io_addressOut_bits(_queues_76_io_addressOut_bits)
	);
	AllocatorBuffer queues_77(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_77_ready),
		.io_addressIn_valid(io_connPE_77_valid),
		.io_addressIn_bits(io_connPE_77_bits),
		.io_addressOut_ready(_networkUnits_77_io_peAddress_ready),
		.io_addressOut_valid(_queues_77_io_addressOut_valid),
		.io_addressOut_bits(_queues_77_io_addressOut_bits)
	);
	AllocatorBuffer queues_78(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_78_ready),
		.io_addressIn_valid(io_connPE_78_valid),
		.io_addressIn_bits(io_connPE_78_bits),
		.io_addressOut_ready(_networkUnits_78_io_peAddress_ready),
		.io_addressOut_valid(_queues_78_io_addressOut_valid),
		.io_addressOut_bits(_queues_78_io_addressOut_bits)
	);
	AllocatorBuffer queues_79(
		.clock(clock),
		.reset(reset),
		.io_addressIn_ready(io_connPE_79_ready),
		.io_addressIn_valid(io_connPE_79_valid),
		.io_addressIn_bits(io_connPE_79_bits),
		.io_addressOut_ready(_networkUnits_79_io_peAddress_ready),
		.io_addressOut_valid(_queues_79_io_addressOut_valid),
		.io_addressOut_bits(_queues_79_io_addressOut_bits)
	);
endmodule
module ram_16x64 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [3:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [63:0] R0_data;
	input [3:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [63:0] W0_data;
	reg [63:0] Memory [0:15];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue16_UInt (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits;
	reg [3:0] enq_ptr_value;
	reg [3:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 4'h0;
			deq_ptr_value <= 4'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 4'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 4'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_16x64 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module ram_16x128 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [3:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [127:0] R0_data;
	input [3:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [127:0] W0_data;
	reg [127:0] Memory [0:15];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (R0_en ? Memory[R0_addr] : 128'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue16_UInt_2 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [127:0] io_enq_bits;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [127:0] io_deq_bits;
	reg [3:0] enq_ptr_value;
	reg [3:0] deq_ptr_value;
	reg maybe_full;
	wire ptr_match = enq_ptr_value == deq_ptr_value;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	always @(posedge clock)
		if (reset) begin
			enq_ptr_value <= 4'h0;
			deq_ptr_value <= 4'h0;
			maybe_full <= 1'h0;
		end
		else begin : sv2v_autoblock_1
			reg do_deq;
			do_deq = io_deq_ready & ~empty;
			if (do_enq)
				enq_ptr_value <= enq_ptr_value + 4'h1;
			if (do_deq)
				deq_ptr_value <= deq_ptr_value + 4'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	ram_16x128 ram_ext(
		.R0_addr(deq_ptr_value),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits),
		.W0_addr(enq_ptr_value),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module ArgumentServer (
	clock,
	reset,
	io_connNetwork_ready,
	io_connNetwork_valid,
	io_connNetwork_bits,
	io_connStealNtw_ctrl_serveStealReq_valid,
	io_connStealNtw_ctrl_serveStealReq_ready,
	io_connStealNtw_data_qOutTask_ready,
	io_connStealNtw_data_qOutTask_valid,
	io_connStealNtw_data_qOutTask_bits,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	io_read_address_task_ready,
	io_read_address_task_valid,
	io_read_address_task_bits,
	io_read_data_task_ready,
	io_read_data_task_valid,
	io_read_data_task_bits
);
	input clock;
	input reset;
	output wire io_connNetwork_ready;
	input io_connNetwork_valid;
	input [63:0] io_connNetwork_bits;
	output wire io_connStealNtw_ctrl_serveStealReq_valid;
	input io_connStealNtw_ctrl_serveStealReq_ready;
	input io_connStealNtw_data_qOutTask_ready;
	output wire io_connStealNtw_data_qOutTask_valid;
	output wire [127:0] io_connStealNtw_data_qOutTask_bits;
	input io_read_address_ready;
	output wire io_read_address_valid;
	output wire [63:0] io_read_address_bits;
	output wire io_read_data_ready;
	input io_read_data_valid;
	input [31:0] io_read_data_bits;
	input io_write_address_ready;
	output wire io_write_address_valid;
	output wire [63:0] io_write_address_bits;
	input io_write_data_ready;
	output wire io_write_data_valid;
	output wire [31:0] io_write_data_bits;
	input io_read_address_task_ready;
	output wire io_read_address_task_valid;
	output wire [63:0] io_read_address_task_bits;
	output wire io_read_data_task_ready;
	input io_read_data_task_valid;
	input [31:0] io_read_data_task_bits;
	wire _readyTasksQueue_io_enq_ready;
	wire _readyTasksQueue_io_deq_valid;
	wire [127:0] _readyTasksQueue_io_deq_bits;
	wire _addressesOfReadyTasks_io_enq_ready;
	wire _addressesOfReadyTasks_io_deq_valid;
	wire [63:0] _addressesOfReadyTasks_io_deq_bits;
	wire _addrNtwInQueue_io_deq_valid;
	wire [63:0] _addrNtwInQueue_io_deq_bits;
	reg [3:0] counterStateReg;
	reg [63:0] counterReg;
	reg [63:0] currReadAddr;
	reg [63:0] counterAddr;
	reg [63:0] addrMask;
	reg helpGarbageCollector;
	wire _GEN = counterStateReg == 4'h1;
	wire _GEN_0 = counterStateReg == 4'h2;
	wire _GEN_1 = counterStateReg == 4'h3;
	wire _GEN_2 = _GEN | _GEN_0;
	wire _GEN_3 = counterStateReg == 4'h4;
	wire _GEN_4 = counterStateReg == 4'h5;
	wire _GEN_5 = counterStateReg == 4'h7;
	wire _GEN_6 = ((_GEN | _GEN_0) | _GEN_1) | _GEN_3;
	reg [3:0] taskReadAddressStateReg;
	reg [63:0] taskAddr;
	wire _GEN_7 = taskReadAddressStateReg == 4'h6;
	wire _GEN_8 = taskReadAddressStateReg == 4'h8;
	reg [3:0] taskReadStateReg;
	reg [1:0] taskReadCount;
	reg [31:0] taskRegisters_0;
	reg [31:0] taskRegisters_1;
	reg [31:0] taskRegisters_2;
	reg [31:0] taskRegisters_3;
	wire io_read_data_task_ready_0 = taskReadStateReg == 4'h9;
	wire _GEN_9 = taskReadStateReg == 4'ha;
	reg [31:0] tasksGivenAwayCount;
	reg [127:0] taskReg;
	reg [3:0] taskWriteStateReg;
	wire _GEN_10 = taskWriteStateReg == 4'hb;
	wire _GEN_11 = taskWriteStateReg == 4'hc;
	wire io_connStealNtw_ctrl_serveStealReq_valid_0 = |tasksGivenAwayCount & (taskWriteStateReg != 4'hc);
	always @(posedge clock)
		if (reset) begin
			counterStateReg <= 4'h1;
			counterReg <= 64'h0000000000000000;
			currReadAddr <= 64'h0000000000000000;
			counterAddr <= 64'h0000000000000000;
			addrMask <= 64'h0000000000000000;
			helpGarbageCollector <= 1'h0;
			taskReadAddressStateReg <= 4'h6;
			taskAddr <= 64'h0000000000000000;
			taskReadStateReg <= 4'h9;
			taskReadCount <= 2'h3;
			taskRegisters_0 <= 32'h00000000;
			taskRegisters_1 <= 32'h00000000;
			taskRegisters_2 <= 32'h00000000;
			taskRegisters_3 <= 32'h00000000;
			tasksGivenAwayCount <= 32'h00000000;
			taskReg <= 128'h00000000000000000000000000000000;
			taskWriteStateReg <= 4'hb;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_12;
			reg _GEN_13;
			reg [1:0] _taskReadCount_T;
			reg _GEN_14;
			_GEN_12 = io_read_data_valid & (io_read_data_bits == 32'h00000001);
			_GEN_13 = _GEN_5 & _addressesOfReadyTasks_io_enq_ready;
			_taskReadCount_T = taskReadCount - 2'h1;
			_GEN_14 = _GEN_11 & io_connStealNtw_data_qOutTask_ready;
			if (_GEN) begin
				if (_addrNtwInQueue_io_deq_valid)
					counterStateReg <= 4'h2;
			end
			else if (_GEN_0) begin
				if (io_read_address_ready)
					counterStateReg <= 4'h3;
			end
			else if (_GEN_1) begin
				if (_GEN_12)
					counterStateReg <= 4'h7;
				else if (io_read_data_valid)
					counterStateReg <= 4'h4;
			end
			else if (_GEN_3) begin
				if (io_write_address_ready)
					counterStateReg <= 4'h5;
			end
			else if (_GEN_4) begin
				if (io_write_data_ready)
					counterStateReg <= 4'h1;
			end
			else if (_GEN_13)
				counterStateReg <= 4'h4;
			if (((_GEN_2 | ~_GEN_1) | _GEN_12) | ~io_read_data_valid)
				;
			else
				counterReg <= {32'h00000000, io_read_data_bits - 32'h00000001};
			if (_GEN_2 | ~(_GEN_1 & _GEN_12))
				;
			else
				currReadAddr <= counterAddr + 64'h0000000000000004;
			if (_GEN & _addrNtwInQueue_io_deq_valid)
				counterAddr <= _addrNtwInQueue_io_deq_bits & addrMask;
			addrMask <= 64'hfffffffffffffff0;
			if (~_GEN_6) begin
				if (_GEN_4)
					helpGarbageCollector <= ~io_write_data_ready & helpGarbageCollector;
				else
					helpGarbageCollector <= _GEN_13 | helpGarbageCollector;
			end
			if (_GEN_7) begin
				if (_addressesOfReadyTasks_io_deq_valid)
					taskReadAddressStateReg <= 4'h8;
			end
			else if (_GEN_8 & io_read_address_task_ready)
				taskReadAddressStateReg <= 4'h6;
			if (_GEN_7 & _addressesOfReadyTasks_io_deq_valid)
				taskAddr <= _addressesOfReadyTasks_io_deq_bits;
			if (io_read_data_task_ready_0) begin
				if ((taskReadCount == 2'h1) & io_read_data_task_valid)
					taskReadStateReg <= 4'ha;
				if (io_read_data_task_valid)
					taskReadCount <= _taskReadCount_T;
			end
			else if (_GEN_9 & _readyTasksQueue_io_enq_ready) begin
				taskReadStateReg <= 4'h9;
				taskReadCount <= 2'h3;
			end
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 2'h0))
				taskRegisters_0 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 2'h1))
				taskRegisters_1 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (_taskReadCount_T == 2'h2))
				taskRegisters_2 <= io_read_data_task_bits;
			if ((io_read_data_task_ready_0 & io_read_data_task_valid) & (&_taskReadCount_T))
				taskRegisters_3 <= io_read_data_task_bits;
			if (io_connStealNtw_ctrl_serveStealReq_valid_0 & io_connStealNtw_ctrl_serveStealReq_ready)
				tasksGivenAwayCount <= tasksGivenAwayCount - 32'h00000001;
			else if (_GEN_10 | ~_GEN_14)
				;
			else
				tasksGivenAwayCount <= tasksGivenAwayCount + 32'h00000001;
			if (_GEN_10 & _readyTasksQueue_io_deq_valid)
				taskReg <= _readyTasksQueue_io_deq_bits;
			if (_GEN_10) begin
				if (_readyTasksQueue_io_deq_valid)
					taskWriteStateReg <= 4'hc;
			end
			else if (_GEN_14)
				taskWriteStateReg <= 4'hb;
		end
	Queue16_UInt addrNtwInQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(io_connNetwork_ready),
		.io_enq_valid(io_connNetwork_valid),
		.io_enq_bits(io_connNetwork_bits),
		.io_deq_ready(_GEN),
		.io_deq_valid(_addrNtwInQueue_io_deq_valid),
		.io_deq_bits(_addrNtwInQueue_io_deq_bits)
	);
	Queue16_UInt addressesOfReadyTasks(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_addressesOfReadyTasks_io_enq_ready),
		.io_enq_valid(~((((_GEN | _GEN_0) | _GEN_1) | _GEN_3) | _GEN_4) & _GEN_5),
		.io_enq_bits(currReadAddr),
		.io_deq_ready(_GEN_7),
		.io_deq_valid(_addressesOfReadyTasks_io_deq_valid),
		.io_deq_bits(_addressesOfReadyTasks_io_deq_bits)
	);
	Queue16_UInt_2 readyTasksQueue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_readyTasksQueue_io_enq_ready),
		.io_enq_valid(~io_read_data_task_ready_0 & _GEN_9),
		.io_enq_bits({taskRegisters_0, taskRegisters_1, taskRegisters_2, taskRegisters_3}),
		.io_deq_ready(_GEN_10),
		.io_deq_valid(_readyTasksQueue_io_deq_valid),
		.io_deq_bits(_readyTasksQueue_io_deq_bits)
	);
	assign io_connStealNtw_ctrl_serveStealReq_valid = io_connStealNtw_ctrl_serveStealReq_valid_0;
	assign io_connStealNtw_data_qOutTask_valid = ~_GEN_10 & _GEN_11;
	assign io_connStealNtw_data_qOutTask_bits = taskReg;
	assign io_read_address_valid = ~_GEN & _GEN_0;
	assign io_read_address_bits = counterAddr;
	assign io_read_data_ready = ~_GEN_2 & _GEN_1;
	assign io_write_address_valid = ~((_GEN | _GEN_0) | _GEN_1) & _GEN_3;
	assign io_write_address_bits = counterAddr;
	assign io_write_data_valid = ~_GEN_6 & _GEN_4;
	assign io_write_data_bits = (helpGarbageCollector ? 32'h01000000 : counterReg[31:0]);
	assign io_read_address_task_valid = ~_GEN_7 & _GEN_8;
	assign io_read_address_task_bits = (_GEN_7 | ~_GEN_8 ? 64'h0000000000000000 : taskAddr);
	assign io_read_data_task_ready = io_read_data_task_ready_0;
endmodule
module RVtoAXIBridge_6 (
	clock,
	reset,
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	io_write_address_ready,
	io_write_address_valid,
	io_write_address_bits,
	io_write_data_ready,
	io_write_data_valid,
	io_write_data_bits,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data,
	axi_aw_ready,
	axi_aw_valid,
	axi_aw_bits_addr,
	axi_w_ready,
	axi_w_valid,
	axi_w_bits_data,
	axi_b_valid
);
	input clock;
	input reset;
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [31:0] io_read_data_bits;
	output wire io_write_address_ready;
	input io_write_address_valid;
	input [63:0] io_write_address_bits;
	output wire io_write_data_ready;
	input io_write_data_valid;
	input [31:0] io_write_data_bits;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire axi_r_ready;
	input axi_r_valid;
	input [31:0] axi_r_bits_data;
	input axi_aw_ready;
	output wire axi_aw_valid;
	output wire [63:0] axi_aw_bits_addr;
	input axi_w_ready;
	output wire axi_w_valid;
	output wire [31:0] axi_w_bits_data;
	input axi_b_valid;
	reg [1:0] writeDataDone;
	reg writeHandshakeDetector;
	wire axi_w_valid_0 = (io_write_data_valid & axi_w_ready) & ~writeHandshakeDetector;
	always @(posedge clock)
		if (reset) begin
			writeDataDone <= 2'h0;
			writeHandshakeDetector <= 1'h0;
		end
		else begin
			if ((writeDataDone == 2'h0) & axi_w_ready)
				writeDataDone <= 2'h1;
			else if ((writeDataDone == 2'h1) & axi_b_valid)
				writeDataDone <= 2'h0;
			writeHandshakeDetector <= axi_w_valid_0 | (~axi_b_valid & writeHandshakeDetector);
		end
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign io_write_address_ready = axi_aw_ready;
	assign io_write_data_ready = (writeDataDone == 2'h1) & axi_b_valid;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_r_ready = io_read_data_ready;
	assign axi_aw_valid = io_write_address_valid;
	assign axi_aw_bits_addr = io_write_address_bits;
	assign axi_w_valid = axi_w_valid_0;
	assign axi_w_bits_data = io_write_data_bits;
endmodule
module RVtoAXIBridge_22 (
	io_read_address_ready,
	io_read_address_valid,
	io_read_address_bits,
	io_read_data_ready,
	io_read_data_valid,
	io_read_data_bits,
	axi_ar_ready,
	axi_ar_valid,
	axi_ar_bits_addr,
	axi_r_ready,
	axi_r_valid,
	axi_r_bits_data
);
	output wire io_read_address_ready;
	input io_read_address_valid;
	input [63:0] io_read_address_bits;
	input io_read_data_ready;
	output wire io_read_data_valid;
	output wire [31:0] io_read_data_bits;
	input axi_ar_ready;
	output wire axi_ar_valid;
	output wire [63:0] axi_ar_bits_addr;
	output wire axi_r_ready;
	input axi_r_valid;
	input [31:0] axi_r_bits_data;
	assign io_read_address_ready = axi_ar_ready;
	assign io_read_data_valid = axi_r_valid;
	assign io_read_data_bits = axi_r_bits_data;
	assign axi_ar_valid = io_read_address_valid;
	assign axi_ar_bits_addr = io_read_address_bits;
	assign axi_r_ready = io_read_data_ready;
endmodule
module AxisUpscaler_64 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [31:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [63:0] io_dataOut_TDATA;
	reg [63:0] buffer;
	reg readCounter;
	reg stateReg;
	always @(posedge clock)
		if (reset) begin
			buffer <= 64'h0000000000000000;
			readCounter <= 1'h0;
			stateReg <= 1'h0;
		end
		else if (stateReg) begin : sv2v_autoblock_1
			reg _GEN;
			_GEN = stateReg & io_dataOut_TREADY;
			readCounter <= ~_GEN & readCounter;
			stateReg <= ~_GEN & stateReg;
		end
		else begin : sv2v_autoblock_2
			reg _GEN_0;
			reg [158:0] _GEN_1;
			reg [158:0] _GEN_2;
			reg _GEN_3;
			_GEN_0 = io_dataIn_TVALID & ~readCounter;
			_GEN_1 = {127'h00000000000000000000000000000000, io_dataIn_TDATA};
			_GEN_2 = {153'h000000000000000000000000000000000000000, readCounter, 5'h00};
			_GEN_3 = io_dataIn_TVALID & readCounter;
			if (_GEN_0) begin : sv2v_autoblock_3
				reg [158:0] _buffer_T_1;
				_buffer_T_1 = _GEN_1 << _GEN_2;
				buffer <= buffer | _buffer_T_1[63:0];
				readCounter <= readCounter - 1'h1;
			end
			else begin : sv2v_autoblock_4
				reg [158:0] _buffer_T_4;
				_buffer_T_4 = _GEN_1 << _GEN_2;
				buffer <= ({64 {_GEN_3}} & _buffer_T_4[63:0]) | buffer;
			end
			stateReg <= (~_GEN_0 & _GEN_3) | stateReg;
		end
	assign io_dataIn_TREADY = ~stateReg;
	assign io_dataOut_TVALID = stateReg;
	assign io_dataOut_TDATA = buffer;
endmodule
module AxisDataWidthConverter_208 (
	clock,
	reset,
	io_dataIn_TREADY,
	io_dataIn_TVALID,
	io_dataIn_TDATA,
	io_dataOut_TREADY,
	io_dataOut_TVALID,
	io_dataOut_TDATA
);
	input clock;
	input reset;
	output wire io_dataIn_TREADY;
	input io_dataIn_TVALID;
	input [31:0] io_dataIn_TDATA;
	input io_dataOut_TREADY;
	output wire io_dataOut_TVALID;
	output wire [63:0] io_dataOut_TDATA;
	AxisUpscaler_64 upScaler(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(io_dataIn_TREADY),
		.io_dataIn_TVALID(io_dataIn_TVALID),
		.io_dataIn_TDATA(io_dataIn_TDATA),
		.io_dataOut_TREADY(io_dataOut_TREADY),
		.io_dataOut_TVALID(io_dataOut_TVALID),
		.io_dataOut_TDATA(io_dataOut_TDATA)
	);
endmodule
module Counter64 (
	clock,
	reset,
	io_signals_0,
	io_signals_1,
	io_signals_2,
	io_signals_3,
	io_signals_4,
	io_signals_5,
	io_signals_6,
	io_signals_7,
	io_signals_8,
	io_signals_9,
	io_signals_10,
	io_signals_11,
	io_signals_12,
	io_signals_13,
	io_signals_14,
	io_signals_15,
	io_signals_16,
	io_signals_17,
	io_signals_18,
	io_signals_19,
	io_signals_20,
	io_signals_21,
	io_signals_22,
	io_signals_23,
	io_signals_24,
	io_signals_25,
	io_signals_26,
	io_signals_27,
	io_signals_28,
	io_signals_29,
	io_signals_30,
	io_signals_31,
	io_signals_32,
	io_signals_33,
	io_signals_34,
	io_signals_35,
	io_signals_36,
	io_signals_37,
	io_signals_38,
	io_signals_39,
	io_signals_40,
	io_signals_41,
	io_signals_42,
	io_signals_43,
	io_signals_44,
	io_signals_45,
	io_signals_46,
	io_signals_47,
	io_signals_48,
	io_signals_49,
	io_signals_50,
	io_signals_51,
	io_signals_52,
	io_signals_53,
	io_signals_54,
	io_signals_55,
	io_signals_56,
	io_signals_57,
	io_signals_58,
	io_signals_59,
	io_signals_60,
	io_signals_61,
	io_signals_62,
	io_signals_63,
	io_signals_64,
	io_signals_65,
	io_signals_66,
	io_signals_67,
	io_signals_68,
	io_signals_69,
	io_signals_70,
	io_signals_71,
	io_signals_72,
	io_signals_73,
	io_signals_74,
	io_signals_75,
	io_signals_76,
	io_signals_77,
	io_signals_78,
	io_signals_79,
	io_counter
);
	input clock;
	input reset;
	input io_signals_0;
	input io_signals_1;
	input io_signals_2;
	input io_signals_3;
	input io_signals_4;
	input io_signals_5;
	input io_signals_6;
	input io_signals_7;
	input io_signals_8;
	input io_signals_9;
	input io_signals_10;
	input io_signals_11;
	input io_signals_12;
	input io_signals_13;
	input io_signals_14;
	input io_signals_15;
	input io_signals_16;
	input io_signals_17;
	input io_signals_18;
	input io_signals_19;
	input io_signals_20;
	input io_signals_21;
	input io_signals_22;
	input io_signals_23;
	input io_signals_24;
	input io_signals_25;
	input io_signals_26;
	input io_signals_27;
	input io_signals_28;
	input io_signals_29;
	input io_signals_30;
	input io_signals_31;
	input io_signals_32;
	input io_signals_33;
	input io_signals_34;
	input io_signals_35;
	input io_signals_36;
	input io_signals_37;
	input io_signals_38;
	input io_signals_39;
	input io_signals_40;
	input io_signals_41;
	input io_signals_42;
	input io_signals_43;
	input io_signals_44;
	input io_signals_45;
	input io_signals_46;
	input io_signals_47;
	input io_signals_48;
	input io_signals_49;
	input io_signals_50;
	input io_signals_51;
	input io_signals_52;
	input io_signals_53;
	input io_signals_54;
	input io_signals_55;
	input io_signals_56;
	input io_signals_57;
	input io_signals_58;
	input io_signals_59;
	input io_signals_60;
	input io_signals_61;
	input io_signals_62;
	input io_signals_63;
	input io_signals_64;
	input io_signals_65;
	input io_signals_66;
	input io_signals_67;
	input io_signals_68;
	input io_signals_69;
	input io_signals_70;
	input io_signals_71;
	input io_signals_72;
	input io_signals_73;
	input io_signals_74;
	input io_signals_75;
	input io_signals_76;
	input io_signals_77;
	input io_signals_78;
	input io_signals_79;
	output wire [63:0] io_counter;
	reg [63:0] counter;
	always @(posedge clock)
		if (reset)
			counter <= 64'h0000000000000000;
		else
			counter <= counter + {57'h000000000000000, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_0} + {1'h0, io_signals_1}} + {1'h0, ({1'h0, io_signals_2} + {1'h0, io_signals_3}) + {1'h0, io_signals_4}}} + {1'h0, {1'h0, {1'h0, io_signals_5} + {1'h0, io_signals_6}} + {1'h0, ({1'h0, io_signals_7} + {1'h0, io_signals_8}) + {1'h0, io_signals_9}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_10} + {1'h0, io_signals_11}} + {1'h0, ({1'h0, io_signals_12} + {1'h0, io_signals_13}) + {1'h0, io_signals_14}}} + {1'h0, {1'h0, {1'h0, io_signals_15} + {1'h0, io_signals_16}} + {1'h0, ({1'h0, io_signals_17} + {1'h0, io_signals_18}) + {1'h0, io_signals_19}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_20} + {1'h0, io_signals_21}} + {1'h0, ({1'h0, io_signals_22} + {1'h0, io_signals_23}) + {1'h0, io_signals_24}}} + {1'h0, {1'h0, {1'h0, io_signals_25} + {1'h0, io_signals_26}} + {1'h0, ({1'h0, io_signals_27} + {1'h0, io_signals_28}) + {1'h0, io_signals_29}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_30} + {1'h0, io_signals_31}} + {1'h0, ({1'h0, io_signals_32} + {1'h0, io_signals_33}) + {1'h0, io_signals_34}}} + {1'h0, {1'h0, {1'h0, io_signals_35} + {1'h0, io_signals_36}} + {1'h0, ({1'h0, io_signals_37} + {1'h0, io_signals_38}) + {1'h0, io_signals_39}}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_40} + {1'h0, io_signals_41}} + {1'h0, ({1'h0, io_signals_42} + {1'h0, io_signals_43}) + {1'h0, io_signals_44}}} + {1'h0, {1'h0, {1'h0, io_signals_45} + {1'h0, io_signals_46}} + {1'h0, ({1'h0, io_signals_47} + {1'h0, io_signals_48}) + {1'h0, io_signals_49}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_50} + {1'h0, io_signals_51}} + {1'h0, ({1'h0, io_signals_52} + {1'h0, io_signals_53}) + {1'h0, io_signals_54}}} + {1'h0, {1'h0, {1'h0, io_signals_55} + {1'h0, io_signals_56}} + {1'h0, ({1'h0, io_signals_57} + {1'h0, io_signals_58}) + {1'h0, io_signals_59}}}}} + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, io_signals_60} + {1'h0, io_signals_61}} + {1'h0, ({1'h0, io_signals_62} + {1'h0, io_signals_63}) + {1'h0, io_signals_64}}} + {1'h0, {1'h0, {1'h0, io_signals_65} + {1'h0, io_signals_66}} + {1'h0, ({1'h0, io_signals_67} + {1'h0, io_signals_68}) + {1'h0, io_signals_69}}}} + {1'h0, {1'h0, {1'h0, {1'h0, io_signals_70} + {1'h0, io_signals_71}} + {1'h0, ({1'h0, io_signals_72} + {1'h0, io_signals_73}) + {1'h0, io_signals_74}}} + {1'h0, {1'h0, {1'h0, io_signals_75} + {1'h0, io_signals_76}} + {1'h0, ({1'h0, io_signals_77} + {1'h0, io_signals_78}) + {1'h0, io_signals_79}}}}}}};
	assign io_counter = counter;
endmodule
module ArgumentNotifier (
	clock,
	reset,
	io_export_argIn_0_TREADY,
	io_export_argIn_0_TVALID,
	io_export_argIn_0_TDATA,
	io_export_argIn_1_TREADY,
	io_export_argIn_1_TVALID,
	io_export_argIn_1_TDATA,
	io_export_argIn_2_TREADY,
	io_export_argIn_2_TVALID,
	io_export_argIn_2_TDATA,
	io_export_argIn_3_TREADY,
	io_export_argIn_3_TVALID,
	io_export_argIn_3_TDATA,
	io_export_argIn_4_TREADY,
	io_export_argIn_4_TVALID,
	io_export_argIn_4_TDATA,
	io_export_argIn_5_TREADY,
	io_export_argIn_5_TVALID,
	io_export_argIn_5_TDATA,
	io_export_argIn_6_TREADY,
	io_export_argIn_6_TVALID,
	io_export_argIn_6_TDATA,
	io_export_argIn_7_TREADY,
	io_export_argIn_7_TVALID,
	io_export_argIn_7_TDATA,
	io_export_argIn_8_TREADY,
	io_export_argIn_8_TVALID,
	io_export_argIn_8_TDATA,
	io_export_argIn_9_TREADY,
	io_export_argIn_9_TVALID,
	io_export_argIn_9_TDATA,
	io_export_argIn_10_TREADY,
	io_export_argIn_10_TVALID,
	io_export_argIn_10_TDATA,
	io_export_argIn_11_TREADY,
	io_export_argIn_11_TVALID,
	io_export_argIn_11_TDATA,
	io_export_argIn_12_TREADY,
	io_export_argIn_12_TVALID,
	io_export_argIn_12_TDATA,
	io_export_argIn_13_TREADY,
	io_export_argIn_13_TVALID,
	io_export_argIn_13_TDATA,
	io_export_argIn_14_TREADY,
	io_export_argIn_14_TVALID,
	io_export_argIn_14_TDATA,
	io_export_argIn_15_TREADY,
	io_export_argIn_15_TVALID,
	io_export_argIn_15_TDATA,
	io_export_argIn_16_TREADY,
	io_export_argIn_16_TVALID,
	io_export_argIn_16_TDATA,
	io_export_argIn_17_TREADY,
	io_export_argIn_17_TVALID,
	io_export_argIn_17_TDATA,
	io_export_argIn_18_TREADY,
	io_export_argIn_18_TVALID,
	io_export_argIn_18_TDATA,
	io_export_argIn_19_TREADY,
	io_export_argIn_19_TVALID,
	io_export_argIn_19_TDATA,
	io_export_argIn_20_TREADY,
	io_export_argIn_20_TVALID,
	io_export_argIn_20_TDATA,
	io_export_argIn_21_TREADY,
	io_export_argIn_21_TVALID,
	io_export_argIn_21_TDATA,
	io_export_argIn_22_TREADY,
	io_export_argIn_22_TVALID,
	io_export_argIn_22_TDATA,
	io_export_argIn_23_TREADY,
	io_export_argIn_23_TVALID,
	io_export_argIn_23_TDATA,
	io_export_argIn_24_TREADY,
	io_export_argIn_24_TVALID,
	io_export_argIn_24_TDATA,
	io_export_argIn_25_TREADY,
	io_export_argIn_25_TVALID,
	io_export_argIn_25_TDATA,
	io_export_argIn_26_TREADY,
	io_export_argIn_26_TVALID,
	io_export_argIn_26_TDATA,
	io_export_argIn_27_TREADY,
	io_export_argIn_27_TVALID,
	io_export_argIn_27_TDATA,
	io_export_argIn_28_TREADY,
	io_export_argIn_28_TVALID,
	io_export_argIn_28_TDATA,
	io_export_argIn_29_TREADY,
	io_export_argIn_29_TVALID,
	io_export_argIn_29_TDATA,
	io_export_argIn_30_TREADY,
	io_export_argIn_30_TVALID,
	io_export_argIn_30_TDATA,
	io_export_argIn_31_TREADY,
	io_export_argIn_31_TVALID,
	io_export_argIn_31_TDATA,
	io_export_argIn_32_TREADY,
	io_export_argIn_32_TVALID,
	io_export_argIn_32_TDATA,
	io_export_argIn_33_TREADY,
	io_export_argIn_33_TVALID,
	io_export_argIn_33_TDATA,
	io_export_argIn_34_TREADY,
	io_export_argIn_34_TVALID,
	io_export_argIn_34_TDATA,
	io_export_argIn_35_TREADY,
	io_export_argIn_35_TVALID,
	io_export_argIn_35_TDATA,
	io_export_argIn_36_TREADY,
	io_export_argIn_36_TVALID,
	io_export_argIn_36_TDATA,
	io_export_argIn_37_TREADY,
	io_export_argIn_37_TVALID,
	io_export_argIn_37_TDATA,
	io_export_argIn_38_TREADY,
	io_export_argIn_38_TVALID,
	io_export_argIn_38_TDATA,
	io_export_argIn_39_TREADY,
	io_export_argIn_39_TVALID,
	io_export_argIn_39_TDATA,
	io_export_argIn_40_TREADY,
	io_export_argIn_40_TVALID,
	io_export_argIn_40_TDATA,
	io_export_argIn_41_TREADY,
	io_export_argIn_41_TVALID,
	io_export_argIn_41_TDATA,
	io_export_argIn_42_TREADY,
	io_export_argIn_42_TVALID,
	io_export_argIn_42_TDATA,
	io_export_argIn_43_TREADY,
	io_export_argIn_43_TVALID,
	io_export_argIn_43_TDATA,
	io_export_argIn_44_TREADY,
	io_export_argIn_44_TVALID,
	io_export_argIn_44_TDATA,
	io_export_argIn_45_TREADY,
	io_export_argIn_45_TVALID,
	io_export_argIn_45_TDATA,
	io_export_argIn_46_TREADY,
	io_export_argIn_46_TVALID,
	io_export_argIn_46_TDATA,
	io_export_argIn_47_TREADY,
	io_export_argIn_47_TVALID,
	io_export_argIn_47_TDATA,
	io_export_argIn_48_TREADY,
	io_export_argIn_48_TVALID,
	io_export_argIn_48_TDATA,
	io_export_argIn_49_TREADY,
	io_export_argIn_49_TVALID,
	io_export_argIn_49_TDATA,
	io_export_argIn_50_TREADY,
	io_export_argIn_50_TVALID,
	io_export_argIn_50_TDATA,
	io_export_argIn_51_TREADY,
	io_export_argIn_51_TVALID,
	io_export_argIn_51_TDATA,
	io_export_argIn_52_TREADY,
	io_export_argIn_52_TVALID,
	io_export_argIn_52_TDATA,
	io_export_argIn_53_TREADY,
	io_export_argIn_53_TVALID,
	io_export_argIn_53_TDATA,
	io_export_argIn_54_TREADY,
	io_export_argIn_54_TVALID,
	io_export_argIn_54_TDATA,
	io_export_argIn_55_TREADY,
	io_export_argIn_55_TVALID,
	io_export_argIn_55_TDATA,
	io_export_argIn_56_TREADY,
	io_export_argIn_56_TVALID,
	io_export_argIn_56_TDATA,
	io_export_argIn_57_TREADY,
	io_export_argIn_57_TVALID,
	io_export_argIn_57_TDATA,
	io_export_argIn_58_TREADY,
	io_export_argIn_58_TVALID,
	io_export_argIn_58_TDATA,
	io_export_argIn_59_TREADY,
	io_export_argIn_59_TVALID,
	io_export_argIn_59_TDATA,
	io_export_argIn_60_TREADY,
	io_export_argIn_60_TVALID,
	io_export_argIn_60_TDATA,
	io_export_argIn_61_TREADY,
	io_export_argIn_61_TVALID,
	io_export_argIn_61_TDATA,
	io_export_argIn_62_TREADY,
	io_export_argIn_62_TVALID,
	io_export_argIn_62_TDATA,
	io_export_argIn_63_TREADY,
	io_export_argIn_63_TVALID,
	io_export_argIn_63_TDATA,
	io_export_argIn_64_TREADY,
	io_export_argIn_64_TVALID,
	io_export_argIn_64_TDATA,
	io_export_argIn_65_TREADY,
	io_export_argIn_65_TVALID,
	io_export_argIn_65_TDATA,
	io_export_argIn_66_TREADY,
	io_export_argIn_66_TVALID,
	io_export_argIn_66_TDATA,
	io_export_argIn_67_TREADY,
	io_export_argIn_67_TVALID,
	io_export_argIn_67_TDATA,
	io_export_argIn_68_TREADY,
	io_export_argIn_68_TVALID,
	io_export_argIn_68_TDATA,
	io_export_argIn_69_TREADY,
	io_export_argIn_69_TVALID,
	io_export_argIn_69_TDATA,
	io_export_argIn_70_TREADY,
	io_export_argIn_70_TVALID,
	io_export_argIn_70_TDATA,
	io_export_argIn_71_TREADY,
	io_export_argIn_71_TVALID,
	io_export_argIn_71_TDATA,
	io_export_argIn_72_TREADY,
	io_export_argIn_72_TVALID,
	io_export_argIn_72_TDATA,
	io_export_argIn_73_TREADY,
	io_export_argIn_73_TVALID,
	io_export_argIn_73_TDATA,
	io_export_argIn_74_TREADY,
	io_export_argIn_74_TVALID,
	io_export_argIn_74_TDATA,
	io_export_argIn_75_TREADY,
	io_export_argIn_75_TVALID,
	io_export_argIn_75_TDATA,
	io_export_argIn_76_TREADY,
	io_export_argIn_76_TVALID,
	io_export_argIn_76_TDATA,
	io_export_argIn_77_TREADY,
	io_export_argIn_77_TVALID,
	io_export_argIn_77_TDATA,
	io_export_argIn_78_TREADY,
	io_export_argIn_78_TVALID,
	io_export_argIn_78_TDATA,
	io_export_argIn_79_TREADY,
	io_export_argIn_79_TVALID,
	io_export_argIn_79_TDATA,
	connStealNtw_0_ctrl_serveStealReq_valid,
	connStealNtw_0_ctrl_serveStealReq_ready,
	connStealNtw_0_data_qOutTask_ready,
	connStealNtw_0_data_qOutTask_valid,
	connStealNtw_0_data_qOutTask_bits,
	connStealNtw_1_ctrl_serveStealReq_valid,
	connStealNtw_1_ctrl_serveStealReq_ready,
	connStealNtw_1_data_qOutTask_ready,
	connStealNtw_1_data_qOutTask_valid,
	connStealNtw_1_data_qOutTask_bits,
	connStealNtw_2_ctrl_serveStealReq_valid,
	connStealNtw_2_ctrl_serveStealReq_ready,
	connStealNtw_2_data_qOutTask_ready,
	connStealNtw_2_data_qOutTask_valid,
	connStealNtw_2_data_qOutTask_bits,
	connStealNtw_3_ctrl_serveStealReq_valid,
	connStealNtw_3_ctrl_serveStealReq_ready,
	connStealNtw_3_data_qOutTask_ready,
	connStealNtw_3_data_qOutTask_valid,
	connStealNtw_3_data_qOutTask_bits,
	connStealNtw_4_ctrl_serveStealReq_valid,
	connStealNtw_4_ctrl_serveStealReq_ready,
	connStealNtw_4_data_qOutTask_ready,
	connStealNtw_4_data_qOutTask_valid,
	connStealNtw_4_data_qOutTask_bits,
	connStealNtw_5_ctrl_serveStealReq_valid,
	connStealNtw_5_ctrl_serveStealReq_ready,
	connStealNtw_5_data_qOutTask_ready,
	connStealNtw_5_data_qOutTask_valid,
	connStealNtw_5_data_qOutTask_bits,
	connStealNtw_6_ctrl_serveStealReq_valid,
	connStealNtw_6_ctrl_serveStealReq_ready,
	connStealNtw_6_data_qOutTask_ready,
	connStealNtw_6_data_qOutTask_valid,
	connStealNtw_6_data_qOutTask_bits,
	connStealNtw_7_ctrl_serveStealReq_valid,
	connStealNtw_7_ctrl_serveStealReq_ready,
	connStealNtw_7_data_qOutTask_ready,
	connStealNtw_7_data_qOutTask_valid,
	connStealNtw_7_data_qOutTask_bits,
	connStealNtw_8_ctrl_serveStealReq_valid,
	connStealNtw_8_ctrl_serveStealReq_ready,
	connStealNtw_8_data_qOutTask_ready,
	connStealNtw_8_data_qOutTask_valid,
	connStealNtw_8_data_qOutTask_bits,
	connStealNtw_9_ctrl_serveStealReq_valid,
	connStealNtw_9_ctrl_serveStealReq_ready,
	connStealNtw_9_data_qOutTask_ready,
	connStealNtw_9_data_qOutTask_valid,
	connStealNtw_9_data_qOutTask_bits,
	connStealNtw_10_ctrl_serveStealReq_valid,
	connStealNtw_10_ctrl_serveStealReq_ready,
	connStealNtw_10_data_qOutTask_ready,
	connStealNtw_10_data_qOutTask_valid,
	connStealNtw_10_data_qOutTask_bits,
	connStealNtw_11_ctrl_serveStealReq_valid,
	connStealNtw_11_ctrl_serveStealReq_ready,
	connStealNtw_11_data_qOutTask_ready,
	connStealNtw_11_data_qOutTask_valid,
	connStealNtw_11_data_qOutTask_bits,
	connStealNtw_12_ctrl_serveStealReq_valid,
	connStealNtw_12_ctrl_serveStealReq_ready,
	connStealNtw_12_data_qOutTask_ready,
	connStealNtw_12_data_qOutTask_valid,
	connStealNtw_12_data_qOutTask_bits,
	connStealNtw_13_ctrl_serveStealReq_valid,
	connStealNtw_13_ctrl_serveStealReq_ready,
	connStealNtw_13_data_qOutTask_ready,
	connStealNtw_13_data_qOutTask_valid,
	connStealNtw_13_data_qOutTask_bits,
	connStealNtw_14_ctrl_serveStealReq_valid,
	connStealNtw_14_ctrl_serveStealReq_ready,
	connStealNtw_14_data_qOutTask_ready,
	connStealNtw_14_data_qOutTask_valid,
	connStealNtw_14_data_qOutTask_bits,
	connStealNtw_15_ctrl_serveStealReq_valid,
	connStealNtw_15_ctrl_serveStealReq_ready,
	connStealNtw_15_data_qOutTask_ready,
	connStealNtw_15_data_qOutTask_valid,
	connStealNtw_15_data_qOutTask_bits,
	axi_full_argRoute_0_ar_ready,
	axi_full_argRoute_0_ar_valid,
	axi_full_argRoute_0_ar_bits_addr,
	axi_full_argRoute_0_r_ready,
	axi_full_argRoute_0_r_valid,
	axi_full_argRoute_0_r_bits_data,
	axi_full_argRoute_0_aw_ready,
	axi_full_argRoute_0_aw_valid,
	axi_full_argRoute_0_aw_bits_addr,
	axi_full_argRoute_0_w_ready,
	axi_full_argRoute_0_w_valid,
	axi_full_argRoute_0_w_bits_data,
	axi_full_argRoute_0_b_valid,
	axi_full_argRoute_1_ar_ready,
	axi_full_argRoute_1_ar_valid,
	axi_full_argRoute_1_ar_bits_addr,
	axi_full_argRoute_1_r_ready,
	axi_full_argRoute_1_r_valid,
	axi_full_argRoute_1_r_bits_data,
	axi_full_argRoute_1_aw_ready,
	axi_full_argRoute_1_aw_valid,
	axi_full_argRoute_1_aw_bits_addr,
	axi_full_argRoute_1_w_ready,
	axi_full_argRoute_1_w_valid,
	axi_full_argRoute_1_w_bits_data,
	axi_full_argRoute_1_b_valid,
	axi_full_argRoute_2_ar_ready,
	axi_full_argRoute_2_ar_valid,
	axi_full_argRoute_2_ar_bits_addr,
	axi_full_argRoute_2_r_ready,
	axi_full_argRoute_2_r_valid,
	axi_full_argRoute_2_r_bits_data,
	axi_full_argRoute_2_aw_ready,
	axi_full_argRoute_2_aw_valid,
	axi_full_argRoute_2_aw_bits_addr,
	axi_full_argRoute_2_w_ready,
	axi_full_argRoute_2_w_valid,
	axi_full_argRoute_2_w_bits_data,
	axi_full_argRoute_2_b_valid,
	axi_full_argRoute_3_ar_ready,
	axi_full_argRoute_3_ar_valid,
	axi_full_argRoute_3_ar_bits_addr,
	axi_full_argRoute_3_r_ready,
	axi_full_argRoute_3_r_valid,
	axi_full_argRoute_3_r_bits_data,
	axi_full_argRoute_3_aw_ready,
	axi_full_argRoute_3_aw_valid,
	axi_full_argRoute_3_aw_bits_addr,
	axi_full_argRoute_3_w_ready,
	axi_full_argRoute_3_w_valid,
	axi_full_argRoute_3_w_bits_data,
	axi_full_argRoute_3_b_valid,
	axi_full_argRoute_4_ar_ready,
	axi_full_argRoute_4_ar_valid,
	axi_full_argRoute_4_ar_bits_addr,
	axi_full_argRoute_4_r_ready,
	axi_full_argRoute_4_r_valid,
	axi_full_argRoute_4_r_bits_data,
	axi_full_argRoute_4_aw_ready,
	axi_full_argRoute_4_aw_valid,
	axi_full_argRoute_4_aw_bits_addr,
	axi_full_argRoute_4_w_ready,
	axi_full_argRoute_4_w_valid,
	axi_full_argRoute_4_w_bits_data,
	axi_full_argRoute_4_b_valid,
	axi_full_argRoute_5_ar_ready,
	axi_full_argRoute_5_ar_valid,
	axi_full_argRoute_5_ar_bits_addr,
	axi_full_argRoute_5_r_ready,
	axi_full_argRoute_5_r_valid,
	axi_full_argRoute_5_r_bits_data,
	axi_full_argRoute_5_aw_ready,
	axi_full_argRoute_5_aw_valid,
	axi_full_argRoute_5_aw_bits_addr,
	axi_full_argRoute_5_w_ready,
	axi_full_argRoute_5_w_valid,
	axi_full_argRoute_5_w_bits_data,
	axi_full_argRoute_5_b_valid,
	axi_full_argRoute_6_ar_ready,
	axi_full_argRoute_6_ar_valid,
	axi_full_argRoute_6_ar_bits_addr,
	axi_full_argRoute_6_r_ready,
	axi_full_argRoute_6_r_valid,
	axi_full_argRoute_6_r_bits_data,
	axi_full_argRoute_6_aw_ready,
	axi_full_argRoute_6_aw_valid,
	axi_full_argRoute_6_aw_bits_addr,
	axi_full_argRoute_6_w_ready,
	axi_full_argRoute_6_w_valid,
	axi_full_argRoute_6_w_bits_data,
	axi_full_argRoute_6_b_valid,
	axi_full_argRoute_7_ar_ready,
	axi_full_argRoute_7_ar_valid,
	axi_full_argRoute_7_ar_bits_addr,
	axi_full_argRoute_7_r_ready,
	axi_full_argRoute_7_r_valid,
	axi_full_argRoute_7_r_bits_data,
	axi_full_argRoute_7_aw_ready,
	axi_full_argRoute_7_aw_valid,
	axi_full_argRoute_7_aw_bits_addr,
	axi_full_argRoute_7_w_ready,
	axi_full_argRoute_7_w_valid,
	axi_full_argRoute_7_w_bits_data,
	axi_full_argRoute_7_b_valid,
	axi_full_argRoute_8_ar_ready,
	axi_full_argRoute_8_ar_valid,
	axi_full_argRoute_8_ar_bits_addr,
	axi_full_argRoute_8_r_ready,
	axi_full_argRoute_8_r_valid,
	axi_full_argRoute_8_r_bits_data,
	axi_full_argRoute_8_aw_ready,
	axi_full_argRoute_8_aw_valid,
	axi_full_argRoute_8_aw_bits_addr,
	axi_full_argRoute_8_w_ready,
	axi_full_argRoute_8_w_valid,
	axi_full_argRoute_8_w_bits_data,
	axi_full_argRoute_8_b_valid,
	axi_full_argRoute_9_ar_ready,
	axi_full_argRoute_9_ar_valid,
	axi_full_argRoute_9_ar_bits_addr,
	axi_full_argRoute_9_r_ready,
	axi_full_argRoute_9_r_valid,
	axi_full_argRoute_9_r_bits_data,
	axi_full_argRoute_9_aw_ready,
	axi_full_argRoute_9_aw_valid,
	axi_full_argRoute_9_aw_bits_addr,
	axi_full_argRoute_9_w_ready,
	axi_full_argRoute_9_w_valid,
	axi_full_argRoute_9_w_bits_data,
	axi_full_argRoute_9_b_valid,
	axi_full_argRoute_10_ar_ready,
	axi_full_argRoute_10_ar_valid,
	axi_full_argRoute_10_ar_bits_addr,
	axi_full_argRoute_10_r_ready,
	axi_full_argRoute_10_r_valid,
	axi_full_argRoute_10_r_bits_data,
	axi_full_argRoute_10_aw_ready,
	axi_full_argRoute_10_aw_valid,
	axi_full_argRoute_10_aw_bits_addr,
	axi_full_argRoute_10_w_ready,
	axi_full_argRoute_10_w_valid,
	axi_full_argRoute_10_w_bits_data,
	axi_full_argRoute_10_b_valid,
	axi_full_argRoute_11_ar_ready,
	axi_full_argRoute_11_ar_valid,
	axi_full_argRoute_11_ar_bits_addr,
	axi_full_argRoute_11_r_ready,
	axi_full_argRoute_11_r_valid,
	axi_full_argRoute_11_r_bits_data,
	axi_full_argRoute_11_aw_ready,
	axi_full_argRoute_11_aw_valid,
	axi_full_argRoute_11_aw_bits_addr,
	axi_full_argRoute_11_w_ready,
	axi_full_argRoute_11_w_valid,
	axi_full_argRoute_11_w_bits_data,
	axi_full_argRoute_11_b_valid,
	axi_full_argRoute_12_ar_ready,
	axi_full_argRoute_12_ar_valid,
	axi_full_argRoute_12_ar_bits_addr,
	axi_full_argRoute_12_r_ready,
	axi_full_argRoute_12_r_valid,
	axi_full_argRoute_12_r_bits_data,
	axi_full_argRoute_12_aw_ready,
	axi_full_argRoute_12_aw_valid,
	axi_full_argRoute_12_aw_bits_addr,
	axi_full_argRoute_12_w_ready,
	axi_full_argRoute_12_w_valid,
	axi_full_argRoute_12_w_bits_data,
	axi_full_argRoute_12_b_valid,
	axi_full_argRoute_13_ar_ready,
	axi_full_argRoute_13_ar_valid,
	axi_full_argRoute_13_ar_bits_addr,
	axi_full_argRoute_13_r_ready,
	axi_full_argRoute_13_r_valid,
	axi_full_argRoute_13_r_bits_data,
	axi_full_argRoute_13_aw_ready,
	axi_full_argRoute_13_aw_valid,
	axi_full_argRoute_13_aw_bits_addr,
	axi_full_argRoute_13_w_ready,
	axi_full_argRoute_13_w_valid,
	axi_full_argRoute_13_w_bits_data,
	axi_full_argRoute_13_b_valid,
	axi_full_argRoute_14_ar_ready,
	axi_full_argRoute_14_ar_valid,
	axi_full_argRoute_14_ar_bits_addr,
	axi_full_argRoute_14_r_ready,
	axi_full_argRoute_14_r_valid,
	axi_full_argRoute_14_r_bits_data,
	axi_full_argRoute_14_aw_ready,
	axi_full_argRoute_14_aw_valid,
	axi_full_argRoute_14_aw_bits_addr,
	axi_full_argRoute_14_w_ready,
	axi_full_argRoute_14_w_valid,
	axi_full_argRoute_14_w_bits_data,
	axi_full_argRoute_14_b_valid,
	axi_full_argRoute_15_ar_ready,
	axi_full_argRoute_15_ar_valid,
	axi_full_argRoute_15_ar_bits_addr,
	axi_full_argRoute_15_r_ready,
	axi_full_argRoute_15_r_valid,
	axi_full_argRoute_15_r_bits_data,
	axi_full_argRoute_15_aw_ready,
	axi_full_argRoute_15_aw_valid,
	axi_full_argRoute_15_aw_bits_addr,
	axi_full_argRoute_15_w_ready,
	axi_full_argRoute_15_w_valid,
	axi_full_argRoute_15_w_bits_data,
	axi_full_argRoute_15_b_valid,
	axi_full_argRoute_16_ar_ready,
	axi_full_argRoute_16_ar_valid,
	axi_full_argRoute_16_ar_bits_addr,
	axi_full_argRoute_16_r_ready,
	axi_full_argRoute_16_r_valid,
	axi_full_argRoute_16_r_bits_data,
	axi_full_argRoute_17_ar_ready,
	axi_full_argRoute_17_ar_valid,
	axi_full_argRoute_17_ar_bits_addr,
	axi_full_argRoute_17_r_ready,
	axi_full_argRoute_17_r_valid,
	axi_full_argRoute_17_r_bits_data,
	axi_full_argRoute_18_ar_ready,
	axi_full_argRoute_18_ar_valid,
	axi_full_argRoute_18_ar_bits_addr,
	axi_full_argRoute_18_r_ready,
	axi_full_argRoute_18_r_valid,
	axi_full_argRoute_18_r_bits_data,
	axi_full_argRoute_19_ar_ready,
	axi_full_argRoute_19_ar_valid,
	axi_full_argRoute_19_ar_bits_addr,
	axi_full_argRoute_19_r_ready,
	axi_full_argRoute_19_r_valid,
	axi_full_argRoute_19_r_bits_data,
	axi_full_argRoute_20_ar_ready,
	axi_full_argRoute_20_ar_valid,
	axi_full_argRoute_20_ar_bits_addr,
	axi_full_argRoute_20_r_ready,
	axi_full_argRoute_20_r_valid,
	axi_full_argRoute_20_r_bits_data,
	axi_full_argRoute_21_ar_ready,
	axi_full_argRoute_21_ar_valid,
	axi_full_argRoute_21_ar_bits_addr,
	axi_full_argRoute_21_r_ready,
	axi_full_argRoute_21_r_valid,
	axi_full_argRoute_21_r_bits_data,
	axi_full_argRoute_22_ar_ready,
	axi_full_argRoute_22_ar_valid,
	axi_full_argRoute_22_ar_bits_addr,
	axi_full_argRoute_22_r_ready,
	axi_full_argRoute_22_r_valid,
	axi_full_argRoute_22_r_bits_data,
	axi_full_argRoute_23_ar_ready,
	axi_full_argRoute_23_ar_valid,
	axi_full_argRoute_23_ar_bits_addr,
	axi_full_argRoute_23_r_ready,
	axi_full_argRoute_23_r_valid,
	axi_full_argRoute_23_r_bits_data,
	axi_full_argRoute_24_ar_ready,
	axi_full_argRoute_24_ar_valid,
	axi_full_argRoute_24_ar_bits_addr,
	axi_full_argRoute_24_r_ready,
	axi_full_argRoute_24_r_valid,
	axi_full_argRoute_24_r_bits_data,
	axi_full_argRoute_25_ar_ready,
	axi_full_argRoute_25_ar_valid,
	axi_full_argRoute_25_ar_bits_addr,
	axi_full_argRoute_25_r_ready,
	axi_full_argRoute_25_r_valid,
	axi_full_argRoute_25_r_bits_data,
	axi_full_argRoute_26_ar_ready,
	axi_full_argRoute_26_ar_valid,
	axi_full_argRoute_26_ar_bits_addr,
	axi_full_argRoute_26_r_ready,
	axi_full_argRoute_26_r_valid,
	axi_full_argRoute_26_r_bits_data,
	axi_full_argRoute_27_ar_ready,
	axi_full_argRoute_27_ar_valid,
	axi_full_argRoute_27_ar_bits_addr,
	axi_full_argRoute_27_r_ready,
	axi_full_argRoute_27_r_valid,
	axi_full_argRoute_27_r_bits_data,
	axi_full_argRoute_28_ar_ready,
	axi_full_argRoute_28_ar_valid,
	axi_full_argRoute_28_ar_bits_addr,
	axi_full_argRoute_28_r_ready,
	axi_full_argRoute_28_r_valid,
	axi_full_argRoute_28_r_bits_data,
	axi_full_argRoute_29_ar_ready,
	axi_full_argRoute_29_ar_valid,
	axi_full_argRoute_29_ar_bits_addr,
	axi_full_argRoute_29_r_ready,
	axi_full_argRoute_29_r_valid,
	axi_full_argRoute_29_r_bits_data,
	axi_full_argRoute_30_ar_ready,
	axi_full_argRoute_30_ar_valid,
	axi_full_argRoute_30_ar_bits_addr,
	axi_full_argRoute_30_r_ready,
	axi_full_argRoute_30_r_valid,
	axi_full_argRoute_30_r_bits_data,
	axi_full_argRoute_31_ar_ready,
	axi_full_argRoute_31_ar_valid,
	axi_full_argRoute_31_ar_bits_addr,
	axi_full_argRoute_31_r_ready,
	axi_full_argRoute_31_r_valid,
	axi_full_argRoute_31_r_bits_data
);
	input clock;
	input reset;
	output wire io_export_argIn_0_TREADY;
	input io_export_argIn_0_TVALID;
	input [31:0] io_export_argIn_0_TDATA;
	output wire io_export_argIn_1_TREADY;
	input io_export_argIn_1_TVALID;
	input [31:0] io_export_argIn_1_TDATA;
	output wire io_export_argIn_2_TREADY;
	input io_export_argIn_2_TVALID;
	input [31:0] io_export_argIn_2_TDATA;
	output wire io_export_argIn_3_TREADY;
	input io_export_argIn_3_TVALID;
	input [31:0] io_export_argIn_3_TDATA;
	output wire io_export_argIn_4_TREADY;
	input io_export_argIn_4_TVALID;
	input [31:0] io_export_argIn_4_TDATA;
	output wire io_export_argIn_5_TREADY;
	input io_export_argIn_5_TVALID;
	input [31:0] io_export_argIn_5_TDATA;
	output wire io_export_argIn_6_TREADY;
	input io_export_argIn_6_TVALID;
	input [31:0] io_export_argIn_6_TDATA;
	output wire io_export_argIn_7_TREADY;
	input io_export_argIn_7_TVALID;
	input [31:0] io_export_argIn_7_TDATA;
	output wire io_export_argIn_8_TREADY;
	input io_export_argIn_8_TVALID;
	input [31:0] io_export_argIn_8_TDATA;
	output wire io_export_argIn_9_TREADY;
	input io_export_argIn_9_TVALID;
	input [31:0] io_export_argIn_9_TDATA;
	output wire io_export_argIn_10_TREADY;
	input io_export_argIn_10_TVALID;
	input [31:0] io_export_argIn_10_TDATA;
	output wire io_export_argIn_11_TREADY;
	input io_export_argIn_11_TVALID;
	input [31:0] io_export_argIn_11_TDATA;
	output wire io_export_argIn_12_TREADY;
	input io_export_argIn_12_TVALID;
	input [31:0] io_export_argIn_12_TDATA;
	output wire io_export_argIn_13_TREADY;
	input io_export_argIn_13_TVALID;
	input [31:0] io_export_argIn_13_TDATA;
	output wire io_export_argIn_14_TREADY;
	input io_export_argIn_14_TVALID;
	input [31:0] io_export_argIn_14_TDATA;
	output wire io_export_argIn_15_TREADY;
	input io_export_argIn_15_TVALID;
	input [31:0] io_export_argIn_15_TDATA;
	output wire io_export_argIn_16_TREADY;
	input io_export_argIn_16_TVALID;
	input [31:0] io_export_argIn_16_TDATA;
	output wire io_export_argIn_17_TREADY;
	input io_export_argIn_17_TVALID;
	input [31:0] io_export_argIn_17_TDATA;
	output wire io_export_argIn_18_TREADY;
	input io_export_argIn_18_TVALID;
	input [31:0] io_export_argIn_18_TDATA;
	output wire io_export_argIn_19_TREADY;
	input io_export_argIn_19_TVALID;
	input [31:0] io_export_argIn_19_TDATA;
	output wire io_export_argIn_20_TREADY;
	input io_export_argIn_20_TVALID;
	input [31:0] io_export_argIn_20_TDATA;
	output wire io_export_argIn_21_TREADY;
	input io_export_argIn_21_TVALID;
	input [31:0] io_export_argIn_21_TDATA;
	output wire io_export_argIn_22_TREADY;
	input io_export_argIn_22_TVALID;
	input [31:0] io_export_argIn_22_TDATA;
	output wire io_export_argIn_23_TREADY;
	input io_export_argIn_23_TVALID;
	input [31:0] io_export_argIn_23_TDATA;
	output wire io_export_argIn_24_TREADY;
	input io_export_argIn_24_TVALID;
	input [31:0] io_export_argIn_24_TDATA;
	output wire io_export_argIn_25_TREADY;
	input io_export_argIn_25_TVALID;
	input [31:0] io_export_argIn_25_TDATA;
	output wire io_export_argIn_26_TREADY;
	input io_export_argIn_26_TVALID;
	input [31:0] io_export_argIn_26_TDATA;
	output wire io_export_argIn_27_TREADY;
	input io_export_argIn_27_TVALID;
	input [31:0] io_export_argIn_27_TDATA;
	output wire io_export_argIn_28_TREADY;
	input io_export_argIn_28_TVALID;
	input [31:0] io_export_argIn_28_TDATA;
	output wire io_export_argIn_29_TREADY;
	input io_export_argIn_29_TVALID;
	input [31:0] io_export_argIn_29_TDATA;
	output wire io_export_argIn_30_TREADY;
	input io_export_argIn_30_TVALID;
	input [31:0] io_export_argIn_30_TDATA;
	output wire io_export_argIn_31_TREADY;
	input io_export_argIn_31_TVALID;
	input [31:0] io_export_argIn_31_TDATA;
	output wire io_export_argIn_32_TREADY;
	input io_export_argIn_32_TVALID;
	input [31:0] io_export_argIn_32_TDATA;
	output wire io_export_argIn_33_TREADY;
	input io_export_argIn_33_TVALID;
	input [31:0] io_export_argIn_33_TDATA;
	output wire io_export_argIn_34_TREADY;
	input io_export_argIn_34_TVALID;
	input [31:0] io_export_argIn_34_TDATA;
	output wire io_export_argIn_35_TREADY;
	input io_export_argIn_35_TVALID;
	input [31:0] io_export_argIn_35_TDATA;
	output wire io_export_argIn_36_TREADY;
	input io_export_argIn_36_TVALID;
	input [31:0] io_export_argIn_36_TDATA;
	output wire io_export_argIn_37_TREADY;
	input io_export_argIn_37_TVALID;
	input [31:0] io_export_argIn_37_TDATA;
	output wire io_export_argIn_38_TREADY;
	input io_export_argIn_38_TVALID;
	input [31:0] io_export_argIn_38_TDATA;
	output wire io_export_argIn_39_TREADY;
	input io_export_argIn_39_TVALID;
	input [31:0] io_export_argIn_39_TDATA;
	output wire io_export_argIn_40_TREADY;
	input io_export_argIn_40_TVALID;
	input [31:0] io_export_argIn_40_TDATA;
	output wire io_export_argIn_41_TREADY;
	input io_export_argIn_41_TVALID;
	input [31:0] io_export_argIn_41_TDATA;
	output wire io_export_argIn_42_TREADY;
	input io_export_argIn_42_TVALID;
	input [31:0] io_export_argIn_42_TDATA;
	output wire io_export_argIn_43_TREADY;
	input io_export_argIn_43_TVALID;
	input [31:0] io_export_argIn_43_TDATA;
	output wire io_export_argIn_44_TREADY;
	input io_export_argIn_44_TVALID;
	input [31:0] io_export_argIn_44_TDATA;
	output wire io_export_argIn_45_TREADY;
	input io_export_argIn_45_TVALID;
	input [31:0] io_export_argIn_45_TDATA;
	output wire io_export_argIn_46_TREADY;
	input io_export_argIn_46_TVALID;
	input [31:0] io_export_argIn_46_TDATA;
	output wire io_export_argIn_47_TREADY;
	input io_export_argIn_47_TVALID;
	input [31:0] io_export_argIn_47_TDATA;
	output wire io_export_argIn_48_TREADY;
	input io_export_argIn_48_TVALID;
	input [31:0] io_export_argIn_48_TDATA;
	output wire io_export_argIn_49_TREADY;
	input io_export_argIn_49_TVALID;
	input [31:0] io_export_argIn_49_TDATA;
	output wire io_export_argIn_50_TREADY;
	input io_export_argIn_50_TVALID;
	input [31:0] io_export_argIn_50_TDATA;
	output wire io_export_argIn_51_TREADY;
	input io_export_argIn_51_TVALID;
	input [31:0] io_export_argIn_51_TDATA;
	output wire io_export_argIn_52_TREADY;
	input io_export_argIn_52_TVALID;
	input [31:0] io_export_argIn_52_TDATA;
	output wire io_export_argIn_53_TREADY;
	input io_export_argIn_53_TVALID;
	input [31:0] io_export_argIn_53_TDATA;
	output wire io_export_argIn_54_TREADY;
	input io_export_argIn_54_TVALID;
	input [31:0] io_export_argIn_54_TDATA;
	output wire io_export_argIn_55_TREADY;
	input io_export_argIn_55_TVALID;
	input [31:0] io_export_argIn_55_TDATA;
	output wire io_export_argIn_56_TREADY;
	input io_export_argIn_56_TVALID;
	input [31:0] io_export_argIn_56_TDATA;
	output wire io_export_argIn_57_TREADY;
	input io_export_argIn_57_TVALID;
	input [31:0] io_export_argIn_57_TDATA;
	output wire io_export_argIn_58_TREADY;
	input io_export_argIn_58_TVALID;
	input [31:0] io_export_argIn_58_TDATA;
	output wire io_export_argIn_59_TREADY;
	input io_export_argIn_59_TVALID;
	input [31:0] io_export_argIn_59_TDATA;
	output wire io_export_argIn_60_TREADY;
	input io_export_argIn_60_TVALID;
	input [31:0] io_export_argIn_60_TDATA;
	output wire io_export_argIn_61_TREADY;
	input io_export_argIn_61_TVALID;
	input [31:0] io_export_argIn_61_TDATA;
	output wire io_export_argIn_62_TREADY;
	input io_export_argIn_62_TVALID;
	input [31:0] io_export_argIn_62_TDATA;
	output wire io_export_argIn_63_TREADY;
	input io_export_argIn_63_TVALID;
	input [31:0] io_export_argIn_63_TDATA;
	output wire io_export_argIn_64_TREADY;
	input io_export_argIn_64_TVALID;
	input [31:0] io_export_argIn_64_TDATA;
	output wire io_export_argIn_65_TREADY;
	input io_export_argIn_65_TVALID;
	input [31:0] io_export_argIn_65_TDATA;
	output wire io_export_argIn_66_TREADY;
	input io_export_argIn_66_TVALID;
	input [31:0] io_export_argIn_66_TDATA;
	output wire io_export_argIn_67_TREADY;
	input io_export_argIn_67_TVALID;
	input [31:0] io_export_argIn_67_TDATA;
	output wire io_export_argIn_68_TREADY;
	input io_export_argIn_68_TVALID;
	input [31:0] io_export_argIn_68_TDATA;
	output wire io_export_argIn_69_TREADY;
	input io_export_argIn_69_TVALID;
	input [31:0] io_export_argIn_69_TDATA;
	output wire io_export_argIn_70_TREADY;
	input io_export_argIn_70_TVALID;
	input [31:0] io_export_argIn_70_TDATA;
	output wire io_export_argIn_71_TREADY;
	input io_export_argIn_71_TVALID;
	input [31:0] io_export_argIn_71_TDATA;
	output wire io_export_argIn_72_TREADY;
	input io_export_argIn_72_TVALID;
	input [31:0] io_export_argIn_72_TDATA;
	output wire io_export_argIn_73_TREADY;
	input io_export_argIn_73_TVALID;
	input [31:0] io_export_argIn_73_TDATA;
	output wire io_export_argIn_74_TREADY;
	input io_export_argIn_74_TVALID;
	input [31:0] io_export_argIn_74_TDATA;
	output wire io_export_argIn_75_TREADY;
	input io_export_argIn_75_TVALID;
	input [31:0] io_export_argIn_75_TDATA;
	output wire io_export_argIn_76_TREADY;
	input io_export_argIn_76_TVALID;
	input [31:0] io_export_argIn_76_TDATA;
	output wire io_export_argIn_77_TREADY;
	input io_export_argIn_77_TVALID;
	input [31:0] io_export_argIn_77_TDATA;
	output wire io_export_argIn_78_TREADY;
	input io_export_argIn_78_TVALID;
	input [31:0] io_export_argIn_78_TDATA;
	output wire io_export_argIn_79_TREADY;
	input io_export_argIn_79_TVALID;
	input [31:0] io_export_argIn_79_TDATA;
	output wire connStealNtw_0_ctrl_serveStealReq_valid;
	input connStealNtw_0_ctrl_serveStealReq_ready;
	input connStealNtw_0_data_qOutTask_ready;
	output wire connStealNtw_0_data_qOutTask_valid;
	output wire [127:0] connStealNtw_0_data_qOutTask_bits;
	output wire connStealNtw_1_ctrl_serveStealReq_valid;
	input connStealNtw_1_ctrl_serveStealReq_ready;
	input connStealNtw_1_data_qOutTask_ready;
	output wire connStealNtw_1_data_qOutTask_valid;
	output wire [127:0] connStealNtw_1_data_qOutTask_bits;
	output wire connStealNtw_2_ctrl_serveStealReq_valid;
	input connStealNtw_2_ctrl_serveStealReq_ready;
	input connStealNtw_2_data_qOutTask_ready;
	output wire connStealNtw_2_data_qOutTask_valid;
	output wire [127:0] connStealNtw_2_data_qOutTask_bits;
	output wire connStealNtw_3_ctrl_serveStealReq_valid;
	input connStealNtw_3_ctrl_serveStealReq_ready;
	input connStealNtw_3_data_qOutTask_ready;
	output wire connStealNtw_3_data_qOutTask_valid;
	output wire [127:0] connStealNtw_3_data_qOutTask_bits;
	output wire connStealNtw_4_ctrl_serveStealReq_valid;
	input connStealNtw_4_ctrl_serveStealReq_ready;
	input connStealNtw_4_data_qOutTask_ready;
	output wire connStealNtw_4_data_qOutTask_valid;
	output wire [127:0] connStealNtw_4_data_qOutTask_bits;
	output wire connStealNtw_5_ctrl_serveStealReq_valid;
	input connStealNtw_5_ctrl_serveStealReq_ready;
	input connStealNtw_5_data_qOutTask_ready;
	output wire connStealNtw_5_data_qOutTask_valid;
	output wire [127:0] connStealNtw_5_data_qOutTask_bits;
	output wire connStealNtw_6_ctrl_serveStealReq_valid;
	input connStealNtw_6_ctrl_serveStealReq_ready;
	input connStealNtw_6_data_qOutTask_ready;
	output wire connStealNtw_6_data_qOutTask_valid;
	output wire [127:0] connStealNtw_6_data_qOutTask_bits;
	output wire connStealNtw_7_ctrl_serveStealReq_valid;
	input connStealNtw_7_ctrl_serveStealReq_ready;
	input connStealNtw_7_data_qOutTask_ready;
	output wire connStealNtw_7_data_qOutTask_valid;
	output wire [127:0] connStealNtw_7_data_qOutTask_bits;
	output wire connStealNtw_8_ctrl_serveStealReq_valid;
	input connStealNtw_8_ctrl_serveStealReq_ready;
	input connStealNtw_8_data_qOutTask_ready;
	output wire connStealNtw_8_data_qOutTask_valid;
	output wire [127:0] connStealNtw_8_data_qOutTask_bits;
	output wire connStealNtw_9_ctrl_serveStealReq_valid;
	input connStealNtw_9_ctrl_serveStealReq_ready;
	input connStealNtw_9_data_qOutTask_ready;
	output wire connStealNtw_9_data_qOutTask_valid;
	output wire [127:0] connStealNtw_9_data_qOutTask_bits;
	output wire connStealNtw_10_ctrl_serveStealReq_valid;
	input connStealNtw_10_ctrl_serveStealReq_ready;
	input connStealNtw_10_data_qOutTask_ready;
	output wire connStealNtw_10_data_qOutTask_valid;
	output wire [127:0] connStealNtw_10_data_qOutTask_bits;
	output wire connStealNtw_11_ctrl_serveStealReq_valid;
	input connStealNtw_11_ctrl_serveStealReq_ready;
	input connStealNtw_11_data_qOutTask_ready;
	output wire connStealNtw_11_data_qOutTask_valid;
	output wire [127:0] connStealNtw_11_data_qOutTask_bits;
	output wire connStealNtw_12_ctrl_serveStealReq_valid;
	input connStealNtw_12_ctrl_serveStealReq_ready;
	input connStealNtw_12_data_qOutTask_ready;
	output wire connStealNtw_12_data_qOutTask_valid;
	output wire [127:0] connStealNtw_12_data_qOutTask_bits;
	output wire connStealNtw_13_ctrl_serveStealReq_valid;
	input connStealNtw_13_ctrl_serveStealReq_ready;
	input connStealNtw_13_data_qOutTask_ready;
	output wire connStealNtw_13_data_qOutTask_valid;
	output wire [127:0] connStealNtw_13_data_qOutTask_bits;
	output wire connStealNtw_14_ctrl_serveStealReq_valid;
	input connStealNtw_14_ctrl_serveStealReq_ready;
	input connStealNtw_14_data_qOutTask_ready;
	output wire connStealNtw_14_data_qOutTask_valid;
	output wire [127:0] connStealNtw_14_data_qOutTask_bits;
	output wire connStealNtw_15_ctrl_serveStealReq_valid;
	input connStealNtw_15_ctrl_serveStealReq_ready;
	input connStealNtw_15_data_qOutTask_ready;
	output wire connStealNtw_15_data_qOutTask_valid;
	output wire [127:0] connStealNtw_15_data_qOutTask_bits;
	input axi_full_argRoute_0_ar_ready;
	output wire axi_full_argRoute_0_ar_valid;
	output wire [63:0] axi_full_argRoute_0_ar_bits_addr;
	output wire axi_full_argRoute_0_r_ready;
	input axi_full_argRoute_0_r_valid;
	input [31:0] axi_full_argRoute_0_r_bits_data;
	input axi_full_argRoute_0_aw_ready;
	output wire axi_full_argRoute_0_aw_valid;
	output wire [63:0] axi_full_argRoute_0_aw_bits_addr;
	input axi_full_argRoute_0_w_ready;
	output wire axi_full_argRoute_0_w_valid;
	output wire [31:0] axi_full_argRoute_0_w_bits_data;
	input axi_full_argRoute_0_b_valid;
	input axi_full_argRoute_1_ar_ready;
	output wire axi_full_argRoute_1_ar_valid;
	output wire [63:0] axi_full_argRoute_1_ar_bits_addr;
	output wire axi_full_argRoute_1_r_ready;
	input axi_full_argRoute_1_r_valid;
	input [31:0] axi_full_argRoute_1_r_bits_data;
	input axi_full_argRoute_1_aw_ready;
	output wire axi_full_argRoute_1_aw_valid;
	output wire [63:0] axi_full_argRoute_1_aw_bits_addr;
	input axi_full_argRoute_1_w_ready;
	output wire axi_full_argRoute_1_w_valid;
	output wire [31:0] axi_full_argRoute_1_w_bits_data;
	input axi_full_argRoute_1_b_valid;
	input axi_full_argRoute_2_ar_ready;
	output wire axi_full_argRoute_2_ar_valid;
	output wire [63:0] axi_full_argRoute_2_ar_bits_addr;
	output wire axi_full_argRoute_2_r_ready;
	input axi_full_argRoute_2_r_valid;
	input [31:0] axi_full_argRoute_2_r_bits_data;
	input axi_full_argRoute_2_aw_ready;
	output wire axi_full_argRoute_2_aw_valid;
	output wire [63:0] axi_full_argRoute_2_aw_bits_addr;
	input axi_full_argRoute_2_w_ready;
	output wire axi_full_argRoute_2_w_valid;
	output wire [31:0] axi_full_argRoute_2_w_bits_data;
	input axi_full_argRoute_2_b_valid;
	input axi_full_argRoute_3_ar_ready;
	output wire axi_full_argRoute_3_ar_valid;
	output wire [63:0] axi_full_argRoute_3_ar_bits_addr;
	output wire axi_full_argRoute_3_r_ready;
	input axi_full_argRoute_3_r_valid;
	input [31:0] axi_full_argRoute_3_r_bits_data;
	input axi_full_argRoute_3_aw_ready;
	output wire axi_full_argRoute_3_aw_valid;
	output wire [63:0] axi_full_argRoute_3_aw_bits_addr;
	input axi_full_argRoute_3_w_ready;
	output wire axi_full_argRoute_3_w_valid;
	output wire [31:0] axi_full_argRoute_3_w_bits_data;
	input axi_full_argRoute_3_b_valid;
	input axi_full_argRoute_4_ar_ready;
	output wire axi_full_argRoute_4_ar_valid;
	output wire [63:0] axi_full_argRoute_4_ar_bits_addr;
	output wire axi_full_argRoute_4_r_ready;
	input axi_full_argRoute_4_r_valid;
	input [31:0] axi_full_argRoute_4_r_bits_data;
	input axi_full_argRoute_4_aw_ready;
	output wire axi_full_argRoute_4_aw_valid;
	output wire [63:0] axi_full_argRoute_4_aw_bits_addr;
	input axi_full_argRoute_4_w_ready;
	output wire axi_full_argRoute_4_w_valid;
	output wire [31:0] axi_full_argRoute_4_w_bits_data;
	input axi_full_argRoute_4_b_valid;
	input axi_full_argRoute_5_ar_ready;
	output wire axi_full_argRoute_5_ar_valid;
	output wire [63:0] axi_full_argRoute_5_ar_bits_addr;
	output wire axi_full_argRoute_5_r_ready;
	input axi_full_argRoute_5_r_valid;
	input [31:0] axi_full_argRoute_5_r_bits_data;
	input axi_full_argRoute_5_aw_ready;
	output wire axi_full_argRoute_5_aw_valid;
	output wire [63:0] axi_full_argRoute_5_aw_bits_addr;
	input axi_full_argRoute_5_w_ready;
	output wire axi_full_argRoute_5_w_valid;
	output wire [31:0] axi_full_argRoute_5_w_bits_data;
	input axi_full_argRoute_5_b_valid;
	input axi_full_argRoute_6_ar_ready;
	output wire axi_full_argRoute_6_ar_valid;
	output wire [63:0] axi_full_argRoute_6_ar_bits_addr;
	output wire axi_full_argRoute_6_r_ready;
	input axi_full_argRoute_6_r_valid;
	input [31:0] axi_full_argRoute_6_r_bits_data;
	input axi_full_argRoute_6_aw_ready;
	output wire axi_full_argRoute_6_aw_valid;
	output wire [63:0] axi_full_argRoute_6_aw_bits_addr;
	input axi_full_argRoute_6_w_ready;
	output wire axi_full_argRoute_6_w_valid;
	output wire [31:0] axi_full_argRoute_6_w_bits_data;
	input axi_full_argRoute_6_b_valid;
	input axi_full_argRoute_7_ar_ready;
	output wire axi_full_argRoute_7_ar_valid;
	output wire [63:0] axi_full_argRoute_7_ar_bits_addr;
	output wire axi_full_argRoute_7_r_ready;
	input axi_full_argRoute_7_r_valid;
	input [31:0] axi_full_argRoute_7_r_bits_data;
	input axi_full_argRoute_7_aw_ready;
	output wire axi_full_argRoute_7_aw_valid;
	output wire [63:0] axi_full_argRoute_7_aw_bits_addr;
	input axi_full_argRoute_7_w_ready;
	output wire axi_full_argRoute_7_w_valid;
	output wire [31:0] axi_full_argRoute_7_w_bits_data;
	input axi_full_argRoute_7_b_valid;
	input axi_full_argRoute_8_ar_ready;
	output wire axi_full_argRoute_8_ar_valid;
	output wire [63:0] axi_full_argRoute_8_ar_bits_addr;
	output wire axi_full_argRoute_8_r_ready;
	input axi_full_argRoute_8_r_valid;
	input [31:0] axi_full_argRoute_8_r_bits_data;
	input axi_full_argRoute_8_aw_ready;
	output wire axi_full_argRoute_8_aw_valid;
	output wire [63:0] axi_full_argRoute_8_aw_bits_addr;
	input axi_full_argRoute_8_w_ready;
	output wire axi_full_argRoute_8_w_valid;
	output wire [31:0] axi_full_argRoute_8_w_bits_data;
	input axi_full_argRoute_8_b_valid;
	input axi_full_argRoute_9_ar_ready;
	output wire axi_full_argRoute_9_ar_valid;
	output wire [63:0] axi_full_argRoute_9_ar_bits_addr;
	output wire axi_full_argRoute_9_r_ready;
	input axi_full_argRoute_9_r_valid;
	input [31:0] axi_full_argRoute_9_r_bits_data;
	input axi_full_argRoute_9_aw_ready;
	output wire axi_full_argRoute_9_aw_valid;
	output wire [63:0] axi_full_argRoute_9_aw_bits_addr;
	input axi_full_argRoute_9_w_ready;
	output wire axi_full_argRoute_9_w_valid;
	output wire [31:0] axi_full_argRoute_9_w_bits_data;
	input axi_full_argRoute_9_b_valid;
	input axi_full_argRoute_10_ar_ready;
	output wire axi_full_argRoute_10_ar_valid;
	output wire [63:0] axi_full_argRoute_10_ar_bits_addr;
	output wire axi_full_argRoute_10_r_ready;
	input axi_full_argRoute_10_r_valid;
	input [31:0] axi_full_argRoute_10_r_bits_data;
	input axi_full_argRoute_10_aw_ready;
	output wire axi_full_argRoute_10_aw_valid;
	output wire [63:0] axi_full_argRoute_10_aw_bits_addr;
	input axi_full_argRoute_10_w_ready;
	output wire axi_full_argRoute_10_w_valid;
	output wire [31:0] axi_full_argRoute_10_w_bits_data;
	input axi_full_argRoute_10_b_valid;
	input axi_full_argRoute_11_ar_ready;
	output wire axi_full_argRoute_11_ar_valid;
	output wire [63:0] axi_full_argRoute_11_ar_bits_addr;
	output wire axi_full_argRoute_11_r_ready;
	input axi_full_argRoute_11_r_valid;
	input [31:0] axi_full_argRoute_11_r_bits_data;
	input axi_full_argRoute_11_aw_ready;
	output wire axi_full_argRoute_11_aw_valid;
	output wire [63:0] axi_full_argRoute_11_aw_bits_addr;
	input axi_full_argRoute_11_w_ready;
	output wire axi_full_argRoute_11_w_valid;
	output wire [31:0] axi_full_argRoute_11_w_bits_data;
	input axi_full_argRoute_11_b_valid;
	input axi_full_argRoute_12_ar_ready;
	output wire axi_full_argRoute_12_ar_valid;
	output wire [63:0] axi_full_argRoute_12_ar_bits_addr;
	output wire axi_full_argRoute_12_r_ready;
	input axi_full_argRoute_12_r_valid;
	input [31:0] axi_full_argRoute_12_r_bits_data;
	input axi_full_argRoute_12_aw_ready;
	output wire axi_full_argRoute_12_aw_valid;
	output wire [63:0] axi_full_argRoute_12_aw_bits_addr;
	input axi_full_argRoute_12_w_ready;
	output wire axi_full_argRoute_12_w_valid;
	output wire [31:0] axi_full_argRoute_12_w_bits_data;
	input axi_full_argRoute_12_b_valid;
	input axi_full_argRoute_13_ar_ready;
	output wire axi_full_argRoute_13_ar_valid;
	output wire [63:0] axi_full_argRoute_13_ar_bits_addr;
	output wire axi_full_argRoute_13_r_ready;
	input axi_full_argRoute_13_r_valid;
	input [31:0] axi_full_argRoute_13_r_bits_data;
	input axi_full_argRoute_13_aw_ready;
	output wire axi_full_argRoute_13_aw_valid;
	output wire [63:0] axi_full_argRoute_13_aw_bits_addr;
	input axi_full_argRoute_13_w_ready;
	output wire axi_full_argRoute_13_w_valid;
	output wire [31:0] axi_full_argRoute_13_w_bits_data;
	input axi_full_argRoute_13_b_valid;
	input axi_full_argRoute_14_ar_ready;
	output wire axi_full_argRoute_14_ar_valid;
	output wire [63:0] axi_full_argRoute_14_ar_bits_addr;
	output wire axi_full_argRoute_14_r_ready;
	input axi_full_argRoute_14_r_valid;
	input [31:0] axi_full_argRoute_14_r_bits_data;
	input axi_full_argRoute_14_aw_ready;
	output wire axi_full_argRoute_14_aw_valid;
	output wire [63:0] axi_full_argRoute_14_aw_bits_addr;
	input axi_full_argRoute_14_w_ready;
	output wire axi_full_argRoute_14_w_valid;
	output wire [31:0] axi_full_argRoute_14_w_bits_data;
	input axi_full_argRoute_14_b_valid;
	input axi_full_argRoute_15_ar_ready;
	output wire axi_full_argRoute_15_ar_valid;
	output wire [63:0] axi_full_argRoute_15_ar_bits_addr;
	output wire axi_full_argRoute_15_r_ready;
	input axi_full_argRoute_15_r_valid;
	input [31:0] axi_full_argRoute_15_r_bits_data;
	input axi_full_argRoute_15_aw_ready;
	output wire axi_full_argRoute_15_aw_valid;
	output wire [63:0] axi_full_argRoute_15_aw_bits_addr;
	input axi_full_argRoute_15_w_ready;
	output wire axi_full_argRoute_15_w_valid;
	output wire [31:0] axi_full_argRoute_15_w_bits_data;
	input axi_full_argRoute_15_b_valid;
	input axi_full_argRoute_16_ar_ready;
	output wire axi_full_argRoute_16_ar_valid;
	output wire [63:0] axi_full_argRoute_16_ar_bits_addr;
	output wire axi_full_argRoute_16_r_ready;
	input axi_full_argRoute_16_r_valid;
	input [31:0] axi_full_argRoute_16_r_bits_data;
	input axi_full_argRoute_17_ar_ready;
	output wire axi_full_argRoute_17_ar_valid;
	output wire [63:0] axi_full_argRoute_17_ar_bits_addr;
	output wire axi_full_argRoute_17_r_ready;
	input axi_full_argRoute_17_r_valid;
	input [31:0] axi_full_argRoute_17_r_bits_data;
	input axi_full_argRoute_18_ar_ready;
	output wire axi_full_argRoute_18_ar_valid;
	output wire [63:0] axi_full_argRoute_18_ar_bits_addr;
	output wire axi_full_argRoute_18_r_ready;
	input axi_full_argRoute_18_r_valid;
	input [31:0] axi_full_argRoute_18_r_bits_data;
	input axi_full_argRoute_19_ar_ready;
	output wire axi_full_argRoute_19_ar_valid;
	output wire [63:0] axi_full_argRoute_19_ar_bits_addr;
	output wire axi_full_argRoute_19_r_ready;
	input axi_full_argRoute_19_r_valid;
	input [31:0] axi_full_argRoute_19_r_bits_data;
	input axi_full_argRoute_20_ar_ready;
	output wire axi_full_argRoute_20_ar_valid;
	output wire [63:0] axi_full_argRoute_20_ar_bits_addr;
	output wire axi_full_argRoute_20_r_ready;
	input axi_full_argRoute_20_r_valid;
	input [31:0] axi_full_argRoute_20_r_bits_data;
	input axi_full_argRoute_21_ar_ready;
	output wire axi_full_argRoute_21_ar_valid;
	output wire [63:0] axi_full_argRoute_21_ar_bits_addr;
	output wire axi_full_argRoute_21_r_ready;
	input axi_full_argRoute_21_r_valid;
	input [31:0] axi_full_argRoute_21_r_bits_data;
	input axi_full_argRoute_22_ar_ready;
	output wire axi_full_argRoute_22_ar_valid;
	output wire [63:0] axi_full_argRoute_22_ar_bits_addr;
	output wire axi_full_argRoute_22_r_ready;
	input axi_full_argRoute_22_r_valid;
	input [31:0] axi_full_argRoute_22_r_bits_data;
	input axi_full_argRoute_23_ar_ready;
	output wire axi_full_argRoute_23_ar_valid;
	output wire [63:0] axi_full_argRoute_23_ar_bits_addr;
	output wire axi_full_argRoute_23_r_ready;
	input axi_full_argRoute_23_r_valid;
	input [31:0] axi_full_argRoute_23_r_bits_data;
	input axi_full_argRoute_24_ar_ready;
	output wire axi_full_argRoute_24_ar_valid;
	output wire [63:0] axi_full_argRoute_24_ar_bits_addr;
	output wire axi_full_argRoute_24_r_ready;
	input axi_full_argRoute_24_r_valid;
	input [31:0] axi_full_argRoute_24_r_bits_data;
	input axi_full_argRoute_25_ar_ready;
	output wire axi_full_argRoute_25_ar_valid;
	output wire [63:0] axi_full_argRoute_25_ar_bits_addr;
	output wire axi_full_argRoute_25_r_ready;
	input axi_full_argRoute_25_r_valid;
	input [31:0] axi_full_argRoute_25_r_bits_data;
	input axi_full_argRoute_26_ar_ready;
	output wire axi_full_argRoute_26_ar_valid;
	output wire [63:0] axi_full_argRoute_26_ar_bits_addr;
	output wire axi_full_argRoute_26_r_ready;
	input axi_full_argRoute_26_r_valid;
	input [31:0] axi_full_argRoute_26_r_bits_data;
	input axi_full_argRoute_27_ar_ready;
	output wire axi_full_argRoute_27_ar_valid;
	output wire [63:0] axi_full_argRoute_27_ar_bits_addr;
	output wire axi_full_argRoute_27_r_ready;
	input axi_full_argRoute_27_r_valid;
	input [31:0] axi_full_argRoute_27_r_bits_data;
	input axi_full_argRoute_28_ar_ready;
	output wire axi_full_argRoute_28_ar_valid;
	output wire [63:0] axi_full_argRoute_28_ar_bits_addr;
	output wire axi_full_argRoute_28_r_ready;
	input axi_full_argRoute_28_r_valid;
	input [31:0] axi_full_argRoute_28_r_bits_data;
	input axi_full_argRoute_29_ar_ready;
	output wire axi_full_argRoute_29_ar_valid;
	output wire [63:0] axi_full_argRoute_29_ar_bits_addr;
	output wire axi_full_argRoute_29_r_ready;
	input axi_full_argRoute_29_r_valid;
	input [31:0] axi_full_argRoute_29_r_bits_data;
	input axi_full_argRoute_30_ar_ready;
	output wire axi_full_argRoute_30_ar_valid;
	output wire [63:0] axi_full_argRoute_30_ar_bits_addr;
	output wire axi_full_argRoute_30_r_ready;
	input axi_full_argRoute_30_r_valid;
	input [31:0] axi_full_argRoute_30_r_bits_data;
	input axi_full_argRoute_31_ar_ready;
	output wire axi_full_argRoute_31_ar_valid;
	output wire [63:0] axi_full_argRoute_31_ar_bits_addr;
	output wire axi_full_argRoute_31_r_ready;
	input axi_full_argRoute_31_r_valid;
	input [31:0] axi_full_argRoute_31_r_bits_data;
	wire _axis_stream_converters_in_79_io_dataIn_TREADY;
	wire _axis_stream_converters_in_79_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_79_io_dataOut_TDATA;
	wire _axis_stream_converters_in_78_io_dataIn_TREADY;
	wire _axis_stream_converters_in_78_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_78_io_dataOut_TDATA;
	wire _axis_stream_converters_in_77_io_dataIn_TREADY;
	wire _axis_stream_converters_in_77_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_77_io_dataOut_TDATA;
	wire _axis_stream_converters_in_76_io_dataIn_TREADY;
	wire _axis_stream_converters_in_76_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_76_io_dataOut_TDATA;
	wire _axis_stream_converters_in_75_io_dataIn_TREADY;
	wire _axis_stream_converters_in_75_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_75_io_dataOut_TDATA;
	wire _axis_stream_converters_in_74_io_dataIn_TREADY;
	wire _axis_stream_converters_in_74_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_74_io_dataOut_TDATA;
	wire _axis_stream_converters_in_73_io_dataIn_TREADY;
	wire _axis_stream_converters_in_73_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_73_io_dataOut_TDATA;
	wire _axis_stream_converters_in_72_io_dataIn_TREADY;
	wire _axis_stream_converters_in_72_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_72_io_dataOut_TDATA;
	wire _axis_stream_converters_in_71_io_dataIn_TREADY;
	wire _axis_stream_converters_in_71_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_71_io_dataOut_TDATA;
	wire _axis_stream_converters_in_70_io_dataIn_TREADY;
	wire _axis_stream_converters_in_70_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_70_io_dataOut_TDATA;
	wire _axis_stream_converters_in_69_io_dataIn_TREADY;
	wire _axis_stream_converters_in_69_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_69_io_dataOut_TDATA;
	wire _axis_stream_converters_in_68_io_dataIn_TREADY;
	wire _axis_stream_converters_in_68_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_68_io_dataOut_TDATA;
	wire _axis_stream_converters_in_67_io_dataIn_TREADY;
	wire _axis_stream_converters_in_67_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_67_io_dataOut_TDATA;
	wire _axis_stream_converters_in_66_io_dataIn_TREADY;
	wire _axis_stream_converters_in_66_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_66_io_dataOut_TDATA;
	wire _axis_stream_converters_in_65_io_dataIn_TREADY;
	wire _axis_stream_converters_in_65_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_65_io_dataOut_TDATA;
	wire _axis_stream_converters_in_64_io_dataIn_TREADY;
	wire _axis_stream_converters_in_64_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_64_io_dataOut_TDATA;
	wire _axis_stream_converters_in_63_io_dataIn_TREADY;
	wire _axis_stream_converters_in_63_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_63_io_dataOut_TDATA;
	wire _axis_stream_converters_in_62_io_dataIn_TREADY;
	wire _axis_stream_converters_in_62_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_62_io_dataOut_TDATA;
	wire _axis_stream_converters_in_61_io_dataIn_TREADY;
	wire _axis_stream_converters_in_61_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_61_io_dataOut_TDATA;
	wire _axis_stream_converters_in_60_io_dataIn_TREADY;
	wire _axis_stream_converters_in_60_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_60_io_dataOut_TDATA;
	wire _axis_stream_converters_in_59_io_dataIn_TREADY;
	wire _axis_stream_converters_in_59_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_59_io_dataOut_TDATA;
	wire _axis_stream_converters_in_58_io_dataIn_TREADY;
	wire _axis_stream_converters_in_58_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_58_io_dataOut_TDATA;
	wire _axis_stream_converters_in_57_io_dataIn_TREADY;
	wire _axis_stream_converters_in_57_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_57_io_dataOut_TDATA;
	wire _axis_stream_converters_in_56_io_dataIn_TREADY;
	wire _axis_stream_converters_in_56_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_56_io_dataOut_TDATA;
	wire _axis_stream_converters_in_55_io_dataIn_TREADY;
	wire _axis_stream_converters_in_55_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_55_io_dataOut_TDATA;
	wire _axis_stream_converters_in_54_io_dataIn_TREADY;
	wire _axis_stream_converters_in_54_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_54_io_dataOut_TDATA;
	wire _axis_stream_converters_in_53_io_dataIn_TREADY;
	wire _axis_stream_converters_in_53_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_53_io_dataOut_TDATA;
	wire _axis_stream_converters_in_52_io_dataIn_TREADY;
	wire _axis_stream_converters_in_52_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_52_io_dataOut_TDATA;
	wire _axis_stream_converters_in_51_io_dataIn_TREADY;
	wire _axis_stream_converters_in_51_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_51_io_dataOut_TDATA;
	wire _axis_stream_converters_in_50_io_dataIn_TREADY;
	wire _axis_stream_converters_in_50_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_50_io_dataOut_TDATA;
	wire _axis_stream_converters_in_49_io_dataIn_TREADY;
	wire _axis_stream_converters_in_49_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_49_io_dataOut_TDATA;
	wire _axis_stream_converters_in_48_io_dataIn_TREADY;
	wire _axis_stream_converters_in_48_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_48_io_dataOut_TDATA;
	wire _axis_stream_converters_in_47_io_dataIn_TREADY;
	wire _axis_stream_converters_in_47_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_47_io_dataOut_TDATA;
	wire _axis_stream_converters_in_46_io_dataIn_TREADY;
	wire _axis_stream_converters_in_46_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_46_io_dataOut_TDATA;
	wire _axis_stream_converters_in_45_io_dataIn_TREADY;
	wire _axis_stream_converters_in_45_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_45_io_dataOut_TDATA;
	wire _axis_stream_converters_in_44_io_dataIn_TREADY;
	wire _axis_stream_converters_in_44_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_44_io_dataOut_TDATA;
	wire _axis_stream_converters_in_43_io_dataIn_TREADY;
	wire _axis_stream_converters_in_43_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_43_io_dataOut_TDATA;
	wire _axis_stream_converters_in_42_io_dataIn_TREADY;
	wire _axis_stream_converters_in_42_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_42_io_dataOut_TDATA;
	wire _axis_stream_converters_in_41_io_dataIn_TREADY;
	wire _axis_stream_converters_in_41_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_41_io_dataOut_TDATA;
	wire _axis_stream_converters_in_40_io_dataIn_TREADY;
	wire _axis_stream_converters_in_40_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_40_io_dataOut_TDATA;
	wire _axis_stream_converters_in_39_io_dataIn_TREADY;
	wire _axis_stream_converters_in_39_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_39_io_dataOut_TDATA;
	wire _axis_stream_converters_in_38_io_dataIn_TREADY;
	wire _axis_stream_converters_in_38_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_38_io_dataOut_TDATA;
	wire _axis_stream_converters_in_37_io_dataIn_TREADY;
	wire _axis_stream_converters_in_37_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_37_io_dataOut_TDATA;
	wire _axis_stream_converters_in_36_io_dataIn_TREADY;
	wire _axis_stream_converters_in_36_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_36_io_dataOut_TDATA;
	wire _axis_stream_converters_in_35_io_dataIn_TREADY;
	wire _axis_stream_converters_in_35_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_35_io_dataOut_TDATA;
	wire _axis_stream_converters_in_34_io_dataIn_TREADY;
	wire _axis_stream_converters_in_34_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_34_io_dataOut_TDATA;
	wire _axis_stream_converters_in_33_io_dataIn_TREADY;
	wire _axis_stream_converters_in_33_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_33_io_dataOut_TDATA;
	wire _axis_stream_converters_in_32_io_dataIn_TREADY;
	wire _axis_stream_converters_in_32_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_32_io_dataOut_TDATA;
	wire _axis_stream_converters_in_31_io_dataIn_TREADY;
	wire _axis_stream_converters_in_31_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_31_io_dataOut_TDATA;
	wire _axis_stream_converters_in_30_io_dataIn_TREADY;
	wire _axis_stream_converters_in_30_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_30_io_dataOut_TDATA;
	wire _axis_stream_converters_in_29_io_dataIn_TREADY;
	wire _axis_stream_converters_in_29_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_29_io_dataOut_TDATA;
	wire _axis_stream_converters_in_28_io_dataIn_TREADY;
	wire _axis_stream_converters_in_28_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_28_io_dataOut_TDATA;
	wire _axis_stream_converters_in_27_io_dataIn_TREADY;
	wire _axis_stream_converters_in_27_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_27_io_dataOut_TDATA;
	wire _axis_stream_converters_in_26_io_dataIn_TREADY;
	wire _axis_stream_converters_in_26_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_26_io_dataOut_TDATA;
	wire _axis_stream_converters_in_25_io_dataIn_TREADY;
	wire _axis_stream_converters_in_25_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_25_io_dataOut_TDATA;
	wire _axis_stream_converters_in_24_io_dataIn_TREADY;
	wire _axis_stream_converters_in_24_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_24_io_dataOut_TDATA;
	wire _axis_stream_converters_in_23_io_dataIn_TREADY;
	wire _axis_stream_converters_in_23_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_23_io_dataOut_TDATA;
	wire _axis_stream_converters_in_22_io_dataIn_TREADY;
	wire _axis_stream_converters_in_22_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_22_io_dataOut_TDATA;
	wire _axis_stream_converters_in_21_io_dataIn_TREADY;
	wire _axis_stream_converters_in_21_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_21_io_dataOut_TDATA;
	wire _axis_stream_converters_in_20_io_dataIn_TREADY;
	wire _axis_stream_converters_in_20_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_20_io_dataOut_TDATA;
	wire _axis_stream_converters_in_19_io_dataIn_TREADY;
	wire _axis_stream_converters_in_19_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_19_io_dataOut_TDATA;
	wire _axis_stream_converters_in_18_io_dataIn_TREADY;
	wire _axis_stream_converters_in_18_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_18_io_dataOut_TDATA;
	wire _axis_stream_converters_in_17_io_dataIn_TREADY;
	wire _axis_stream_converters_in_17_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_17_io_dataOut_TDATA;
	wire _axis_stream_converters_in_16_io_dataIn_TREADY;
	wire _axis_stream_converters_in_16_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_16_io_dataOut_TDATA;
	wire _axis_stream_converters_in_15_io_dataIn_TREADY;
	wire _axis_stream_converters_in_15_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_15_io_dataOut_TDATA;
	wire _axis_stream_converters_in_14_io_dataIn_TREADY;
	wire _axis_stream_converters_in_14_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_14_io_dataOut_TDATA;
	wire _axis_stream_converters_in_13_io_dataIn_TREADY;
	wire _axis_stream_converters_in_13_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_13_io_dataOut_TDATA;
	wire _axis_stream_converters_in_12_io_dataIn_TREADY;
	wire _axis_stream_converters_in_12_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_12_io_dataOut_TDATA;
	wire _axis_stream_converters_in_11_io_dataIn_TREADY;
	wire _axis_stream_converters_in_11_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_11_io_dataOut_TDATA;
	wire _axis_stream_converters_in_10_io_dataIn_TREADY;
	wire _axis_stream_converters_in_10_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_10_io_dataOut_TDATA;
	wire _axis_stream_converters_in_9_io_dataIn_TREADY;
	wire _axis_stream_converters_in_9_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_9_io_dataOut_TDATA;
	wire _axis_stream_converters_in_8_io_dataIn_TREADY;
	wire _axis_stream_converters_in_8_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_8_io_dataOut_TDATA;
	wire _axis_stream_converters_in_7_io_dataIn_TREADY;
	wire _axis_stream_converters_in_7_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_7_io_dataOut_TDATA;
	wire _axis_stream_converters_in_6_io_dataIn_TREADY;
	wire _axis_stream_converters_in_6_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_6_io_dataOut_TDATA;
	wire _axis_stream_converters_in_5_io_dataIn_TREADY;
	wire _axis_stream_converters_in_5_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_5_io_dataOut_TDATA;
	wire _axis_stream_converters_in_4_io_dataIn_TREADY;
	wire _axis_stream_converters_in_4_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_4_io_dataOut_TDATA;
	wire _axis_stream_converters_in_3_io_dataIn_TREADY;
	wire _axis_stream_converters_in_3_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_3_io_dataOut_TDATA;
	wire _axis_stream_converters_in_2_io_dataIn_TREADY;
	wire _axis_stream_converters_in_2_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_2_io_dataOut_TDATA;
	wire _axis_stream_converters_in_1_io_dataIn_TREADY;
	wire _axis_stream_converters_in_1_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_1_io_dataOut_TDATA;
	wire _axis_stream_converters_in_0_io_dataIn_TREADY;
	wire _axis_stream_converters_in_0_io_dataOut_TVALID;
	wire [63:0] _axis_stream_converters_in_0_io_dataOut_TDATA;
	wire _argRouteRvmReadOnly_15_io_read_address_ready;
	wire _argRouteRvmReadOnly_15_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_15_io_read_data_bits;
	wire _argRouteRvmReadOnly_14_io_read_address_ready;
	wire _argRouteRvmReadOnly_14_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_14_io_read_data_bits;
	wire _argRouteRvmReadOnly_13_io_read_address_ready;
	wire _argRouteRvmReadOnly_13_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_13_io_read_data_bits;
	wire _argRouteRvmReadOnly_12_io_read_address_ready;
	wire _argRouteRvmReadOnly_12_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_12_io_read_data_bits;
	wire _argRouteRvmReadOnly_11_io_read_address_ready;
	wire _argRouteRvmReadOnly_11_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_11_io_read_data_bits;
	wire _argRouteRvmReadOnly_10_io_read_address_ready;
	wire _argRouteRvmReadOnly_10_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_10_io_read_data_bits;
	wire _argRouteRvmReadOnly_9_io_read_address_ready;
	wire _argRouteRvmReadOnly_9_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_9_io_read_data_bits;
	wire _argRouteRvmReadOnly_8_io_read_address_ready;
	wire _argRouteRvmReadOnly_8_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_8_io_read_data_bits;
	wire _argRouteRvmReadOnly_7_io_read_address_ready;
	wire _argRouteRvmReadOnly_7_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_7_io_read_data_bits;
	wire _argRouteRvmReadOnly_6_io_read_address_ready;
	wire _argRouteRvmReadOnly_6_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_6_io_read_data_bits;
	wire _argRouteRvmReadOnly_5_io_read_address_ready;
	wire _argRouteRvmReadOnly_5_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_5_io_read_data_bits;
	wire _argRouteRvmReadOnly_4_io_read_address_ready;
	wire _argRouteRvmReadOnly_4_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_4_io_read_data_bits;
	wire _argRouteRvmReadOnly_3_io_read_address_ready;
	wire _argRouteRvmReadOnly_3_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_3_io_read_data_bits;
	wire _argRouteRvmReadOnly_2_io_read_address_ready;
	wire _argRouteRvmReadOnly_2_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_2_io_read_data_bits;
	wire _argRouteRvmReadOnly_1_io_read_address_ready;
	wire _argRouteRvmReadOnly_1_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_1_io_read_data_bits;
	wire _argRouteRvmReadOnly_0_io_read_address_ready;
	wire _argRouteRvmReadOnly_0_io_read_data_valid;
	wire [31:0] _argRouteRvmReadOnly_0_io_read_data_bits;
	wire _argRouteRvm_15_io_read_address_ready;
	wire _argRouteRvm_15_io_read_data_valid;
	wire [31:0] _argRouteRvm_15_io_read_data_bits;
	wire _argRouteRvm_15_io_write_address_ready;
	wire _argRouteRvm_15_io_write_data_ready;
	wire _argRouteRvm_14_io_read_address_ready;
	wire _argRouteRvm_14_io_read_data_valid;
	wire [31:0] _argRouteRvm_14_io_read_data_bits;
	wire _argRouteRvm_14_io_write_address_ready;
	wire _argRouteRvm_14_io_write_data_ready;
	wire _argRouteRvm_13_io_read_address_ready;
	wire _argRouteRvm_13_io_read_data_valid;
	wire [31:0] _argRouteRvm_13_io_read_data_bits;
	wire _argRouteRvm_13_io_write_address_ready;
	wire _argRouteRvm_13_io_write_data_ready;
	wire _argRouteRvm_12_io_read_address_ready;
	wire _argRouteRvm_12_io_read_data_valid;
	wire [31:0] _argRouteRvm_12_io_read_data_bits;
	wire _argRouteRvm_12_io_write_address_ready;
	wire _argRouteRvm_12_io_write_data_ready;
	wire _argRouteRvm_11_io_read_address_ready;
	wire _argRouteRvm_11_io_read_data_valid;
	wire [31:0] _argRouteRvm_11_io_read_data_bits;
	wire _argRouteRvm_11_io_write_address_ready;
	wire _argRouteRvm_11_io_write_data_ready;
	wire _argRouteRvm_10_io_read_address_ready;
	wire _argRouteRvm_10_io_read_data_valid;
	wire [31:0] _argRouteRvm_10_io_read_data_bits;
	wire _argRouteRvm_10_io_write_address_ready;
	wire _argRouteRvm_10_io_write_data_ready;
	wire _argRouteRvm_9_io_read_address_ready;
	wire _argRouteRvm_9_io_read_data_valid;
	wire [31:0] _argRouteRvm_9_io_read_data_bits;
	wire _argRouteRvm_9_io_write_address_ready;
	wire _argRouteRvm_9_io_write_data_ready;
	wire _argRouteRvm_8_io_read_address_ready;
	wire _argRouteRvm_8_io_read_data_valid;
	wire [31:0] _argRouteRvm_8_io_read_data_bits;
	wire _argRouteRvm_8_io_write_address_ready;
	wire _argRouteRvm_8_io_write_data_ready;
	wire _argRouteRvm_7_io_read_address_ready;
	wire _argRouteRvm_7_io_read_data_valid;
	wire [31:0] _argRouteRvm_7_io_read_data_bits;
	wire _argRouteRvm_7_io_write_address_ready;
	wire _argRouteRvm_7_io_write_data_ready;
	wire _argRouteRvm_6_io_read_address_ready;
	wire _argRouteRvm_6_io_read_data_valid;
	wire [31:0] _argRouteRvm_6_io_read_data_bits;
	wire _argRouteRvm_6_io_write_address_ready;
	wire _argRouteRvm_6_io_write_data_ready;
	wire _argRouteRvm_5_io_read_address_ready;
	wire _argRouteRvm_5_io_read_data_valid;
	wire [31:0] _argRouteRvm_5_io_read_data_bits;
	wire _argRouteRvm_5_io_write_address_ready;
	wire _argRouteRvm_5_io_write_data_ready;
	wire _argRouteRvm_4_io_read_address_ready;
	wire _argRouteRvm_4_io_read_data_valid;
	wire [31:0] _argRouteRvm_4_io_read_data_bits;
	wire _argRouteRvm_4_io_write_address_ready;
	wire _argRouteRvm_4_io_write_data_ready;
	wire _argRouteRvm_3_io_read_address_ready;
	wire _argRouteRvm_3_io_read_data_valid;
	wire [31:0] _argRouteRvm_3_io_read_data_bits;
	wire _argRouteRvm_3_io_write_address_ready;
	wire _argRouteRvm_3_io_write_data_ready;
	wire _argRouteRvm_2_io_read_address_ready;
	wire _argRouteRvm_2_io_read_data_valid;
	wire [31:0] _argRouteRvm_2_io_read_data_bits;
	wire _argRouteRvm_2_io_write_address_ready;
	wire _argRouteRvm_2_io_write_data_ready;
	wire _argRouteRvm_1_io_read_address_ready;
	wire _argRouteRvm_1_io_read_data_valid;
	wire [31:0] _argRouteRvm_1_io_read_data_bits;
	wire _argRouteRvm_1_io_write_address_ready;
	wire _argRouteRvm_1_io_write_data_ready;
	wire _argRouteRvm_0_io_read_address_ready;
	wire _argRouteRvm_0_io_read_data_valid;
	wire [31:0] _argRouteRvm_0_io_read_data_bits;
	wire _argRouteRvm_0_io_write_address_ready;
	wire _argRouteRvm_0_io_write_data_ready;
	wire _argRouteServers_15_io_connNetwork_ready;
	wire _argRouteServers_15_io_read_address_valid;
	wire [63:0] _argRouteServers_15_io_read_address_bits;
	wire _argRouteServers_15_io_read_data_ready;
	wire _argRouteServers_15_io_write_address_valid;
	wire [63:0] _argRouteServers_15_io_write_address_bits;
	wire _argRouteServers_15_io_write_data_valid;
	wire [31:0] _argRouteServers_15_io_write_data_bits;
	wire _argRouteServers_15_io_read_address_task_valid;
	wire [63:0] _argRouteServers_15_io_read_address_task_bits;
	wire _argRouteServers_15_io_read_data_task_ready;
	wire _argRouteServers_14_io_connNetwork_ready;
	wire _argRouteServers_14_io_read_address_valid;
	wire [63:0] _argRouteServers_14_io_read_address_bits;
	wire _argRouteServers_14_io_read_data_ready;
	wire _argRouteServers_14_io_write_address_valid;
	wire [63:0] _argRouteServers_14_io_write_address_bits;
	wire _argRouteServers_14_io_write_data_valid;
	wire [31:0] _argRouteServers_14_io_write_data_bits;
	wire _argRouteServers_14_io_read_address_task_valid;
	wire [63:0] _argRouteServers_14_io_read_address_task_bits;
	wire _argRouteServers_14_io_read_data_task_ready;
	wire _argRouteServers_13_io_connNetwork_ready;
	wire _argRouteServers_13_io_read_address_valid;
	wire [63:0] _argRouteServers_13_io_read_address_bits;
	wire _argRouteServers_13_io_read_data_ready;
	wire _argRouteServers_13_io_write_address_valid;
	wire [63:0] _argRouteServers_13_io_write_address_bits;
	wire _argRouteServers_13_io_write_data_valid;
	wire [31:0] _argRouteServers_13_io_write_data_bits;
	wire _argRouteServers_13_io_read_address_task_valid;
	wire [63:0] _argRouteServers_13_io_read_address_task_bits;
	wire _argRouteServers_13_io_read_data_task_ready;
	wire _argRouteServers_12_io_connNetwork_ready;
	wire _argRouteServers_12_io_read_address_valid;
	wire [63:0] _argRouteServers_12_io_read_address_bits;
	wire _argRouteServers_12_io_read_data_ready;
	wire _argRouteServers_12_io_write_address_valid;
	wire [63:0] _argRouteServers_12_io_write_address_bits;
	wire _argRouteServers_12_io_write_data_valid;
	wire [31:0] _argRouteServers_12_io_write_data_bits;
	wire _argRouteServers_12_io_read_address_task_valid;
	wire [63:0] _argRouteServers_12_io_read_address_task_bits;
	wire _argRouteServers_12_io_read_data_task_ready;
	wire _argRouteServers_11_io_connNetwork_ready;
	wire _argRouteServers_11_io_read_address_valid;
	wire [63:0] _argRouteServers_11_io_read_address_bits;
	wire _argRouteServers_11_io_read_data_ready;
	wire _argRouteServers_11_io_write_address_valid;
	wire [63:0] _argRouteServers_11_io_write_address_bits;
	wire _argRouteServers_11_io_write_data_valid;
	wire [31:0] _argRouteServers_11_io_write_data_bits;
	wire _argRouteServers_11_io_read_address_task_valid;
	wire [63:0] _argRouteServers_11_io_read_address_task_bits;
	wire _argRouteServers_11_io_read_data_task_ready;
	wire _argRouteServers_10_io_connNetwork_ready;
	wire _argRouteServers_10_io_read_address_valid;
	wire [63:0] _argRouteServers_10_io_read_address_bits;
	wire _argRouteServers_10_io_read_data_ready;
	wire _argRouteServers_10_io_write_address_valid;
	wire [63:0] _argRouteServers_10_io_write_address_bits;
	wire _argRouteServers_10_io_write_data_valid;
	wire [31:0] _argRouteServers_10_io_write_data_bits;
	wire _argRouteServers_10_io_read_address_task_valid;
	wire [63:0] _argRouteServers_10_io_read_address_task_bits;
	wire _argRouteServers_10_io_read_data_task_ready;
	wire _argRouteServers_9_io_connNetwork_ready;
	wire _argRouteServers_9_io_read_address_valid;
	wire [63:0] _argRouteServers_9_io_read_address_bits;
	wire _argRouteServers_9_io_read_data_ready;
	wire _argRouteServers_9_io_write_address_valid;
	wire [63:0] _argRouteServers_9_io_write_address_bits;
	wire _argRouteServers_9_io_write_data_valid;
	wire [31:0] _argRouteServers_9_io_write_data_bits;
	wire _argRouteServers_9_io_read_address_task_valid;
	wire [63:0] _argRouteServers_9_io_read_address_task_bits;
	wire _argRouteServers_9_io_read_data_task_ready;
	wire _argRouteServers_8_io_connNetwork_ready;
	wire _argRouteServers_8_io_read_address_valid;
	wire [63:0] _argRouteServers_8_io_read_address_bits;
	wire _argRouteServers_8_io_read_data_ready;
	wire _argRouteServers_8_io_write_address_valid;
	wire [63:0] _argRouteServers_8_io_write_address_bits;
	wire _argRouteServers_8_io_write_data_valid;
	wire [31:0] _argRouteServers_8_io_write_data_bits;
	wire _argRouteServers_8_io_read_address_task_valid;
	wire [63:0] _argRouteServers_8_io_read_address_task_bits;
	wire _argRouteServers_8_io_read_data_task_ready;
	wire _argRouteServers_7_io_connNetwork_ready;
	wire _argRouteServers_7_io_read_address_valid;
	wire [63:0] _argRouteServers_7_io_read_address_bits;
	wire _argRouteServers_7_io_read_data_ready;
	wire _argRouteServers_7_io_write_address_valid;
	wire [63:0] _argRouteServers_7_io_write_address_bits;
	wire _argRouteServers_7_io_write_data_valid;
	wire [31:0] _argRouteServers_7_io_write_data_bits;
	wire _argRouteServers_7_io_read_address_task_valid;
	wire [63:0] _argRouteServers_7_io_read_address_task_bits;
	wire _argRouteServers_7_io_read_data_task_ready;
	wire _argRouteServers_6_io_connNetwork_ready;
	wire _argRouteServers_6_io_read_address_valid;
	wire [63:0] _argRouteServers_6_io_read_address_bits;
	wire _argRouteServers_6_io_read_data_ready;
	wire _argRouteServers_6_io_write_address_valid;
	wire [63:0] _argRouteServers_6_io_write_address_bits;
	wire _argRouteServers_6_io_write_data_valid;
	wire [31:0] _argRouteServers_6_io_write_data_bits;
	wire _argRouteServers_6_io_read_address_task_valid;
	wire [63:0] _argRouteServers_6_io_read_address_task_bits;
	wire _argRouteServers_6_io_read_data_task_ready;
	wire _argRouteServers_5_io_connNetwork_ready;
	wire _argRouteServers_5_io_read_address_valid;
	wire [63:0] _argRouteServers_5_io_read_address_bits;
	wire _argRouteServers_5_io_read_data_ready;
	wire _argRouteServers_5_io_write_address_valid;
	wire [63:0] _argRouteServers_5_io_write_address_bits;
	wire _argRouteServers_5_io_write_data_valid;
	wire [31:0] _argRouteServers_5_io_write_data_bits;
	wire _argRouteServers_5_io_read_address_task_valid;
	wire [63:0] _argRouteServers_5_io_read_address_task_bits;
	wire _argRouteServers_5_io_read_data_task_ready;
	wire _argRouteServers_4_io_connNetwork_ready;
	wire _argRouteServers_4_io_read_address_valid;
	wire [63:0] _argRouteServers_4_io_read_address_bits;
	wire _argRouteServers_4_io_read_data_ready;
	wire _argRouteServers_4_io_write_address_valid;
	wire [63:0] _argRouteServers_4_io_write_address_bits;
	wire _argRouteServers_4_io_write_data_valid;
	wire [31:0] _argRouteServers_4_io_write_data_bits;
	wire _argRouteServers_4_io_read_address_task_valid;
	wire [63:0] _argRouteServers_4_io_read_address_task_bits;
	wire _argRouteServers_4_io_read_data_task_ready;
	wire _argRouteServers_3_io_connNetwork_ready;
	wire _argRouteServers_3_io_read_address_valid;
	wire [63:0] _argRouteServers_3_io_read_address_bits;
	wire _argRouteServers_3_io_read_data_ready;
	wire _argRouteServers_3_io_write_address_valid;
	wire [63:0] _argRouteServers_3_io_write_address_bits;
	wire _argRouteServers_3_io_write_data_valid;
	wire [31:0] _argRouteServers_3_io_write_data_bits;
	wire _argRouteServers_3_io_read_address_task_valid;
	wire [63:0] _argRouteServers_3_io_read_address_task_bits;
	wire _argRouteServers_3_io_read_data_task_ready;
	wire _argRouteServers_2_io_connNetwork_ready;
	wire _argRouteServers_2_io_read_address_valid;
	wire [63:0] _argRouteServers_2_io_read_address_bits;
	wire _argRouteServers_2_io_read_data_ready;
	wire _argRouteServers_2_io_write_address_valid;
	wire [63:0] _argRouteServers_2_io_write_address_bits;
	wire _argRouteServers_2_io_write_data_valid;
	wire [31:0] _argRouteServers_2_io_write_data_bits;
	wire _argRouteServers_2_io_read_address_task_valid;
	wire [63:0] _argRouteServers_2_io_read_address_task_bits;
	wire _argRouteServers_2_io_read_data_task_ready;
	wire _argRouteServers_1_io_connNetwork_ready;
	wire _argRouteServers_1_io_read_address_valid;
	wire [63:0] _argRouteServers_1_io_read_address_bits;
	wire _argRouteServers_1_io_read_data_ready;
	wire _argRouteServers_1_io_write_address_valid;
	wire [63:0] _argRouteServers_1_io_write_address_bits;
	wire _argRouteServers_1_io_write_data_valid;
	wire [31:0] _argRouteServers_1_io_write_data_bits;
	wire _argRouteServers_1_io_read_address_task_valid;
	wire [63:0] _argRouteServers_1_io_read_address_task_bits;
	wire _argRouteServers_1_io_read_data_task_ready;
	wire _argRouteServers_0_io_connNetwork_ready;
	wire _argRouteServers_0_io_read_address_valid;
	wire [63:0] _argRouteServers_0_io_read_address_bits;
	wire _argRouteServers_0_io_read_data_ready;
	wire _argRouteServers_0_io_write_address_valid;
	wire [63:0] _argRouteServers_0_io_write_address_bits;
	wire _argRouteServers_0_io_write_data_valid;
	wire [31:0] _argRouteServers_0_io_write_data_bits;
	wire _argRouteServers_0_io_read_address_task_valid;
	wire [63:0] _argRouteServers_0_io_read_address_task_bits;
	wire _argRouteServers_0_io_read_data_task_ready;
	wire _argSide_io_connVAS_0_valid;
	wire [63:0] _argSide_io_connVAS_0_bits;
	wire _argSide_io_connVAS_1_valid;
	wire [63:0] _argSide_io_connVAS_1_bits;
	wire _argSide_io_connVAS_2_valid;
	wire [63:0] _argSide_io_connVAS_2_bits;
	wire _argSide_io_connVAS_3_valid;
	wire [63:0] _argSide_io_connVAS_3_bits;
	wire _argSide_io_connVAS_4_valid;
	wire [63:0] _argSide_io_connVAS_4_bits;
	wire _argSide_io_connVAS_5_valid;
	wire [63:0] _argSide_io_connVAS_5_bits;
	wire _argSide_io_connVAS_6_valid;
	wire [63:0] _argSide_io_connVAS_6_bits;
	wire _argSide_io_connVAS_7_valid;
	wire [63:0] _argSide_io_connVAS_7_bits;
	wire _argSide_io_connVAS_8_valid;
	wire [63:0] _argSide_io_connVAS_8_bits;
	wire _argSide_io_connVAS_9_valid;
	wire [63:0] _argSide_io_connVAS_9_bits;
	wire _argSide_io_connVAS_10_valid;
	wire [63:0] _argSide_io_connVAS_10_bits;
	wire _argSide_io_connVAS_11_valid;
	wire [63:0] _argSide_io_connVAS_11_bits;
	wire _argSide_io_connVAS_12_valid;
	wire [63:0] _argSide_io_connVAS_12_bits;
	wire _argSide_io_connVAS_13_valid;
	wire [63:0] _argSide_io_connVAS_13_bits;
	wire _argSide_io_connVAS_14_valid;
	wire [63:0] _argSide_io_connVAS_14_bits;
	wire _argSide_io_connVAS_15_valid;
	wire [63:0] _argSide_io_connVAS_15_bits;
	wire _argSide_io_connPE_0_ready;
	wire _argSide_io_connPE_1_ready;
	wire _argSide_io_connPE_2_ready;
	wire _argSide_io_connPE_3_ready;
	wire _argSide_io_connPE_4_ready;
	wire _argSide_io_connPE_5_ready;
	wire _argSide_io_connPE_6_ready;
	wire _argSide_io_connPE_7_ready;
	wire _argSide_io_connPE_8_ready;
	wire _argSide_io_connPE_9_ready;
	wire _argSide_io_connPE_10_ready;
	wire _argSide_io_connPE_11_ready;
	wire _argSide_io_connPE_12_ready;
	wire _argSide_io_connPE_13_ready;
	wire _argSide_io_connPE_14_ready;
	wire _argSide_io_connPE_15_ready;
	wire _argSide_io_connPE_16_ready;
	wire _argSide_io_connPE_17_ready;
	wire _argSide_io_connPE_18_ready;
	wire _argSide_io_connPE_19_ready;
	wire _argSide_io_connPE_20_ready;
	wire _argSide_io_connPE_21_ready;
	wire _argSide_io_connPE_22_ready;
	wire _argSide_io_connPE_23_ready;
	wire _argSide_io_connPE_24_ready;
	wire _argSide_io_connPE_25_ready;
	wire _argSide_io_connPE_26_ready;
	wire _argSide_io_connPE_27_ready;
	wire _argSide_io_connPE_28_ready;
	wire _argSide_io_connPE_29_ready;
	wire _argSide_io_connPE_30_ready;
	wire _argSide_io_connPE_31_ready;
	wire _argSide_io_connPE_32_ready;
	wire _argSide_io_connPE_33_ready;
	wire _argSide_io_connPE_34_ready;
	wire _argSide_io_connPE_35_ready;
	wire _argSide_io_connPE_36_ready;
	wire _argSide_io_connPE_37_ready;
	wire _argSide_io_connPE_38_ready;
	wire _argSide_io_connPE_39_ready;
	wire _argSide_io_connPE_40_ready;
	wire _argSide_io_connPE_41_ready;
	wire _argSide_io_connPE_42_ready;
	wire _argSide_io_connPE_43_ready;
	wire _argSide_io_connPE_44_ready;
	wire _argSide_io_connPE_45_ready;
	wire _argSide_io_connPE_46_ready;
	wire _argSide_io_connPE_47_ready;
	wire _argSide_io_connPE_48_ready;
	wire _argSide_io_connPE_49_ready;
	wire _argSide_io_connPE_50_ready;
	wire _argSide_io_connPE_51_ready;
	wire _argSide_io_connPE_52_ready;
	wire _argSide_io_connPE_53_ready;
	wire _argSide_io_connPE_54_ready;
	wire _argSide_io_connPE_55_ready;
	wire _argSide_io_connPE_56_ready;
	wire _argSide_io_connPE_57_ready;
	wire _argSide_io_connPE_58_ready;
	wire _argSide_io_connPE_59_ready;
	wire _argSide_io_connPE_60_ready;
	wire _argSide_io_connPE_61_ready;
	wire _argSide_io_connPE_62_ready;
	wire _argSide_io_connPE_63_ready;
	wire _argSide_io_connPE_64_ready;
	wire _argSide_io_connPE_65_ready;
	wire _argSide_io_connPE_66_ready;
	wire _argSide_io_connPE_67_ready;
	wire _argSide_io_connPE_68_ready;
	wire _argSide_io_connPE_69_ready;
	wire _argSide_io_connPE_70_ready;
	wire _argSide_io_connPE_71_ready;
	wire _argSide_io_connPE_72_ready;
	wire _argSide_io_connPE_73_ready;
	wire _argSide_io_connPE_74_ready;
	wire _argSide_io_connPE_75_ready;
	wire _argSide_io_connPE_76_ready;
	wire _argSide_io_connPE_77_ready;
	wire _argSide_io_connPE_78_ready;
	wire _argSide_io_connPE_79_ready;
	ArgumentNotifierNetwork argSide(
		.clock(clock),
		.reset(reset),
		.io_connVAS_0_ready(_argRouteServers_0_io_connNetwork_ready),
		.io_connVAS_0_valid(_argSide_io_connVAS_0_valid),
		.io_connVAS_0_bits(_argSide_io_connVAS_0_bits),
		.io_connVAS_1_ready(_argRouteServers_1_io_connNetwork_ready),
		.io_connVAS_1_valid(_argSide_io_connVAS_1_valid),
		.io_connVAS_1_bits(_argSide_io_connVAS_1_bits),
		.io_connVAS_2_ready(_argRouteServers_2_io_connNetwork_ready),
		.io_connVAS_2_valid(_argSide_io_connVAS_2_valid),
		.io_connVAS_2_bits(_argSide_io_connVAS_2_bits),
		.io_connVAS_3_ready(_argRouteServers_3_io_connNetwork_ready),
		.io_connVAS_3_valid(_argSide_io_connVAS_3_valid),
		.io_connVAS_3_bits(_argSide_io_connVAS_3_bits),
		.io_connVAS_4_ready(_argRouteServers_4_io_connNetwork_ready),
		.io_connVAS_4_valid(_argSide_io_connVAS_4_valid),
		.io_connVAS_4_bits(_argSide_io_connVAS_4_bits),
		.io_connVAS_5_ready(_argRouteServers_5_io_connNetwork_ready),
		.io_connVAS_5_valid(_argSide_io_connVAS_5_valid),
		.io_connVAS_5_bits(_argSide_io_connVAS_5_bits),
		.io_connVAS_6_ready(_argRouteServers_6_io_connNetwork_ready),
		.io_connVAS_6_valid(_argSide_io_connVAS_6_valid),
		.io_connVAS_6_bits(_argSide_io_connVAS_6_bits),
		.io_connVAS_7_ready(_argRouteServers_7_io_connNetwork_ready),
		.io_connVAS_7_valid(_argSide_io_connVAS_7_valid),
		.io_connVAS_7_bits(_argSide_io_connVAS_7_bits),
		.io_connVAS_8_ready(_argRouteServers_8_io_connNetwork_ready),
		.io_connVAS_8_valid(_argSide_io_connVAS_8_valid),
		.io_connVAS_8_bits(_argSide_io_connVAS_8_bits),
		.io_connVAS_9_ready(_argRouteServers_9_io_connNetwork_ready),
		.io_connVAS_9_valid(_argSide_io_connVAS_9_valid),
		.io_connVAS_9_bits(_argSide_io_connVAS_9_bits),
		.io_connVAS_10_ready(_argRouteServers_10_io_connNetwork_ready),
		.io_connVAS_10_valid(_argSide_io_connVAS_10_valid),
		.io_connVAS_10_bits(_argSide_io_connVAS_10_bits),
		.io_connVAS_11_ready(_argRouteServers_11_io_connNetwork_ready),
		.io_connVAS_11_valid(_argSide_io_connVAS_11_valid),
		.io_connVAS_11_bits(_argSide_io_connVAS_11_bits),
		.io_connVAS_12_ready(_argRouteServers_12_io_connNetwork_ready),
		.io_connVAS_12_valid(_argSide_io_connVAS_12_valid),
		.io_connVAS_12_bits(_argSide_io_connVAS_12_bits),
		.io_connVAS_13_ready(_argRouteServers_13_io_connNetwork_ready),
		.io_connVAS_13_valid(_argSide_io_connVAS_13_valid),
		.io_connVAS_13_bits(_argSide_io_connVAS_13_bits),
		.io_connVAS_14_ready(_argRouteServers_14_io_connNetwork_ready),
		.io_connVAS_14_valid(_argSide_io_connVAS_14_valid),
		.io_connVAS_14_bits(_argSide_io_connVAS_14_bits),
		.io_connVAS_15_ready(_argRouteServers_15_io_connNetwork_ready),
		.io_connVAS_15_valid(_argSide_io_connVAS_15_valid),
		.io_connVAS_15_bits(_argSide_io_connVAS_15_bits),
		.io_connPE_0_ready(_argSide_io_connPE_0_ready),
		.io_connPE_0_valid(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_connPE_0_bits(_axis_stream_converters_in_0_io_dataOut_TDATA),
		.io_connPE_1_ready(_argSide_io_connPE_1_ready),
		.io_connPE_1_valid(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_connPE_1_bits(_axis_stream_converters_in_1_io_dataOut_TDATA),
		.io_connPE_2_ready(_argSide_io_connPE_2_ready),
		.io_connPE_2_valid(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_connPE_2_bits(_axis_stream_converters_in_2_io_dataOut_TDATA),
		.io_connPE_3_ready(_argSide_io_connPE_3_ready),
		.io_connPE_3_valid(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_connPE_3_bits(_axis_stream_converters_in_3_io_dataOut_TDATA),
		.io_connPE_4_ready(_argSide_io_connPE_4_ready),
		.io_connPE_4_valid(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_connPE_4_bits(_axis_stream_converters_in_4_io_dataOut_TDATA),
		.io_connPE_5_ready(_argSide_io_connPE_5_ready),
		.io_connPE_5_valid(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_connPE_5_bits(_axis_stream_converters_in_5_io_dataOut_TDATA),
		.io_connPE_6_ready(_argSide_io_connPE_6_ready),
		.io_connPE_6_valid(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_connPE_6_bits(_axis_stream_converters_in_6_io_dataOut_TDATA),
		.io_connPE_7_ready(_argSide_io_connPE_7_ready),
		.io_connPE_7_valid(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_connPE_7_bits(_axis_stream_converters_in_7_io_dataOut_TDATA),
		.io_connPE_8_ready(_argSide_io_connPE_8_ready),
		.io_connPE_8_valid(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_connPE_8_bits(_axis_stream_converters_in_8_io_dataOut_TDATA),
		.io_connPE_9_ready(_argSide_io_connPE_9_ready),
		.io_connPE_9_valid(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_connPE_9_bits(_axis_stream_converters_in_9_io_dataOut_TDATA),
		.io_connPE_10_ready(_argSide_io_connPE_10_ready),
		.io_connPE_10_valid(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_connPE_10_bits(_axis_stream_converters_in_10_io_dataOut_TDATA),
		.io_connPE_11_ready(_argSide_io_connPE_11_ready),
		.io_connPE_11_valid(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_connPE_11_bits(_axis_stream_converters_in_11_io_dataOut_TDATA),
		.io_connPE_12_ready(_argSide_io_connPE_12_ready),
		.io_connPE_12_valid(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_connPE_12_bits(_axis_stream_converters_in_12_io_dataOut_TDATA),
		.io_connPE_13_ready(_argSide_io_connPE_13_ready),
		.io_connPE_13_valid(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_connPE_13_bits(_axis_stream_converters_in_13_io_dataOut_TDATA),
		.io_connPE_14_ready(_argSide_io_connPE_14_ready),
		.io_connPE_14_valid(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_connPE_14_bits(_axis_stream_converters_in_14_io_dataOut_TDATA),
		.io_connPE_15_ready(_argSide_io_connPE_15_ready),
		.io_connPE_15_valid(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_connPE_15_bits(_axis_stream_converters_in_15_io_dataOut_TDATA),
		.io_connPE_16_ready(_argSide_io_connPE_16_ready),
		.io_connPE_16_valid(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_connPE_16_bits(_axis_stream_converters_in_16_io_dataOut_TDATA),
		.io_connPE_17_ready(_argSide_io_connPE_17_ready),
		.io_connPE_17_valid(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_connPE_17_bits(_axis_stream_converters_in_17_io_dataOut_TDATA),
		.io_connPE_18_ready(_argSide_io_connPE_18_ready),
		.io_connPE_18_valid(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_connPE_18_bits(_axis_stream_converters_in_18_io_dataOut_TDATA),
		.io_connPE_19_ready(_argSide_io_connPE_19_ready),
		.io_connPE_19_valid(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_connPE_19_bits(_axis_stream_converters_in_19_io_dataOut_TDATA),
		.io_connPE_20_ready(_argSide_io_connPE_20_ready),
		.io_connPE_20_valid(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_connPE_20_bits(_axis_stream_converters_in_20_io_dataOut_TDATA),
		.io_connPE_21_ready(_argSide_io_connPE_21_ready),
		.io_connPE_21_valid(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_connPE_21_bits(_axis_stream_converters_in_21_io_dataOut_TDATA),
		.io_connPE_22_ready(_argSide_io_connPE_22_ready),
		.io_connPE_22_valid(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_connPE_22_bits(_axis_stream_converters_in_22_io_dataOut_TDATA),
		.io_connPE_23_ready(_argSide_io_connPE_23_ready),
		.io_connPE_23_valid(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_connPE_23_bits(_axis_stream_converters_in_23_io_dataOut_TDATA),
		.io_connPE_24_ready(_argSide_io_connPE_24_ready),
		.io_connPE_24_valid(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_connPE_24_bits(_axis_stream_converters_in_24_io_dataOut_TDATA),
		.io_connPE_25_ready(_argSide_io_connPE_25_ready),
		.io_connPE_25_valid(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_connPE_25_bits(_axis_stream_converters_in_25_io_dataOut_TDATA),
		.io_connPE_26_ready(_argSide_io_connPE_26_ready),
		.io_connPE_26_valid(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_connPE_26_bits(_axis_stream_converters_in_26_io_dataOut_TDATA),
		.io_connPE_27_ready(_argSide_io_connPE_27_ready),
		.io_connPE_27_valid(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_connPE_27_bits(_axis_stream_converters_in_27_io_dataOut_TDATA),
		.io_connPE_28_ready(_argSide_io_connPE_28_ready),
		.io_connPE_28_valid(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_connPE_28_bits(_axis_stream_converters_in_28_io_dataOut_TDATA),
		.io_connPE_29_ready(_argSide_io_connPE_29_ready),
		.io_connPE_29_valid(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_connPE_29_bits(_axis_stream_converters_in_29_io_dataOut_TDATA),
		.io_connPE_30_ready(_argSide_io_connPE_30_ready),
		.io_connPE_30_valid(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_connPE_30_bits(_axis_stream_converters_in_30_io_dataOut_TDATA),
		.io_connPE_31_ready(_argSide_io_connPE_31_ready),
		.io_connPE_31_valid(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_connPE_31_bits(_axis_stream_converters_in_31_io_dataOut_TDATA),
		.io_connPE_32_ready(_argSide_io_connPE_32_ready),
		.io_connPE_32_valid(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_connPE_32_bits(_axis_stream_converters_in_32_io_dataOut_TDATA),
		.io_connPE_33_ready(_argSide_io_connPE_33_ready),
		.io_connPE_33_valid(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_connPE_33_bits(_axis_stream_converters_in_33_io_dataOut_TDATA),
		.io_connPE_34_ready(_argSide_io_connPE_34_ready),
		.io_connPE_34_valid(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_connPE_34_bits(_axis_stream_converters_in_34_io_dataOut_TDATA),
		.io_connPE_35_ready(_argSide_io_connPE_35_ready),
		.io_connPE_35_valid(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_connPE_35_bits(_axis_stream_converters_in_35_io_dataOut_TDATA),
		.io_connPE_36_ready(_argSide_io_connPE_36_ready),
		.io_connPE_36_valid(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_connPE_36_bits(_axis_stream_converters_in_36_io_dataOut_TDATA),
		.io_connPE_37_ready(_argSide_io_connPE_37_ready),
		.io_connPE_37_valid(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_connPE_37_bits(_axis_stream_converters_in_37_io_dataOut_TDATA),
		.io_connPE_38_ready(_argSide_io_connPE_38_ready),
		.io_connPE_38_valid(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_connPE_38_bits(_axis_stream_converters_in_38_io_dataOut_TDATA),
		.io_connPE_39_ready(_argSide_io_connPE_39_ready),
		.io_connPE_39_valid(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_connPE_39_bits(_axis_stream_converters_in_39_io_dataOut_TDATA),
		.io_connPE_40_ready(_argSide_io_connPE_40_ready),
		.io_connPE_40_valid(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_connPE_40_bits(_axis_stream_converters_in_40_io_dataOut_TDATA),
		.io_connPE_41_ready(_argSide_io_connPE_41_ready),
		.io_connPE_41_valid(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_connPE_41_bits(_axis_stream_converters_in_41_io_dataOut_TDATA),
		.io_connPE_42_ready(_argSide_io_connPE_42_ready),
		.io_connPE_42_valid(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_connPE_42_bits(_axis_stream_converters_in_42_io_dataOut_TDATA),
		.io_connPE_43_ready(_argSide_io_connPE_43_ready),
		.io_connPE_43_valid(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_connPE_43_bits(_axis_stream_converters_in_43_io_dataOut_TDATA),
		.io_connPE_44_ready(_argSide_io_connPE_44_ready),
		.io_connPE_44_valid(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_connPE_44_bits(_axis_stream_converters_in_44_io_dataOut_TDATA),
		.io_connPE_45_ready(_argSide_io_connPE_45_ready),
		.io_connPE_45_valid(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_connPE_45_bits(_axis_stream_converters_in_45_io_dataOut_TDATA),
		.io_connPE_46_ready(_argSide_io_connPE_46_ready),
		.io_connPE_46_valid(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_connPE_46_bits(_axis_stream_converters_in_46_io_dataOut_TDATA),
		.io_connPE_47_ready(_argSide_io_connPE_47_ready),
		.io_connPE_47_valid(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_connPE_47_bits(_axis_stream_converters_in_47_io_dataOut_TDATA),
		.io_connPE_48_ready(_argSide_io_connPE_48_ready),
		.io_connPE_48_valid(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_connPE_48_bits(_axis_stream_converters_in_48_io_dataOut_TDATA),
		.io_connPE_49_ready(_argSide_io_connPE_49_ready),
		.io_connPE_49_valid(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_connPE_49_bits(_axis_stream_converters_in_49_io_dataOut_TDATA),
		.io_connPE_50_ready(_argSide_io_connPE_50_ready),
		.io_connPE_50_valid(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_connPE_50_bits(_axis_stream_converters_in_50_io_dataOut_TDATA),
		.io_connPE_51_ready(_argSide_io_connPE_51_ready),
		.io_connPE_51_valid(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_connPE_51_bits(_axis_stream_converters_in_51_io_dataOut_TDATA),
		.io_connPE_52_ready(_argSide_io_connPE_52_ready),
		.io_connPE_52_valid(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_connPE_52_bits(_axis_stream_converters_in_52_io_dataOut_TDATA),
		.io_connPE_53_ready(_argSide_io_connPE_53_ready),
		.io_connPE_53_valid(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_connPE_53_bits(_axis_stream_converters_in_53_io_dataOut_TDATA),
		.io_connPE_54_ready(_argSide_io_connPE_54_ready),
		.io_connPE_54_valid(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_connPE_54_bits(_axis_stream_converters_in_54_io_dataOut_TDATA),
		.io_connPE_55_ready(_argSide_io_connPE_55_ready),
		.io_connPE_55_valid(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_connPE_55_bits(_axis_stream_converters_in_55_io_dataOut_TDATA),
		.io_connPE_56_ready(_argSide_io_connPE_56_ready),
		.io_connPE_56_valid(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_connPE_56_bits(_axis_stream_converters_in_56_io_dataOut_TDATA),
		.io_connPE_57_ready(_argSide_io_connPE_57_ready),
		.io_connPE_57_valid(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_connPE_57_bits(_axis_stream_converters_in_57_io_dataOut_TDATA),
		.io_connPE_58_ready(_argSide_io_connPE_58_ready),
		.io_connPE_58_valid(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_connPE_58_bits(_axis_stream_converters_in_58_io_dataOut_TDATA),
		.io_connPE_59_ready(_argSide_io_connPE_59_ready),
		.io_connPE_59_valid(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_connPE_59_bits(_axis_stream_converters_in_59_io_dataOut_TDATA),
		.io_connPE_60_ready(_argSide_io_connPE_60_ready),
		.io_connPE_60_valid(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_connPE_60_bits(_axis_stream_converters_in_60_io_dataOut_TDATA),
		.io_connPE_61_ready(_argSide_io_connPE_61_ready),
		.io_connPE_61_valid(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_connPE_61_bits(_axis_stream_converters_in_61_io_dataOut_TDATA),
		.io_connPE_62_ready(_argSide_io_connPE_62_ready),
		.io_connPE_62_valid(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_connPE_62_bits(_axis_stream_converters_in_62_io_dataOut_TDATA),
		.io_connPE_63_ready(_argSide_io_connPE_63_ready),
		.io_connPE_63_valid(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_connPE_63_bits(_axis_stream_converters_in_63_io_dataOut_TDATA),
		.io_connPE_64_ready(_argSide_io_connPE_64_ready),
		.io_connPE_64_valid(_axis_stream_converters_in_64_io_dataOut_TVALID),
		.io_connPE_64_bits(_axis_stream_converters_in_64_io_dataOut_TDATA),
		.io_connPE_65_ready(_argSide_io_connPE_65_ready),
		.io_connPE_65_valid(_axis_stream_converters_in_65_io_dataOut_TVALID),
		.io_connPE_65_bits(_axis_stream_converters_in_65_io_dataOut_TDATA),
		.io_connPE_66_ready(_argSide_io_connPE_66_ready),
		.io_connPE_66_valid(_axis_stream_converters_in_66_io_dataOut_TVALID),
		.io_connPE_66_bits(_axis_stream_converters_in_66_io_dataOut_TDATA),
		.io_connPE_67_ready(_argSide_io_connPE_67_ready),
		.io_connPE_67_valid(_axis_stream_converters_in_67_io_dataOut_TVALID),
		.io_connPE_67_bits(_axis_stream_converters_in_67_io_dataOut_TDATA),
		.io_connPE_68_ready(_argSide_io_connPE_68_ready),
		.io_connPE_68_valid(_axis_stream_converters_in_68_io_dataOut_TVALID),
		.io_connPE_68_bits(_axis_stream_converters_in_68_io_dataOut_TDATA),
		.io_connPE_69_ready(_argSide_io_connPE_69_ready),
		.io_connPE_69_valid(_axis_stream_converters_in_69_io_dataOut_TVALID),
		.io_connPE_69_bits(_axis_stream_converters_in_69_io_dataOut_TDATA),
		.io_connPE_70_ready(_argSide_io_connPE_70_ready),
		.io_connPE_70_valid(_axis_stream_converters_in_70_io_dataOut_TVALID),
		.io_connPE_70_bits(_axis_stream_converters_in_70_io_dataOut_TDATA),
		.io_connPE_71_ready(_argSide_io_connPE_71_ready),
		.io_connPE_71_valid(_axis_stream_converters_in_71_io_dataOut_TVALID),
		.io_connPE_71_bits(_axis_stream_converters_in_71_io_dataOut_TDATA),
		.io_connPE_72_ready(_argSide_io_connPE_72_ready),
		.io_connPE_72_valid(_axis_stream_converters_in_72_io_dataOut_TVALID),
		.io_connPE_72_bits(_axis_stream_converters_in_72_io_dataOut_TDATA),
		.io_connPE_73_ready(_argSide_io_connPE_73_ready),
		.io_connPE_73_valid(_axis_stream_converters_in_73_io_dataOut_TVALID),
		.io_connPE_73_bits(_axis_stream_converters_in_73_io_dataOut_TDATA),
		.io_connPE_74_ready(_argSide_io_connPE_74_ready),
		.io_connPE_74_valid(_axis_stream_converters_in_74_io_dataOut_TVALID),
		.io_connPE_74_bits(_axis_stream_converters_in_74_io_dataOut_TDATA),
		.io_connPE_75_ready(_argSide_io_connPE_75_ready),
		.io_connPE_75_valid(_axis_stream_converters_in_75_io_dataOut_TVALID),
		.io_connPE_75_bits(_axis_stream_converters_in_75_io_dataOut_TDATA),
		.io_connPE_76_ready(_argSide_io_connPE_76_ready),
		.io_connPE_76_valid(_axis_stream_converters_in_76_io_dataOut_TVALID),
		.io_connPE_76_bits(_axis_stream_converters_in_76_io_dataOut_TDATA),
		.io_connPE_77_ready(_argSide_io_connPE_77_ready),
		.io_connPE_77_valid(_axis_stream_converters_in_77_io_dataOut_TVALID),
		.io_connPE_77_bits(_axis_stream_converters_in_77_io_dataOut_TDATA),
		.io_connPE_78_ready(_argSide_io_connPE_78_ready),
		.io_connPE_78_valid(_axis_stream_converters_in_78_io_dataOut_TVALID),
		.io_connPE_78_bits(_axis_stream_converters_in_78_io_dataOut_TDATA),
		.io_connPE_79_ready(_argSide_io_connPE_79_ready),
		.io_connPE_79_valid(_axis_stream_converters_in_79_io_dataOut_TVALID),
		.io_connPE_79_bits(_axis_stream_converters_in_79_io_dataOut_TDATA)
	);
	ArgumentServer argRouteServers_0(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_0_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_0_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_0_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_0_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_0_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_0_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_0_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_0_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_0_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_0_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_0_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_0_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_0_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_0_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_0_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_0_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_0_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_0_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_0_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_0_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_0_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_0_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_0_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_0_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_0_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_0_io_read_data_bits)
	);
	ArgumentServer argRouteServers_1(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_1_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_1_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_1_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_1_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_1_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_1_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_1_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_1_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_1_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_1_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_1_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_1_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_1_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_1_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_1_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_1_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_1_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_1_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_1_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_1_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_1_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_1_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_1_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_1_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_1_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_1_io_read_data_bits)
	);
	ArgumentServer argRouteServers_2(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_2_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_2_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_2_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_2_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_2_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_2_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_2_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_2_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_2_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_2_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_2_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_2_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_2_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_2_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_2_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_2_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_2_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_2_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_2_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_2_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_2_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_2_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_2_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_2_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_2_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_2_io_read_data_bits)
	);
	ArgumentServer argRouteServers_3(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_3_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_3_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_3_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_3_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_3_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_3_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_3_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_3_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_3_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_3_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_3_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_3_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_3_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_3_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_3_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_3_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_3_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_3_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_3_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_3_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_3_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_3_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_3_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_3_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_3_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_3_io_read_data_bits)
	);
	ArgumentServer argRouteServers_4(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_4_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_4_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_4_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_4_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_4_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_4_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_4_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_4_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_4_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_4_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_4_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_4_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_4_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_4_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_4_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_4_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_4_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_4_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_4_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_4_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_4_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_4_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_4_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_4_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_4_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_4_io_read_data_bits)
	);
	ArgumentServer argRouteServers_5(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_5_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_5_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_5_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_5_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_5_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_5_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_5_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_5_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_5_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_5_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_5_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_5_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_5_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_5_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_5_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_5_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_5_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_5_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_5_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_5_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_5_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_5_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_5_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_5_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_5_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_5_io_read_data_bits)
	);
	ArgumentServer argRouteServers_6(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_6_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_6_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_6_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_6_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_6_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_6_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_6_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_6_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_6_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_6_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_6_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_6_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_6_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_6_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_6_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_6_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_6_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_6_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_6_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_6_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_6_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_6_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_6_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_6_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_6_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_6_io_read_data_bits)
	);
	ArgumentServer argRouteServers_7(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_7_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_7_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_7_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_7_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_7_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_7_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_7_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_7_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_7_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_7_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_7_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_7_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_7_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_7_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_7_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_7_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_7_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_7_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_7_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_7_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_7_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_7_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_7_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_7_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_7_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_7_io_read_data_bits)
	);
	ArgumentServer argRouteServers_8(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_8_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_8_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_8_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_8_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_8_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_8_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_8_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_8_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_8_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_8_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_8_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_8_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_8_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_8_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_8_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_8_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_8_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_8_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_8_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_8_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_8_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_8_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_8_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_8_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_8_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_8_io_read_data_bits)
	);
	ArgumentServer argRouteServers_9(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_9_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_9_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_9_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_9_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_9_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_9_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_9_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_9_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_9_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_9_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_9_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_9_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_9_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_9_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_9_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_9_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_9_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_9_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_9_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_9_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_9_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_9_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_9_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_9_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_9_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_9_io_read_data_bits)
	);
	ArgumentServer argRouteServers_10(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_10_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_10_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_10_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_10_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_10_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_10_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_10_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_10_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_10_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_10_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_10_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_10_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_10_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_10_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_10_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_10_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_10_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_10_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_10_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_10_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_10_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_10_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_10_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_10_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_10_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_10_io_read_data_bits)
	);
	ArgumentServer argRouteServers_11(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_11_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_11_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_11_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_11_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_11_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_11_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_11_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_11_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_11_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_11_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_11_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_11_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_11_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_11_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_11_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_11_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_11_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_11_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_11_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_11_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_11_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_11_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_11_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_11_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_11_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_11_io_read_data_bits)
	);
	ArgumentServer argRouteServers_12(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_12_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_12_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_12_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_12_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_12_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_12_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_12_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_12_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_12_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_12_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_12_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_12_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_12_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_12_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_12_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_12_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_12_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_12_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_12_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_12_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_12_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_12_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_12_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_12_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_12_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_12_io_read_data_bits)
	);
	ArgumentServer argRouteServers_13(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_13_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_13_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_13_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_13_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_13_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_13_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_13_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_13_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_13_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_13_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_13_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_13_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_13_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_13_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_13_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_13_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_13_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_13_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_13_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_13_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_13_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_13_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_13_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_13_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_13_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_13_io_read_data_bits)
	);
	ArgumentServer argRouteServers_14(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_14_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_14_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_14_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_14_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_14_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_14_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_14_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_14_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_14_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_14_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_14_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_14_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_14_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_14_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_14_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_14_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_14_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_14_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_14_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_14_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_14_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_14_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_14_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_14_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_14_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_14_io_read_data_bits)
	);
	ArgumentServer argRouteServers_15(
		.clock(clock),
		.reset(reset),
		.io_connNetwork_ready(_argRouteServers_15_io_connNetwork_ready),
		.io_connNetwork_valid(_argSide_io_connVAS_15_valid),
		.io_connNetwork_bits(_argSide_io_connVAS_15_bits),
		.io_connStealNtw_ctrl_serveStealReq_valid(connStealNtw_15_ctrl_serveStealReq_valid),
		.io_connStealNtw_ctrl_serveStealReq_ready(connStealNtw_15_ctrl_serveStealReq_ready),
		.io_connStealNtw_data_qOutTask_ready(connStealNtw_15_data_qOutTask_ready),
		.io_connStealNtw_data_qOutTask_valid(connStealNtw_15_data_qOutTask_valid),
		.io_connStealNtw_data_qOutTask_bits(connStealNtw_15_data_qOutTask_bits),
		.io_read_address_ready(_argRouteRvm_15_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_15_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_15_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_15_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_15_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_15_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_15_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_15_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_15_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_15_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_15_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_15_io_write_data_bits),
		.io_read_address_task_ready(_argRouteRvmReadOnly_15_io_read_address_ready),
		.io_read_address_task_valid(_argRouteServers_15_io_read_address_task_valid),
		.io_read_address_task_bits(_argRouteServers_15_io_read_address_task_bits),
		.io_read_data_task_ready(_argRouteServers_15_io_read_data_task_ready),
		.io_read_data_task_valid(_argRouteRvmReadOnly_15_io_read_data_valid),
		.io_read_data_task_bits(_argRouteRvmReadOnly_15_io_read_data_bits)
	);
	RVtoAXIBridge_6 argRouteRvm_0(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_0_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_0_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_0_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_0_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_0_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_0_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_0_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_0_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_0_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_0_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_0_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_0_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_0_ar_ready),
		.axi_ar_valid(axi_full_argRoute_0_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_0_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_0_r_ready),
		.axi_r_valid(axi_full_argRoute_0_r_valid),
		.axi_r_bits_data(axi_full_argRoute_0_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_0_aw_ready),
		.axi_aw_valid(axi_full_argRoute_0_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_0_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_0_w_ready),
		.axi_w_valid(axi_full_argRoute_0_w_valid),
		.axi_w_bits_data(axi_full_argRoute_0_w_bits_data),
		.axi_b_valid(axi_full_argRoute_0_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_1(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_1_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_1_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_1_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_1_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_1_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_1_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_1_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_1_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_1_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_1_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_1_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_1_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_1_ar_ready),
		.axi_ar_valid(axi_full_argRoute_1_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_1_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_1_r_ready),
		.axi_r_valid(axi_full_argRoute_1_r_valid),
		.axi_r_bits_data(axi_full_argRoute_1_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_1_aw_ready),
		.axi_aw_valid(axi_full_argRoute_1_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_1_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_1_w_ready),
		.axi_w_valid(axi_full_argRoute_1_w_valid),
		.axi_w_bits_data(axi_full_argRoute_1_w_bits_data),
		.axi_b_valid(axi_full_argRoute_1_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_2(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_2_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_2_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_2_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_2_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_2_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_2_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_2_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_2_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_2_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_2_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_2_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_2_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_2_ar_ready),
		.axi_ar_valid(axi_full_argRoute_2_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_2_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_2_r_ready),
		.axi_r_valid(axi_full_argRoute_2_r_valid),
		.axi_r_bits_data(axi_full_argRoute_2_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_2_aw_ready),
		.axi_aw_valid(axi_full_argRoute_2_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_2_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_2_w_ready),
		.axi_w_valid(axi_full_argRoute_2_w_valid),
		.axi_w_bits_data(axi_full_argRoute_2_w_bits_data),
		.axi_b_valid(axi_full_argRoute_2_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_3(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_3_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_3_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_3_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_3_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_3_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_3_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_3_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_3_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_3_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_3_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_3_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_3_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_3_ar_ready),
		.axi_ar_valid(axi_full_argRoute_3_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_3_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_3_r_ready),
		.axi_r_valid(axi_full_argRoute_3_r_valid),
		.axi_r_bits_data(axi_full_argRoute_3_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_3_aw_ready),
		.axi_aw_valid(axi_full_argRoute_3_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_3_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_3_w_ready),
		.axi_w_valid(axi_full_argRoute_3_w_valid),
		.axi_w_bits_data(axi_full_argRoute_3_w_bits_data),
		.axi_b_valid(axi_full_argRoute_3_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_4(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_4_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_4_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_4_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_4_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_4_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_4_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_4_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_4_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_4_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_4_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_4_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_4_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_4_ar_ready),
		.axi_ar_valid(axi_full_argRoute_4_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_4_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_4_r_ready),
		.axi_r_valid(axi_full_argRoute_4_r_valid),
		.axi_r_bits_data(axi_full_argRoute_4_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_4_aw_ready),
		.axi_aw_valid(axi_full_argRoute_4_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_4_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_4_w_ready),
		.axi_w_valid(axi_full_argRoute_4_w_valid),
		.axi_w_bits_data(axi_full_argRoute_4_w_bits_data),
		.axi_b_valid(axi_full_argRoute_4_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_5(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_5_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_5_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_5_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_5_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_5_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_5_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_5_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_5_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_5_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_5_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_5_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_5_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_5_ar_ready),
		.axi_ar_valid(axi_full_argRoute_5_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_5_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_5_r_ready),
		.axi_r_valid(axi_full_argRoute_5_r_valid),
		.axi_r_bits_data(axi_full_argRoute_5_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_5_aw_ready),
		.axi_aw_valid(axi_full_argRoute_5_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_5_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_5_w_ready),
		.axi_w_valid(axi_full_argRoute_5_w_valid),
		.axi_w_bits_data(axi_full_argRoute_5_w_bits_data),
		.axi_b_valid(axi_full_argRoute_5_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_6(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_6_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_6_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_6_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_6_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_6_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_6_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_6_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_6_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_6_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_6_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_6_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_6_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_6_ar_ready),
		.axi_ar_valid(axi_full_argRoute_6_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_6_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_6_r_ready),
		.axi_r_valid(axi_full_argRoute_6_r_valid),
		.axi_r_bits_data(axi_full_argRoute_6_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_6_aw_ready),
		.axi_aw_valid(axi_full_argRoute_6_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_6_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_6_w_ready),
		.axi_w_valid(axi_full_argRoute_6_w_valid),
		.axi_w_bits_data(axi_full_argRoute_6_w_bits_data),
		.axi_b_valid(axi_full_argRoute_6_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_7(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_7_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_7_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_7_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_7_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_7_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_7_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_7_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_7_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_7_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_7_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_7_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_7_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_7_ar_ready),
		.axi_ar_valid(axi_full_argRoute_7_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_7_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_7_r_ready),
		.axi_r_valid(axi_full_argRoute_7_r_valid),
		.axi_r_bits_data(axi_full_argRoute_7_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_7_aw_ready),
		.axi_aw_valid(axi_full_argRoute_7_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_7_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_7_w_ready),
		.axi_w_valid(axi_full_argRoute_7_w_valid),
		.axi_w_bits_data(axi_full_argRoute_7_w_bits_data),
		.axi_b_valid(axi_full_argRoute_7_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_8(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_8_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_8_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_8_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_8_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_8_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_8_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_8_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_8_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_8_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_8_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_8_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_8_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_8_ar_ready),
		.axi_ar_valid(axi_full_argRoute_8_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_8_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_8_r_ready),
		.axi_r_valid(axi_full_argRoute_8_r_valid),
		.axi_r_bits_data(axi_full_argRoute_8_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_8_aw_ready),
		.axi_aw_valid(axi_full_argRoute_8_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_8_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_8_w_ready),
		.axi_w_valid(axi_full_argRoute_8_w_valid),
		.axi_w_bits_data(axi_full_argRoute_8_w_bits_data),
		.axi_b_valid(axi_full_argRoute_8_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_9(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_9_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_9_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_9_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_9_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_9_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_9_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_9_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_9_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_9_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_9_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_9_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_9_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_9_ar_ready),
		.axi_ar_valid(axi_full_argRoute_9_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_9_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_9_r_ready),
		.axi_r_valid(axi_full_argRoute_9_r_valid),
		.axi_r_bits_data(axi_full_argRoute_9_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_9_aw_ready),
		.axi_aw_valid(axi_full_argRoute_9_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_9_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_9_w_ready),
		.axi_w_valid(axi_full_argRoute_9_w_valid),
		.axi_w_bits_data(axi_full_argRoute_9_w_bits_data),
		.axi_b_valid(axi_full_argRoute_9_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_10(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_10_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_10_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_10_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_10_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_10_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_10_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_10_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_10_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_10_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_10_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_10_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_10_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_10_ar_ready),
		.axi_ar_valid(axi_full_argRoute_10_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_10_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_10_r_ready),
		.axi_r_valid(axi_full_argRoute_10_r_valid),
		.axi_r_bits_data(axi_full_argRoute_10_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_10_aw_ready),
		.axi_aw_valid(axi_full_argRoute_10_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_10_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_10_w_ready),
		.axi_w_valid(axi_full_argRoute_10_w_valid),
		.axi_w_bits_data(axi_full_argRoute_10_w_bits_data),
		.axi_b_valid(axi_full_argRoute_10_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_11(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_11_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_11_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_11_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_11_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_11_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_11_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_11_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_11_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_11_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_11_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_11_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_11_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_11_ar_ready),
		.axi_ar_valid(axi_full_argRoute_11_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_11_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_11_r_ready),
		.axi_r_valid(axi_full_argRoute_11_r_valid),
		.axi_r_bits_data(axi_full_argRoute_11_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_11_aw_ready),
		.axi_aw_valid(axi_full_argRoute_11_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_11_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_11_w_ready),
		.axi_w_valid(axi_full_argRoute_11_w_valid),
		.axi_w_bits_data(axi_full_argRoute_11_w_bits_data),
		.axi_b_valid(axi_full_argRoute_11_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_12(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_12_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_12_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_12_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_12_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_12_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_12_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_12_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_12_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_12_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_12_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_12_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_12_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_12_ar_ready),
		.axi_ar_valid(axi_full_argRoute_12_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_12_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_12_r_ready),
		.axi_r_valid(axi_full_argRoute_12_r_valid),
		.axi_r_bits_data(axi_full_argRoute_12_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_12_aw_ready),
		.axi_aw_valid(axi_full_argRoute_12_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_12_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_12_w_ready),
		.axi_w_valid(axi_full_argRoute_12_w_valid),
		.axi_w_bits_data(axi_full_argRoute_12_w_bits_data),
		.axi_b_valid(axi_full_argRoute_12_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_13(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_13_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_13_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_13_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_13_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_13_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_13_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_13_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_13_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_13_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_13_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_13_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_13_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_13_ar_ready),
		.axi_ar_valid(axi_full_argRoute_13_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_13_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_13_r_ready),
		.axi_r_valid(axi_full_argRoute_13_r_valid),
		.axi_r_bits_data(axi_full_argRoute_13_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_13_aw_ready),
		.axi_aw_valid(axi_full_argRoute_13_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_13_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_13_w_ready),
		.axi_w_valid(axi_full_argRoute_13_w_valid),
		.axi_w_bits_data(axi_full_argRoute_13_w_bits_data),
		.axi_b_valid(axi_full_argRoute_13_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_14(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_14_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_14_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_14_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_14_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_14_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_14_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_14_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_14_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_14_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_14_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_14_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_14_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_14_ar_ready),
		.axi_ar_valid(axi_full_argRoute_14_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_14_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_14_r_ready),
		.axi_r_valid(axi_full_argRoute_14_r_valid),
		.axi_r_bits_data(axi_full_argRoute_14_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_14_aw_ready),
		.axi_aw_valid(axi_full_argRoute_14_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_14_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_14_w_ready),
		.axi_w_valid(axi_full_argRoute_14_w_valid),
		.axi_w_bits_data(axi_full_argRoute_14_w_bits_data),
		.axi_b_valid(axi_full_argRoute_14_b_valid)
	);
	RVtoAXIBridge_6 argRouteRvm_15(
		.clock(clock),
		.reset(reset),
		.io_read_address_ready(_argRouteRvm_15_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_15_io_read_address_valid),
		.io_read_address_bits(_argRouteServers_15_io_read_address_bits),
		.io_read_data_ready(_argRouteServers_15_io_read_data_ready),
		.io_read_data_valid(_argRouteRvm_15_io_read_data_valid),
		.io_read_data_bits(_argRouteRvm_15_io_read_data_bits),
		.io_write_address_ready(_argRouteRvm_15_io_write_address_ready),
		.io_write_address_valid(_argRouteServers_15_io_write_address_valid),
		.io_write_address_bits(_argRouteServers_15_io_write_address_bits),
		.io_write_data_ready(_argRouteRvm_15_io_write_data_ready),
		.io_write_data_valid(_argRouteServers_15_io_write_data_valid),
		.io_write_data_bits(_argRouteServers_15_io_write_data_bits),
		.axi_ar_ready(axi_full_argRoute_15_ar_ready),
		.axi_ar_valid(axi_full_argRoute_15_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_15_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_15_r_ready),
		.axi_r_valid(axi_full_argRoute_15_r_valid),
		.axi_r_bits_data(axi_full_argRoute_15_r_bits_data),
		.axi_aw_ready(axi_full_argRoute_15_aw_ready),
		.axi_aw_valid(axi_full_argRoute_15_aw_valid),
		.axi_aw_bits_addr(axi_full_argRoute_15_aw_bits_addr),
		.axi_w_ready(axi_full_argRoute_15_w_ready),
		.axi_w_valid(axi_full_argRoute_15_w_valid),
		.axi_w_bits_data(axi_full_argRoute_15_w_bits_data),
		.axi_b_valid(axi_full_argRoute_15_b_valid)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_0(
		.io_read_address_ready(_argRouteRvmReadOnly_0_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_0_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_0_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_0_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_0_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_0_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_16_ar_ready),
		.axi_ar_valid(axi_full_argRoute_16_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_16_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_16_r_ready),
		.axi_r_valid(axi_full_argRoute_16_r_valid),
		.axi_r_bits_data(axi_full_argRoute_16_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_1(
		.io_read_address_ready(_argRouteRvmReadOnly_1_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_1_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_1_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_1_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_1_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_1_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_17_ar_ready),
		.axi_ar_valid(axi_full_argRoute_17_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_17_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_17_r_ready),
		.axi_r_valid(axi_full_argRoute_17_r_valid),
		.axi_r_bits_data(axi_full_argRoute_17_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_2(
		.io_read_address_ready(_argRouteRvmReadOnly_2_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_2_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_2_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_2_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_2_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_2_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_18_ar_ready),
		.axi_ar_valid(axi_full_argRoute_18_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_18_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_18_r_ready),
		.axi_r_valid(axi_full_argRoute_18_r_valid),
		.axi_r_bits_data(axi_full_argRoute_18_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_3(
		.io_read_address_ready(_argRouteRvmReadOnly_3_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_3_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_3_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_3_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_3_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_3_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_19_ar_ready),
		.axi_ar_valid(axi_full_argRoute_19_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_19_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_19_r_ready),
		.axi_r_valid(axi_full_argRoute_19_r_valid),
		.axi_r_bits_data(axi_full_argRoute_19_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_4(
		.io_read_address_ready(_argRouteRvmReadOnly_4_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_4_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_4_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_4_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_4_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_4_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_20_ar_ready),
		.axi_ar_valid(axi_full_argRoute_20_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_20_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_20_r_ready),
		.axi_r_valid(axi_full_argRoute_20_r_valid),
		.axi_r_bits_data(axi_full_argRoute_20_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_5(
		.io_read_address_ready(_argRouteRvmReadOnly_5_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_5_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_5_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_5_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_5_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_5_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_21_ar_ready),
		.axi_ar_valid(axi_full_argRoute_21_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_21_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_21_r_ready),
		.axi_r_valid(axi_full_argRoute_21_r_valid),
		.axi_r_bits_data(axi_full_argRoute_21_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_6(
		.io_read_address_ready(_argRouteRvmReadOnly_6_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_6_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_6_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_6_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_6_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_6_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_22_ar_ready),
		.axi_ar_valid(axi_full_argRoute_22_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_22_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_22_r_ready),
		.axi_r_valid(axi_full_argRoute_22_r_valid),
		.axi_r_bits_data(axi_full_argRoute_22_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_7(
		.io_read_address_ready(_argRouteRvmReadOnly_7_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_7_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_7_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_7_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_7_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_7_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_23_ar_ready),
		.axi_ar_valid(axi_full_argRoute_23_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_23_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_23_r_ready),
		.axi_r_valid(axi_full_argRoute_23_r_valid),
		.axi_r_bits_data(axi_full_argRoute_23_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_8(
		.io_read_address_ready(_argRouteRvmReadOnly_8_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_8_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_8_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_8_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_8_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_8_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_24_ar_ready),
		.axi_ar_valid(axi_full_argRoute_24_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_24_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_24_r_ready),
		.axi_r_valid(axi_full_argRoute_24_r_valid),
		.axi_r_bits_data(axi_full_argRoute_24_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_9(
		.io_read_address_ready(_argRouteRvmReadOnly_9_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_9_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_9_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_9_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_9_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_9_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_25_ar_ready),
		.axi_ar_valid(axi_full_argRoute_25_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_25_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_25_r_ready),
		.axi_r_valid(axi_full_argRoute_25_r_valid),
		.axi_r_bits_data(axi_full_argRoute_25_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_10(
		.io_read_address_ready(_argRouteRvmReadOnly_10_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_10_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_10_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_10_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_10_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_10_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_26_ar_ready),
		.axi_ar_valid(axi_full_argRoute_26_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_26_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_26_r_ready),
		.axi_r_valid(axi_full_argRoute_26_r_valid),
		.axi_r_bits_data(axi_full_argRoute_26_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_11(
		.io_read_address_ready(_argRouteRvmReadOnly_11_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_11_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_11_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_11_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_11_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_11_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_27_ar_ready),
		.axi_ar_valid(axi_full_argRoute_27_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_27_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_27_r_ready),
		.axi_r_valid(axi_full_argRoute_27_r_valid),
		.axi_r_bits_data(axi_full_argRoute_27_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_12(
		.io_read_address_ready(_argRouteRvmReadOnly_12_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_12_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_12_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_12_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_12_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_12_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_28_ar_ready),
		.axi_ar_valid(axi_full_argRoute_28_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_28_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_28_r_ready),
		.axi_r_valid(axi_full_argRoute_28_r_valid),
		.axi_r_bits_data(axi_full_argRoute_28_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_13(
		.io_read_address_ready(_argRouteRvmReadOnly_13_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_13_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_13_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_13_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_13_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_13_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_29_ar_ready),
		.axi_ar_valid(axi_full_argRoute_29_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_29_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_29_r_ready),
		.axi_r_valid(axi_full_argRoute_29_r_valid),
		.axi_r_bits_data(axi_full_argRoute_29_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_14(
		.io_read_address_ready(_argRouteRvmReadOnly_14_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_14_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_14_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_14_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_14_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_14_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_30_ar_ready),
		.axi_ar_valid(axi_full_argRoute_30_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_30_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_30_r_ready),
		.axi_r_valid(axi_full_argRoute_30_r_valid),
		.axi_r_bits_data(axi_full_argRoute_30_r_bits_data)
	);
	RVtoAXIBridge_22 argRouteRvmReadOnly_15(
		.io_read_address_ready(_argRouteRvmReadOnly_15_io_read_address_ready),
		.io_read_address_valid(_argRouteServers_15_io_read_address_task_valid),
		.io_read_address_bits(_argRouteServers_15_io_read_address_task_bits),
		.io_read_data_ready(_argRouteServers_15_io_read_data_task_ready),
		.io_read_data_valid(_argRouteRvmReadOnly_15_io_read_data_valid),
		.io_read_data_bits(_argRouteRvmReadOnly_15_io_read_data_bits),
		.axi_ar_ready(axi_full_argRoute_31_ar_ready),
		.axi_ar_valid(axi_full_argRoute_31_ar_valid),
		.axi_ar_bits_addr(axi_full_argRoute_31_ar_bits_addr),
		.axi_r_ready(axi_full_argRoute_31_r_ready),
		.axi_r_valid(axi_full_argRoute_31_r_valid),
		.axi_r_bits_data(axi_full_argRoute_31_r_bits_data)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_0(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_0_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_0_TVALID),
		.io_dataIn_TDATA(io_export_argIn_0_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_0_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_0_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_0_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_1(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_1_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_1_TVALID),
		.io_dataIn_TDATA(io_export_argIn_1_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_1_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_1_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_1_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_2(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_2_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_2_TVALID),
		.io_dataIn_TDATA(io_export_argIn_2_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_2_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_2_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_2_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_3(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_3_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_3_TVALID),
		.io_dataIn_TDATA(io_export_argIn_3_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_3_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_3_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_3_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_4(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_4_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_4_TVALID),
		.io_dataIn_TDATA(io_export_argIn_4_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_4_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_4_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_4_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_5(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_5_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_5_TVALID),
		.io_dataIn_TDATA(io_export_argIn_5_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_5_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_5_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_5_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_6(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_6_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_6_TVALID),
		.io_dataIn_TDATA(io_export_argIn_6_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_6_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_6_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_6_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_7(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_7_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_7_TVALID),
		.io_dataIn_TDATA(io_export_argIn_7_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_7_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_7_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_7_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_8(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_8_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_8_TVALID),
		.io_dataIn_TDATA(io_export_argIn_8_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_8_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_8_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_8_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_9(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_9_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_9_TVALID),
		.io_dataIn_TDATA(io_export_argIn_9_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_9_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_9_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_9_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_10(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_10_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_10_TVALID),
		.io_dataIn_TDATA(io_export_argIn_10_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_10_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_10_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_10_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_11(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_11_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_11_TVALID),
		.io_dataIn_TDATA(io_export_argIn_11_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_11_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_11_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_11_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_12(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_12_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_12_TVALID),
		.io_dataIn_TDATA(io_export_argIn_12_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_12_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_12_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_12_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_13(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_13_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_13_TVALID),
		.io_dataIn_TDATA(io_export_argIn_13_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_13_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_13_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_13_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_14(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_14_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_14_TVALID),
		.io_dataIn_TDATA(io_export_argIn_14_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_14_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_14_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_14_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_15(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_15_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_15_TVALID),
		.io_dataIn_TDATA(io_export_argIn_15_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_15_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_15_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_15_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_16(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_16_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_16_TVALID),
		.io_dataIn_TDATA(io_export_argIn_16_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_16_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_16_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_16_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_17(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_17_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_17_TVALID),
		.io_dataIn_TDATA(io_export_argIn_17_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_17_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_17_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_17_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_18(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_18_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_18_TVALID),
		.io_dataIn_TDATA(io_export_argIn_18_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_18_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_18_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_18_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_19(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_19_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_19_TVALID),
		.io_dataIn_TDATA(io_export_argIn_19_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_19_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_19_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_19_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_20(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_20_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_20_TVALID),
		.io_dataIn_TDATA(io_export_argIn_20_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_20_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_20_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_20_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_21(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_21_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_21_TVALID),
		.io_dataIn_TDATA(io_export_argIn_21_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_21_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_21_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_21_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_22(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_22_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_22_TVALID),
		.io_dataIn_TDATA(io_export_argIn_22_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_22_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_22_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_22_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_23(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_23_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_23_TVALID),
		.io_dataIn_TDATA(io_export_argIn_23_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_23_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_23_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_23_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_24(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_24_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_24_TVALID),
		.io_dataIn_TDATA(io_export_argIn_24_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_24_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_24_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_24_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_25(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_25_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_25_TVALID),
		.io_dataIn_TDATA(io_export_argIn_25_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_25_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_25_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_25_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_26(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_26_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_26_TVALID),
		.io_dataIn_TDATA(io_export_argIn_26_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_26_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_26_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_26_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_27(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_27_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_27_TVALID),
		.io_dataIn_TDATA(io_export_argIn_27_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_27_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_27_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_27_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_28(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_28_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_28_TVALID),
		.io_dataIn_TDATA(io_export_argIn_28_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_28_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_28_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_28_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_29(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_29_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_29_TVALID),
		.io_dataIn_TDATA(io_export_argIn_29_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_29_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_29_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_29_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_30(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_30_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_30_TVALID),
		.io_dataIn_TDATA(io_export_argIn_30_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_30_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_30_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_30_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_31(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_31_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_31_TVALID),
		.io_dataIn_TDATA(io_export_argIn_31_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_31_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_31_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_31_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_32(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_32_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_32_TVALID),
		.io_dataIn_TDATA(io_export_argIn_32_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_32_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_32_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_32_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_33(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_33_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_33_TVALID),
		.io_dataIn_TDATA(io_export_argIn_33_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_33_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_33_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_33_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_34(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_34_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_34_TVALID),
		.io_dataIn_TDATA(io_export_argIn_34_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_34_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_34_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_34_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_35(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_35_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_35_TVALID),
		.io_dataIn_TDATA(io_export_argIn_35_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_35_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_35_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_35_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_36(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_36_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_36_TVALID),
		.io_dataIn_TDATA(io_export_argIn_36_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_36_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_36_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_36_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_37(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_37_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_37_TVALID),
		.io_dataIn_TDATA(io_export_argIn_37_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_37_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_37_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_37_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_38(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_38_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_38_TVALID),
		.io_dataIn_TDATA(io_export_argIn_38_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_38_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_38_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_38_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_39(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_39_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_39_TVALID),
		.io_dataIn_TDATA(io_export_argIn_39_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_39_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_39_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_39_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_40(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_40_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_40_TVALID),
		.io_dataIn_TDATA(io_export_argIn_40_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_40_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_40_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_40_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_41(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_41_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_41_TVALID),
		.io_dataIn_TDATA(io_export_argIn_41_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_41_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_41_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_41_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_42(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_42_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_42_TVALID),
		.io_dataIn_TDATA(io_export_argIn_42_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_42_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_42_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_42_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_43(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_43_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_43_TVALID),
		.io_dataIn_TDATA(io_export_argIn_43_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_43_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_43_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_43_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_44(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_44_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_44_TVALID),
		.io_dataIn_TDATA(io_export_argIn_44_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_44_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_44_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_44_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_45(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_45_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_45_TVALID),
		.io_dataIn_TDATA(io_export_argIn_45_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_45_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_45_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_45_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_46(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_46_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_46_TVALID),
		.io_dataIn_TDATA(io_export_argIn_46_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_46_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_46_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_46_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_47(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_47_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_47_TVALID),
		.io_dataIn_TDATA(io_export_argIn_47_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_47_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_47_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_47_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_48(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_48_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_48_TVALID),
		.io_dataIn_TDATA(io_export_argIn_48_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_48_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_48_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_48_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_49(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_49_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_49_TVALID),
		.io_dataIn_TDATA(io_export_argIn_49_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_49_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_49_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_49_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_50(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_50_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_50_TVALID),
		.io_dataIn_TDATA(io_export_argIn_50_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_50_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_50_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_50_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_51(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_51_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_51_TVALID),
		.io_dataIn_TDATA(io_export_argIn_51_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_51_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_51_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_51_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_52(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_52_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_52_TVALID),
		.io_dataIn_TDATA(io_export_argIn_52_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_52_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_52_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_52_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_53(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_53_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_53_TVALID),
		.io_dataIn_TDATA(io_export_argIn_53_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_53_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_53_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_53_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_54(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_54_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_54_TVALID),
		.io_dataIn_TDATA(io_export_argIn_54_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_54_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_54_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_54_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_55(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_55_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_55_TVALID),
		.io_dataIn_TDATA(io_export_argIn_55_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_55_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_55_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_55_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_56(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_56_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_56_TVALID),
		.io_dataIn_TDATA(io_export_argIn_56_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_56_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_56_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_56_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_57(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_57_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_57_TVALID),
		.io_dataIn_TDATA(io_export_argIn_57_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_57_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_57_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_57_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_58(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_58_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_58_TVALID),
		.io_dataIn_TDATA(io_export_argIn_58_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_58_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_58_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_58_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_59(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_59_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_59_TVALID),
		.io_dataIn_TDATA(io_export_argIn_59_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_59_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_59_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_59_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_60(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_60_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_60_TVALID),
		.io_dataIn_TDATA(io_export_argIn_60_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_60_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_60_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_60_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_61(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_61_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_61_TVALID),
		.io_dataIn_TDATA(io_export_argIn_61_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_61_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_61_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_61_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_62(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_62_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_62_TVALID),
		.io_dataIn_TDATA(io_export_argIn_62_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_62_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_62_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_62_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_63(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_63_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_63_TVALID),
		.io_dataIn_TDATA(io_export_argIn_63_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_63_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_63_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_63_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_64(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_64_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_64_TVALID),
		.io_dataIn_TDATA(io_export_argIn_64_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_64_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_64_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_64_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_65(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_65_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_65_TVALID),
		.io_dataIn_TDATA(io_export_argIn_65_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_65_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_65_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_65_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_66(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_66_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_66_TVALID),
		.io_dataIn_TDATA(io_export_argIn_66_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_66_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_66_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_66_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_67(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_67_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_67_TVALID),
		.io_dataIn_TDATA(io_export_argIn_67_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_67_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_67_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_67_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_68(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_68_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_68_TVALID),
		.io_dataIn_TDATA(io_export_argIn_68_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_68_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_68_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_68_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_69(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_69_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_69_TVALID),
		.io_dataIn_TDATA(io_export_argIn_69_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_69_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_69_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_69_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_70(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_70_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_70_TVALID),
		.io_dataIn_TDATA(io_export_argIn_70_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_70_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_70_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_70_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_71(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_71_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_71_TVALID),
		.io_dataIn_TDATA(io_export_argIn_71_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_71_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_71_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_71_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_72(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_72_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_72_TVALID),
		.io_dataIn_TDATA(io_export_argIn_72_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_72_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_72_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_72_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_73(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_73_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_73_TVALID),
		.io_dataIn_TDATA(io_export_argIn_73_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_73_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_73_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_73_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_74(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_74_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_74_TVALID),
		.io_dataIn_TDATA(io_export_argIn_74_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_74_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_74_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_74_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_75(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_75_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_75_TVALID),
		.io_dataIn_TDATA(io_export_argIn_75_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_75_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_75_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_75_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_76(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_76_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_76_TVALID),
		.io_dataIn_TDATA(io_export_argIn_76_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_76_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_76_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_76_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_77(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_77_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_77_TVALID),
		.io_dataIn_TDATA(io_export_argIn_77_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_77_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_77_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_77_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_78(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_78_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_78_TVALID),
		.io_dataIn_TDATA(io_export_argIn_78_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_78_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_78_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_78_io_dataOut_TDATA)
	);
	AxisDataWidthConverter_208 axis_stream_converters_in_79(
		.clock(clock),
		.reset(reset),
		.io_dataIn_TREADY(_axis_stream_converters_in_79_io_dataIn_TREADY),
		.io_dataIn_TVALID(io_export_argIn_79_TVALID),
		.io_dataIn_TDATA(io_export_argIn_79_TDATA),
		.io_dataOut_TREADY(_argSide_io_connPE_79_ready),
		.io_dataOut_TVALID(_axis_stream_converters_in_79_io_dataOut_TVALID),
		.io_dataOut_TDATA(_axis_stream_converters_in_79_io_dataOut_TDATA)
	);
	Counter64 argInCounter(
		.clock(clock),
		.reset(reset),
		.io_signals_0(io_export_argIn_0_TVALID & _axis_stream_converters_in_0_io_dataIn_TREADY),
		.io_signals_1(io_export_argIn_1_TVALID & _axis_stream_converters_in_1_io_dataIn_TREADY),
		.io_signals_2(io_export_argIn_2_TVALID & _axis_stream_converters_in_2_io_dataIn_TREADY),
		.io_signals_3(io_export_argIn_3_TVALID & _axis_stream_converters_in_3_io_dataIn_TREADY),
		.io_signals_4(io_export_argIn_4_TVALID & _axis_stream_converters_in_4_io_dataIn_TREADY),
		.io_signals_5(io_export_argIn_5_TVALID & _axis_stream_converters_in_5_io_dataIn_TREADY),
		.io_signals_6(io_export_argIn_6_TVALID & _axis_stream_converters_in_6_io_dataIn_TREADY),
		.io_signals_7(io_export_argIn_7_TVALID & _axis_stream_converters_in_7_io_dataIn_TREADY),
		.io_signals_8(io_export_argIn_8_TVALID & _axis_stream_converters_in_8_io_dataIn_TREADY),
		.io_signals_9(io_export_argIn_9_TVALID & _axis_stream_converters_in_9_io_dataIn_TREADY),
		.io_signals_10(io_export_argIn_10_TVALID & _axis_stream_converters_in_10_io_dataIn_TREADY),
		.io_signals_11(io_export_argIn_11_TVALID & _axis_stream_converters_in_11_io_dataIn_TREADY),
		.io_signals_12(io_export_argIn_12_TVALID & _axis_stream_converters_in_12_io_dataIn_TREADY),
		.io_signals_13(io_export_argIn_13_TVALID & _axis_stream_converters_in_13_io_dataIn_TREADY),
		.io_signals_14(io_export_argIn_14_TVALID & _axis_stream_converters_in_14_io_dataIn_TREADY),
		.io_signals_15(io_export_argIn_15_TVALID & _axis_stream_converters_in_15_io_dataIn_TREADY),
		.io_signals_16(io_export_argIn_16_TVALID & _axis_stream_converters_in_16_io_dataIn_TREADY),
		.io_signals_17(io_export_argIn_17_TVALID & _axis_stream_converters_in_17_io_dataIn_TREADY),
		.io_signals_18(io_export_argIn_18_TVALID & _axis_stream_converters_in_18_io_dataIn_TREADY),
		.io_signals_19(io_export_argIn_19_TVALID & _axis_stream_converters_in_19_io_dataIn_TREADY),
		.io_signals_20(io_export_argIn_20_TVALID & _axis_stream_converters_in_20_io_dataIn_TREADY),
		.io_signals_21(io_export_argIn_21_TVALID & _axis_stream_converters_in_21_io_dataIn_TREADY),
		.io_signals_22(io_export_argIn_22_TVALID & _axis_stream_converters_in_22_io_dataIn_TREADY),
		.io_signals_23(io_export_argIn_23_TVALID & _axis_stream_converters_in_23_io_dataIn_TREADY),
		.io_signals_24(io_export_argIn_24_TVALID & _axis_stream_converters_in_24_io_dataIn_TREADY),
		.io_signals_25(io_export_argIn_25_TVALID & _axis_stream_converters_in_25_io_dataIn_TREADY),
		.io_signals_26(io_export_argIn_26_TVALID & _axis_stream_converters_in_26_io_dataIn_TREADY),
		.io_signals_27(io_export_argIn_27_TVALID & _axis_stream_converters_in_27_io_dataIn_TREADY),
		.io_signals_28(io_export_argIn_28_TVALID & _axis_stream_converters_in_28_io_dataIn_TREADY),
		.io_signals_29(io_export_argIn_29_TVALID & _axis_stream_converters_in_29_io_dataIn_TREADY),
		.io_signals_30(io_export_argIn_30_TVALID & _axis_stream_converters_in_30_io_dataIn_TREADY),
		.io_signals_31(io_export_argIn_31_TVALID & _axis_stream_converters_in_31_io_dataIn_TREADY),
		.io_signals_32(io_export_argIn_32_TVALID & _axis_stream_converters_in_32_io_dataIn_TREADY),
		.io_signals_33(io_export_argIn_33_TVALID & _axis_stream_converters_in_33_io_dataIn_TREADY),
		.io_signals_34(io_export_argIn_34_TVALID & _axis_stream_converters_in_34_io_dataIn_TREADY),
		.io_signals_35(io_export_argIn_35_TVALID & _axis_stream_converters_in_35_io_dataIn_TREADY),
		.io_signals_36(io_export_argIn_36_TVALID & _axis_stream_converters_in_36_io_dataIn_TREADY),
		.io_signals_37(io_export_argIn_37_TVALID & _axis_stream_converters_in_37_io_dataIn_TREADY),
		.io_signals_38(io_export_argIn_38_TVALID & _axis_stream_converters_in_38_io_dataIn_TREADY),
		.io_signals_39(io_export_argIn_39_TVALID & _axis_stream_converters_in_39_io_dataIn_TREADY),
		.io_signals_40(io_export_argIn_40_TVALID & _axis_stream_converters_in_40_io_dataIn_TREADY),
		.io_signals_41(io_export_argIn_41_TVALID & _axis_stream_converters_in_41_io_dataIn_TREADY),
		.io_signals_42(io_export_argIn_42_TVALID & _axis_stream_converters_in_42_io_dataIn_TREADY),
		.io_signals_43(io_export_argIn_43_TVALID & _axis_stream_converters_in_43_io_dataIn_TREADY),
		.io_signals_44(io_export_argIn_44_TVALID & _axis_stream_converters_in_44_io_dataIn_TREADY),
		.io_signals_45(io_export_argIn_45_TVALID & _axis_stream_converters_in_45_io_dataIn_TREADY),
		.io_signals_46(io_export_argIn_46_TVALID & _axis_stream_converters_in_46_io_dataIn_TREADY),
		.io_signals_47(io_export_argIn_47_TVALID & _axis_stream_converters_in_47_io_dataIn_TREADY),
		.io_signals_48(io_export_argIn_48_TVALID & _axis_stream_converters_in_48_io_dataIn_TREADY),
		.io_signals_49(io_export_argIn_49_TVALID & _axis_stream_converters_in_49_io_dataIn_TREADY),
		.io_signals_50(io_export_argIn_50_TVALID & _axis_stream_converters_in_50_io_dataIn_TREADY),
		.io_signals_51(io_export_argIn_51_TVALID & _axis_stream_converters_in_51_io_dataIn_TREADY),
		.io_signals_52(io_export_argIn_52_TVALID & _axis_stream_converters_in_52_io_dataIn_TREADY),
		.io_signals_53(io_export_argIn_53_TVALID & _axis_stream_converters_in_53_io_dataIn_TREADY),
		.io_signals_54(io_export_argIn_54_TVALID & _axis_stream_converters_in_54_io_dataIn_TREADY),
		.io_signals_55(io_export_argIn_55_TVALID & _axis_stream_converters_in_55_io_dataIn_TREADY),
		.io_signals_56(io_export_argIn_56_TVALID & _axis_stream_converters_in_56_io_dataIn_TREADY),
		.io_signals_57(io_export_argIn_57_TVALID & _axis_stream_converters_in_57_io_dataIn_TREADY),
		.io_signals_58(io_export_argIn_58_TVALID & _axis_stream_converters_in_58_io_dataIn_TREADY),
		.io_signals_59(io_export_argIn_59_TVALID & _axis_stream_converters_in_59_io_dataIn_TREADY),
		.io_signals_60(io_export_argIn_60_TVALID & _axis_stream_converters_in_60_io_dataIn_TREADY),
		.io_signals_61(io_export_argIn_61_TVALID & _axis_stream_converters_in_61_io_dataIn_TREADY),
		.io_signals_62(io_export_argIn_62_TVALID & _axis_stream_converters_in_62_io_dataIn_TREADY),
		.io_signals_63(io_export_argIn_63_TVALID & _axis_stream_converters_in_63_io_dataIn_TREADY),
		.io_signals_64(io_export_argIn_64_TVALID & _axis_stream_converters_in_64_io_dataIn_TREADY),
		.io_signals_65(io_export_argIn_65_TVALID & _axis_stream_converters_in_65_io_dataIn_TREADY),
		.io_signals_66(io_export_argIn_66_TVALID & _axis_stream_converters_in_66_io_dataIn_TREADY),
		.io_signals_67(io_export_argIn_67_TVALID & _axis_stream_converters_in_67_io_dataIn_TREADY),
		.io_signals_68(io_export_argIn_68_TVALID & _axis_stream_converters_in_68_io_dataIn_TREADY),
		.io_signals_69(io_export_argIn_69_TVALID & _axis_stream_converters_in_69_io_dataIn_TREADY),
		.io_signals_70(io_export_argIn_70_TVALID & _axis_stream_converters_in_70_io_dataIn_TREADY),
		.io_signals_71(io_export_argIn_71_TVALID & _axis_stream_converters_in_71_io_dataIn_TREADY),
		.io_signals_72(io_export_argIn_72_TVALID & _axis_stream_converters_in_72_io_dataIn_TREADY),
		.io_signals_73(io_export_argIn_73_TVALID & _axis_stream_converters_in_73_io_dataIn_TREADY),
		.io_signals_74(io_export_argIn_74_TVALID & _axis_stream_converters_in_74_io_dataIn_TREADY),
		.io_signals_75(io_export_argIn_75_TVALID & _axis_stream_converters_in_75_io_dataIn_TREADY),
		.io_signals_76(io_export_argIn_76_TVALID & _axis_stream_converters_in_76_io_dataIn_TREADY),
		.io_signals_77(io_export_argIn_77_TVALID & _axis_stream_converters_in_77_io_dataIn_TREADY),
		.io_signals_78(io_export_argIn_78_TVALID & _axis_stream_converters_in_78_io_dataIn_TREADY),
		.io_signals_79(io_export_argIn_79_TVALID & _axis_stream_converters_in_79_io_dataIn_TREADY),
		.io_counter()
	);
	assign io_export_argIn_0_TREADY = _axis_stream_converters_in_0_io_dataIn_TREADY;
	assign io_export_argIn_1_TREADY = _axis_stream_converters_in_1_io_dataIn_TREADY;
	assign io_export_argIn_2_TREADY = _axis_stream_converters_in_2_io_dataIn_TREADY;
	assign io_export_argIn_3_TREADY = _axis_stream_converters_in_3_io_dataIn_TREADY;
	assign io_export_argIn_4_TREADY = _axis_stream_converters_in_4_io_dataIn_TREADY;
	assign io_export_argIn_5_TREADY = _axis_stream_converters_in_5_io_dataIn_TREADY;
	assign io_export_argIn_6_TREADY = _axis_stream_converters_in_6_io_dataIn_TREADY;
	assign io_export_argIn_7_TREADY = _axis_stream_converters_in_7_io_dataIn_TREADY;
	assign io_export_argIn_8_TREADY = _axis_stream_converters_in_8_io_dataIn_TREADY;
	assign io_export_argIn_9_TREADY = _axis_stream_converters_in_9_io_dataIn_TREADY;
	assign io_export_argIn_10_TREADY = _axis_stream_converters_in_10_io_dataIn_TREADY;
	assign io_export_argIn_11_TREADY = _axis_stream_converters_in_11_io_dataIn_TREADY;
	assign io_export_argIn_12_TREADY = _axis_stream_converters_in_12_io_dataIn_TREADY;
	assign io_export_argIn_13_TREADY = _axis_stream_converters_in_13_io_dataIn_TREADY;
	assign io_export_argIn_14_TREADY = _axis_stream_converters_in_14_io_dataIn_TREADY;
	assign io_export_argIn_15_TREADY = _axis_stream_converters_in_15_io_dataIn_TREADY;
	assign io_export_argIn_16_TREADY = _axis_stream_converters_in_16_io_dataIn_TREADY;
	assign io_export_argIn_17_TREADY = _axis_stream_converters_in_17_io_dataIn_TREADY;
	assign io_export_argIn_18_TREADY = _axis_stream_converters_in_18_io_dataIn_TREADY;
	assign io_export_argIn_19_TREADY = _axis_stream_converters_in_19_io_dataIn_TREADY;
	assign io_export_argIn_20_TREADY = _axis_stream_converters_in_20_io_dataIn_TREADY;
	assign io_export_argIn_21_TREADY = _axis_stream_converters_in_21_io_dataIn_TREADY;
	assign io_export_argIn_22_TREADY = _axis_stream_converters_in_22_io_dataIn_TREADY;
	assign io_export_argIn_23_TREADY = _axis_stream_converters_in_23_io_dataIn_TREADY;
	assign io_export_argIn_24_TREADY = _axis_stream_converters_in_24_io_dataIn_TREADY;
	assign io_export_argIn_25_TREADY = _axis_stream_converters_in_25_io_dataIn_TREADY;
	assign io_export_argIn_26_TREADY = _axis_stream_converters_in_26_io_dataIn_TREADY;
	assign io_export_argIn_27_TREADY = _axis_stream_converters_in_27_io_dataIn_TREADY;
	assign io_export_argIn_28_TREADY = _axis_stream_converters_in_28_io_dataIn_TREADY;
	assign io_export_argIn_29_TREADY = _axis_stream_converters_in_29_io_dataIn_TREADY;
	assign io_export_argIn_30_TREADY = _axis_stream_converters_in_30_io_dataIn_TREADY;
	assign io_export_argIn_31_TREADY = _axis_stream_converters_in_31_io_dataIn_TREADY;
	assign io_export_argIn_32_TREADY = _axis_stream_converters_in_32_io_dataIn_TREADY;
	assign io_export_argIn_33_TREADY = _axis_stream_converters_in_33_io_dataIn_TREADY;
	assign io_export_argIn_34_TREADY = _axis_stream_converters_in_34_io_dataIn_TREADY;
	assign io_export_argIn_35_TREADY = _axis_stream_converters_in_35_io_dataIn_TREADY;
	assign io_export_argIn_36_TREADY = _axis_stream_converters_in_36_io_dataIn_TREADY;
	assign io_export_argIn_37_TREADY = _axis_stream_converters_in_37_io_dataIn_TREADY;
	assign io_export_argIn_38_TREADY = _axis_stream_converters_in_38_io_dataIn_TREADY;
	assign io_export_argIn_39_TREADY = _axis_stream_converters_in_39_io_dataIn_TREADY;
	assign io_export_argIn_40_TREADY = _axis_stream_converters_in_40_io_dataIn_TREADY;
	assign io_export_argIn_41_TREADY = _axis_stream_converters_in_41_io_dataIn_TREADY;
	assign io_export_argIn_42_TREADY = _axis_stream_converters_in_42_io_dataIn_TREADY;
	assign io_export_argIn_43_TREADY = _axis_stream_converters_in_43_io_dataIn_TREADY;
	assign io_export_argIn_44_TREADY = _axis_stream_converters_in_44_io_dataIn_TREADY;
	assign io_export_argIn_45_TREADY = _axis_stream_converters_in_45_io_dataIn_TREADY;
	assign io_export_argIn_46_TREADY = _axis_stream_converters_in_46_io_dataIn_TREADY;
	assign io_export_argIn_47_TREADY = _axis_stream_converters_in_47_io_dataIn_TREADY;
	assign io_export_argIn_48_TREADY = _axis_stream_converters_in_48_io_dataIn_TREADY;
	assign io_export_argIn_49_TREADY = _axis_stream_converters_in_49_io_dataIn_TREADY;
	assign io_export_argIn_50_TREADY = _axis_stream_converters_in_50_io_dataIn_TREADY;
	assign io_export_argIn_51_TREADY = _axis_stream_converters_in_51_io_dataIn_TREADY;
	assign io_export_argIn_52_TREADY = _axis_stream_converters_in_52_io_dataIn_TREADY;
	assign io_export_argIn_53_TREADY = _axis_stream_converters_in_53_io_dataIn_TREADY;
	assign io_export_argIn_54_TREADY = _axis_stream_converters_in_54_io_dataIn_TREADY;
	assign io_export_argIn_55_TREADY = _axis_stream_converters_in_55_io_dataIn_TREADY;
	assign io_export_argIn_56_TREADY = _axis_stream_converters_in_56_io_dataIn_TREADY;
	assign io_export_argIn_57_TREADY = _axis_stream_converters_in_57_io_dataIn_TREADY;
	assign io_export_argIn_58_TREADY = _axis_stream_converters_in_58_io_dataIn_TREADY;
	assign io_export_argIn_59_TREADY = _axis_stream_converters_in_59_io_dataIn_TREADY;
	assign io_export_argIn_60_TREADY = _axis_stream_converters_in_60_io_dataIn_TREADY;
	assign io_export_argIn_61_TREADY = _axis_stream_converters_in_61_io_dataIn_TREADY;
	assign io_export_argIn_62_TREADY = _axis_stream_converters_in_62_io_dataIn_TREADY;
	assign io_export_argIn_63_TREADY = _axis_stream_converters_in_63_io_dataIn_TREADY;
	assign io_export_argIn_64_TREADY = _axis_stream_converters_in_64_io_dataIn_TREADY;
	assign io_export_argIn_65_TREADY = _axis_stream_converters_in_65_io_dataIn_TREADY;
	assign io_export_argIn_66_TREADY = _axis_stream_converters_in_66_io_dataIn_TREADY;
	assign io_export_argIn_67_TREADY = _axis_stream_converters_in_67_io_dataIn_TREADY;
	assign io_export_argIn_68_TREADY = _axis_stream_converters_in_68_io_dataIn_TREADY;
	assign io_export_argIn_69_TREADY = _axis_stream_converters_in_69_io_dataIn_TREADY;
	assign io_export_argIn_70_TREADY = _axis_stream_converters_in_70_io_dataIn_TREADY;
	assign io_export_argIn_71_TREADY = _axis_stream_converters_in_71_io_dataIn_TREADY;
	assign io_export_argIn_72_TREADY = _axis_stream_converters_in_72_io_dataIn_TREADY;
	assign io_export_argIn_73_TREADY = _axis_stream_converters_in_73_io_dataIn_TREADY;
	assign io_export_argIn_74_TREADY = _axis_stream_converters_in_74_io_dataIn_TREADY;
	assign io_export_argIn_75_TREADY = _axis_stream_converters_in_75_io_dataIn_TREADY;
	assign io_export_argIn_76_TREADY = _axis_stream_converters_in_76_io_dataIn_TREADY;
	assign io_export_argIn_77_TREADY = _axis_stream_converters_in_77_io_dataIn_TREADY;
	assign io_export_argIn_78_TREADY = _axis_stream_converters_in_78_io_dataIn_TREADY;
	assign io_export_argIn_79_TREADY = _axis_stream_converters_in_79_io_dataIn_TREADY;
endmodule
module quickSort (
	clock,
	reset,
	s_axil_mgmt_hardcilk_ARREADY,
	s_axil_mgmt_hardcilk_ARVALID,
	s_axil_mgmt_hardcilk_ARADDR,
	s_axil_mgmt_hardcilk_ARPROT,
	s_axil_mgmt_hardcilk_RREADY,
	s_axil_mgmt_hardcilk_RVALID,
	s_axil_mgmt_hardcilk_RDATA,
	s_axil_mgmt_hardcilk_RRESP,
	s_axil_mgmt_hardcilk_AWREADY,
	s_axil_mgmt_hardcilk_AWVALID,
	s_axil_mgmt_hardcilk_AWADDR,
	s_axil_mgmt_hardcilk_AWPROT,
	s_axil_mgmt_hardcilk_WREADY,
	s_axil_mgmt_hardcilk_WVALID,
	s_axil_mgmt_hardcilk_WDATA,
	s_axil_mgmt_hardcilk_WSTRB,
	s_axil_mgmt_hardcilk_BREADY,
	s_axil_mgmt_hardcilk_BVALID,
	s_axil_mgmt_hardcilk_BRESP,
	qsort_0_m_axi_gmem_ARREADY,
	qsort_0_m_axi_gmem_ARVALID,
	qsort_0_m_axi_gmem_ARID,
	qsort_0_m_axi_gmem_ARADDR,
	qsort_0_m_axi_gmem_ARLEN,
	qsort_0_m_axi_gmem_ARSIZE,
	qsort_0_m_axi_gmem_ARBURST,
	qsort_0_m_axi_gmem_ARLOCK,
	qsort_0_m_axi_gmem_ARCACHE,
	qsort_0_m_axi_gmem_ARPROT,
	qsort_0_m_axi_gmem_ARQOS,
	qsort_0_m_axi_gmem_ARREGION,
	qsort_0_m_axi_gmem_ARUSER,
	qsort_0_m_axi_gmem_RREADY,
	qsort_0_m_axi_gmem_RVALID,
	qsort_0_m_axi_gmem_RID,
	qsort_0_m_axi_gmem_RDATA,
	qsort_0_m_axi_gmem_RRESP,
	qsort_0_m_axi_gmem_RLAST,
	qsort_0_m_axi_gmem_RUSER,
	qsort_0_m_axi_gmem_AWREADY,
	qsort_0_m_axi_gmem_AWVALID,
	qsort_0_m_axi_gmem_AWID,
	qsort_0_m_axi_gmem_AWADDR,
	qsort_0_m_axi_gmem_AWLEN,
	qsort_0_m_axi_gmem_AWSIZE,
	qsort_0_m_axi_gmem_AWBURST,
	qsort_0_m_axi_gmem_AWLOCK,
	qsort_0_m_axi_gmem_AWCACHE,
	qsort_0_m_axi_gmem_AWPROT,
	qsort_0_m_axi_gmem_AWQOS,
	qsort_0_m_axi_gmem_AWREGION,
	qsort_0_m_axi_gmem_AWUSER,
	qsort_0_m_axi_gmem_WREADY,
	qsort_0_m_axi_gmem_WVALID,
	qsort_0_m_axi_gmem_WDATA,
	qsort_0_m_axi_gmem_WSTRB,
	qsort_0_m_axi_gmem_WLAST,
	qsort_0_m_axi_gmem_WUSER,
	qsort_0_m_axi_gmem_BREADY,
	qsort_0_m_axi_gmem_BVALID,
	qsort_0_m_axi_gmem_BID,
	qsort_0_m_axi_gmem_BRESP,
	qsort_0_m_axi_gmem_BUSER,
	qsort_0_s_axi_control_ARREADY,
	qsort_0_s_axi_control_ARVALID,
	qsort_0_s_axi_control_ARADDR,
	qsort_0_s_axi_control_RREADY,
	qsort_0_s_axi_control_RVALID,
	qsort_0_s_axi_control_RDATA,
	qsort_0_s_axi_control_RRESP,
	qsort_0_s_axi_control_AWREADY,
	qsort_0_s_axi_control_AWVALID,
	qsort_0_s_axi_control_AWADDR,
	qsort_0_s_axi_control_WREADY,
	qsort_0_s_axi_control_WVALID,
	qsort_0_s_axi_control_WDATA,
	qsort_0_s_axi_control_WSTRB,
	qsort_0_s_axi_control_BREADY,
	qsort_0_s_axi_control_BVALID,
	qsort_0_s_axi_control_BRESP,
	qsort_1_m_axi_gmem_ARREADY,
	qsort_1_m_axi_gmem_ARVALID,
	qsort_1_m_axi_gmem_ARID,
	qsort_1_m_axi_gmem_ARADDR,
	qsort_1_m_axi_gmem_ARLEN,
	qsort_1_m_axi_gmem_ARSIZE,
	qsort_1_m_axi_gmem_ARBURST,
	qsort_1_m_axi_gmem_ARLOCK,
	qsort_1_m_axi_gmem_ARCACHE,
	qsort_1_m_axi_gmem_ARPROT,
	qsort_1_m_axi_gmem_ARQOS,
	qsort_1_m_axi_gmem_ARREGION,
	qsort_1_m_axi_gmem_ARUSER,
	qsort_1_m_axi_gmem_RREADY,
	qsort_1_m_axi_gmem_RVALID,
	qsort_1_m_axi_gmem_RID,
	qsort_1_m_axi_gmem_RDATA,
	qsort_1_m_axi_gmem_RRESP,
	qsort_1_m_axi_gmem_RLAST,
	qsort_1_m_axi_gmem_RUSER,
	qsort_1_m_axi_gmem_AWREADY,
	qsort_1_m_axi_gmem_AWVALID,
	qsort_1_m_axi_gmem_AWID,
	qsort_1_m_axi_gmem_AWADDR,
	qsort_1_m_axi_gmem_AWLEN,
	qsort_1_m_axi_gmem_AWSIZE,
	qsort_1_m_axi_gmem_AWBURST,
	qsort_1_m_axi_gmem_AWLOCK,
	qsort_1_m_axi_gmem_AWCACHE,
	qsort_1_m_axi_gmem_AWPROT,
	qsort_1_m_axi_gmem_AWQOS,
	qsort_1_m_axi_gmem_AWREGION,
	qsort_1_m_axi_gmem_AWUSER,
	qsort_1_m_axi_gmem_WREADY,
	qsort_1_m_axi_gmem_WVALID,
	qsort_1_m_axi_gmem_WDATA,
	qsort_1_m_axi_gmem_WSTRB,
	qsort_1_m_axi_gmem_WLAST,
	qsort_1_m_axi_gmem_WUSER,
	qsort_1_m_axi_gmem_BREADY,
	qsort_1_m_axi_gmem_BVALID,
	qsort_1_m_axi_gmem_BID,
	qsort_1_m_axi_gmem_BRESP,
	qsort_1_m_axi_gmem_BUSER,
	qsort_1_s_axi_control_ARREADY,
	qsort_1_s_axi_control_ARVALID,
	qsort_1_s_axi_control_ARADDR,
	qsort_1_s_axi_control_RREADY,
	qsort_1_s_axi_control_RVALID,
	qsort_1_s_axi_control_RDATA,
	qsort_1_s_axi_control_RRESP,
	qsort_1_s_axi_control_AWREADY,
	qsort_1_s_axi_control_AWVALID,
	qsort_1_s_axi_control_AWADDR,
	qsort_1_s_axi_control_WREADY,
	qsort_1_s_axi_control_WVALID,
	qsort_1_s_axi_control_WDATA,
	qsort_1_s_axi_control_WSTRB,
	qsort_1_s_axi_control_BREADY,
	qsort_1_s_axi_control_BVALID,
	qsort_1_s_axi_control_BRESP,
	qsort_2_m_axi_gmem_ARREADY,
	qsort_2_m_axi_gmem_ARVALID,
	qsort_2_m_axi_gmem_ARID,
	qsort_2_m_axi_gmem_ARADDR,
	qsort_2_m_axi_gmem_ARLEN,
	qsort_2_m_axi_gmem_ARSIZE,
	qsort_2_m_axi_gmem_ARBURST,
	qsort_2_m_axi_gmem_ARLOCK,
	qsort_2_m_axi_gmem_ARCACHE,
	qsort_2_m_axi_gmem_ARPROT,
	qsort_2_m_axi_gmem_ARQOS,
	qsort_2_m_axi_gmem_ARREGION,
	qsort_2_m_axi_gmem_ARUSER,
	qsort_2_m_axi_gmem_RREADY,
	qsort_2_m_axi_gmem_RVALID,
	qsort_2_m_axi_gmem_RID,
	qsort_2_m_axi_gmem_RDATA,
	qsort_2_m_axi_gmem_RRESP,
	qsort_2_m_axi_gmem_RLAST,
	qsort_2_m_axi_gmem_RUSER,
	qsort_2_m_axi_gmem_AWREADY,
	qsort_2_m_axi_gmem_AWVALID,
	qsort_2_m_axi_gmem_AWID,
	qsort_2_m_axi_gmem_AWADDR,
	qsort_2_m_axi_gmem_AWLEN,
	qsort_2_m_axi_gmem_AWSIZE,
	qsort_2_m_axi_gmem_AWBURST,
	qsort_2_m_axi_gmem_AWLOCK,
	qsort_2_m_axi_gmem_AWCACHE,
	qsort_2_m_axi_gmem_AWPROT,
	qsort_2_m_axi_gmem_AWQOS,
	qsort_2_m_axi_gmem_AWREGION,
	qsort_2_m_axi_gmem_AWUSER,
	qsort_2_m_axi_gmem_WREADY,
	qsort_2_m_axi_gmem_WVALID,
	qsort_2_m_axi_gmem_WDATA,
	qsort_2_m_axi_gmem_WSTRB,
	qsort_2_m_axi_gmem_WLAST,
	qsort_2_m_axi_gmem_WUSER,
	qsort_2_m_axi_gmem_BREADY,
	qsort_2_m_axi_gmem_BVALID,
	qsort_2_m_axi_gmem_BID,
	qsort_2_m_axi_gmem_BRESP,
	qsort_2_m_axi_gmem_BUSER,
	qsort_2_s_axi_control_ARREADY,
	qsort_2_s_axi_control_ARVALID,
	qsort_2_s_axi_control_ARADDR,
	qsort_2_s_axi_control_RREADY,
	qsort_2_s_axi_control_RVALID,
	qsort_2_s_axi_control_RDATA,
	qsort_2_s_axi_control_RRESP,
	qsort_2_s_axi_control_AWREADY,
	qsort_2_s_axi_control_AWVALID,
	qsort_2_s_axi_control_AWADDR,
	qsort_2_s_axi_control_WREADY,
	qsort_2_s_axi_control_WVALID,
	qsort_2_s_axi_control_WDATA,
	qsort_2_s_axi_control_WSTRB,
	qsort_2_s_axi_control_BREADY,
	qsort_2_s_axi_control_BVALID,
	qsort_2_s_axi_control_BRESP,
	qsort_3_m_axi_gmem_ARREADY,
	qsort_3_m_axi_gmem_ARVALID,
	qsort_3_m_axi_gmem_ARID,
	qsort_3_m_axi_gmem_ARADDR,
	qsort_3_m_axi_gmem_ARLEN,
	qsort_3_m_axi_gmem_ARSIZE,
	qsort_3_m_axi_gmem_ARBURST,
	qsort_3_m_axi_gmem_ARLOCK,
	qsort_3_m_axi_gmem_ARCACHE,
	qsort_3_m_axi_gmem_ARPROT,
	qsort_3_m_axi_gmem_ARQOS,
	qsort_3_m_axi_gmem_ARREGION,
	qsort_3_m_axi_gmem_ARUSER,
	qsort_3_m_axi_gmem_RREADY,
	qsort_3_m_axi_gmem_RVALID,
	qsort_3_m_axi_gmem_RID,
	qsort_3_m_axi_gmem_RDATA,
	qsort_3_m_axi_gmem_RRESP,
	qsort_3_m_axi_gmem_RLAST,
	qsort_3_m_axi_gmem_RUSER,
	qsort_3_m_axi_gmem_AWREADY,
	qsort_3_m_axi_gmem_AWVALID,
	qsort_3_m_axi_gmem_AWID,
	qsort_3_m_axi_gmem_AWADDR,
	qsort_3_m_axi_gmem_AWLEN,
	qsort_3_m_axi_gmem_AWSIZE,
	qsort_3_m_axi_gmem_AWBURST,
	qsort_3_m_axi_gmem_AWLOCK,
	qsort_3_m_axi_gmem_AWCACHE,
	qsort_3_m_axi_gmem_AWPROT,
	qsort_3_m_axi_gmem_AWQOS,
	qsort_3_m_axi_gmem_AWREGION,
	qsort_3_m_axi_gmem_AWUSER,
	qsort_3_m_axi_gmem_WREADY,
	qsort_3_m_axi_gmem_WVALID,
	qsort_3_m_axi_gmem_WDATA,
	qsort_3_m_axi_gmem_WSTRB,
	qsort_3_m_axi_gmem_WLAST,
	qsort_3_m_axi_gmem_WUSER,
	qsort_3_m_axi_gmem_BREADY,
	qsort_3_m_axi_gmem_BVALID,
	qsort_3_m_axi_gmem_BID,
	qsort_3_m_axi_gmem_BRESP,
	qsort_3_m_axi_gmem_BUSER,
	qsort_3_s_axi_control_ARREADY,
	qsort_3_s_axi_control_ARVALID,
	qsort_3_s_axi_control_ARADDR,
	qsort_3_s_axi_control_RREADY,
	qsort_3_s_axi_control_RVALID,
	qsort_3_s_axi_control_RDATA,
	qsort_3_s_axi_control_RRESP,
	qsort_3_s_axi_control_AWREADY,
	qsort_3_s_axi_control_AWVALID,
	qsort_3_s_axi_control_AWADDR,
	qsort_3_s_axi_control_WREADY,
	qsort_3_s_axi_control_WVALID,
	qsort_3_s_axi_control_WDATA,
	qsort_3_s_axi_control_WSTRB,
	qsort_3_s_axi_control_BREADY,
	qsort_3_s_axi_control_BVALID,
	qsort_3_s_axi_control_BRESP,
	qsort_4_m_axi_gmem_ARREADY,
	qsort_4_m_axi_gmem_ARVALID,
	qsort_4_m_axi_gmem_ARID,
	qsort_4_m_axi_gmem_ARADDR,
	qsort_4_m_axi_gmem_ARLEN,
	qsort_4_m_axi_gmem_ARSIZE,
	qsort_4_m_axi_gmem_ARBURST,
	qsort_4_m_axi_gmem_ARLOCK,
	qsort_4_m_axi_gmem_ARCACHE,
	qsort_4_m_axi_gmem_ARPROT,
	qsort_4_m_axi_gmem_ARQOS,
	qsort_4_m_axi_gmem_ARREGION,
	qsort_4_m_axi_gmem_ARUSER,
	qsort_4_m_axi_gmem_RREADY,
	qsort_4_m_axi_gmem_RVALID,
	qsort_4_m_axi_gmem_RID,
	qsort_4_m_axi_gmem_RDATA,
	qsort_4_m_axi_gmem_RRESP,
	qsort_4_m_axi_gmem_RLAST,
	qsort_4_m_axi_gmem_RUSER,
	qsort_4_m_axi_gmem_AWREADY,
	qsort_4_m_axi_gmem_AWVALID,
	qsort_4_m_axi_gmem_AWID,
	qsort_4_m_axi_gmem_AWADDR,
	qsort_4_m_axi_gmem_AWLEN,
	qsort_4_m_axi_gmem_AWSIZE,
	qsort_4_m_axi_gmem_AWBURST,
	qsort_4_m_axi_gmem_AWLOCK,
	qsort_4_m_axi_gmem_AWCACHE,
	qsort_4_m_axi_gmem_AWPROT,
	qsort_4_m_axi_gmem_AWQOS,
	qsort_4_m_axi_gmem_AWREGION,
	qsort_4_m_axi_gmem_AWUSER,
	qsort_4_m_axi_gmem_WREADY,
	qsort_4_m_axi_gmem_WVALID,
	qsort_4_m_axi_gmem_WDATA,
	qsort_4_m_axi_gmem_WSTRB,
	qsort_4_m_axi_gmem_WLAST,
	qsort_4_m_axi_gmem_WUSER,
	qsort_4_m_axi_gmem_BREADY,
	qsort_4_m_axi_gmem_BVALID,
	qsort_4_m_axi_gmem_BID,
	qsort_4_m_axi_gmem_BRESP,
	qsort_4_m_axi_gmem_BUSER,
	qsort_4_s_axi_control_ARREADY,
	qsort_4_s_axi_control_ARVALID,
	qsort_4_s_axi_control_ARADDR,
	qsort_4_s_axi_control_RREADY,
	qsort_4_s_axi_control_RVALID,
	qsort_4_s_axi_control_RDATA,
	qsort_4_s_axi_control_RRESP,
	qsort_4_s_axi_control_AWREADY,
	qsort_4_s_axi_control_AWVALID,
	qsort_4_s_axi_control_AWADDR,
	qsort_4_s_axi_control_WREADY,
	qsort_4_s_axi_control_WVALID,
	qsort_4_s_axi_control_WDATA,
	qsort_4_s_axi_control_WSTRB,
	qsort_4_s_axi_control_BREADY,
	qsort_4_s_axi_control_BVALID,
	qsort_4_s_axi_control_BRESP,
	qsort_5_m_axi_gmem_ARREADY,
	qsort_5_m_axi_gmem_ARVALID,
	qsort_5_m_axi_gmem_ARID,
	qsort_5_m_axi_gmem_ARADDR,
	qsort_5_m_axi_gmem_ARLEN,
	qsort_5_m_axi_gmem_ARSIZE,
	qsort_5_m_axi_gmem_ARBURST,
	qsort_5_m_axi_gmem_ARLOCK,
	qsort_5_m_axi_gmem_ARCACHE,
	qsort_5_m_axi_gmem_ARPROT,
	qsort_5_m_axi_gmem_ARQOS,
	qsort_5_m_axi_gmem_ARREGION,
	qsort_5_m_axi_gmem_ARUSER,
	qsort_5_m_axi_gmem_RREADY,
	qsort_5_m_axi_gmem_RVALID,
	qsort_5_m_axi_gmem_RID,
	qsort_5_m_axi_gmem_RDATA,
	qsort_5_m_axi_gmem_RRESP,
	qsort_5_m_axi_gmem_RLAST,
	qsort_5_m_axi_gmem_RUSER,
	qsort_5_m_axi_gmem_AWREADY,
	qsort_5_m_axi_gmem_AWVALID,
	qsort_5_m_axi_gmem_AWID,
	qsort_5_m_axi_gmem_AWADDR,
	qsort_5_m_axi_gmem_AWLEN,
	qsort_5_m_axi_gmem_AWSIZE,
	qsort_5_m_axi_gmem_AWBURST,
	qsort_5_m_axi_gmem_AWLOCK,
	qsort_5_m_axi_gmem_AWCACHE,
	qsort_5_m_axi_gmem_AWPROT,
	qsort_5_m_axi_gmem_AWQOS,
	qsort_5_m_axi_gmem_AWREGION,
	qsort_5_m_axi_gmem_AWUSER,
	qsort_5_m_axi_gmem_WREADY,
	qsort_5_m_axi_gmem_WVALID,
	qsort_5_m_axi_gmem_WDATA,
	qsort_5_m_axi_gmem_WSTRB,
	qsort_5_m_axi_gmem_WLAST,
	qsort_5_m_axi_gmem_WUSER,
	qsort_5_m_axi_gmem_BREADY,
	qsort_5_m_axi_gmem_BVALID,
	qsort_5_m_axi_gmem_BID,
	qsort_5_m_axi_gmem_BRESP,
	qsort_5_m_axi_gmem_BUSER,
	qsort_5_s_axi_control_ARREADY,
	qsort_5_s_axi_control_ARVALID,
	qsort_5_s_axi_control_ARADDR,
	qsort_5_s_axi_control_RREADY,
	qsort_5_s_axi_control_RVALID,
	qsort_5_s_axi_control_RDATA,
	qsort_5_s_axi_control_RRESP,
	qsort_5_s_axi_control_AWREADY,
	qsort_5_s_axi_control_AWVALID,
	qsort_5_s_axi_control_AWADDR,
	qsort_5_s_axi_control_WREADY,
	qsort_5_s_axi_control_WVALID,
	qsort_5_s_axi_control_WDATA,
	qsort_5_s_axi_control_WSTRB,
	qsort_5_s_axi_control_BREADY,
	qsort_5_s_axi_control_BVALID,
	qsort_5_s_axi_control_BRESP,
	qsort_6_m_axi_gmem_ARREADY,
	qsort_6_m_axi_gmem_ARVALID,
	qsort_6_m_axi_gmem_ARID,
	qsort_6_m_axi_gmem_ARADDR,
	qsort_6_m_axi_gmem_ARLEN,
	qsort_6_m_axi_gmem_ARSIZE,
	qsort_6_m_axi_gmem_ARBURST,
	qsort_6_m_axi_gmem_ARLOCK,
	qsort_6_m_axi_gmem_ARCACHE,
	qsort_6_m_axi_gmem_ARPROT,
	qsort_6_m_axi_gmem_ARQOS,
	qsort_6_m_axi_gmem_ARREGION,
	qsort_6_m_axi_gmem_ARUSER,
	qsort_6_m_axi_gmem_RREADY,
	qsort_6_m_axi_gmem_RVALID,
	qsort_6_m_axi_gmem_RID,
	qsort_6_m_axi_gmem_RDATA,
	qsort_6_m_axi_gmem_RRESP,
	qsort_6_m_axi_gmem_RLAST,
	qsort_6_m_axi_gmem_RUSER,
	qsort_6_m_axi_gmem_AWREADY,
	qsort_6_m_axi_gmem_AWVALID,
	qsort_6_m_axi_gmem_AWID,
	qsort_6_m_axi_gmem_AWADDR,
	qsort_6_m_axi_gmem_AWLEN,
	qsort_6_m_axi_gmem_AWSIZE,
	qsort_6_m_axi_gmem_AWBURST,
	qsort_6_m_axi_gmem_AWLOCK,
	qsort_6_m_axi_gmem_AWCACHE,
	qsort_6_m_axi_gmem_AWPROT,
	qsort_6_m_axi_gmem_AWQOS,
	qsort_6_m_axi_gmem_AWREGION,
	qsort_6_m_axi_gmem_AWUSER,
	qsort_6_m_axi_gmem_WREADY,
	qsort_6_m_axi_gmem_WVALID,
	qsort_6_m_axi_gmem_WDATA,
	qsort_6_m_axi_gmem_WSTRB,
	qsort_6_m_axi_gmem_WLAST,
	qsort_6_m_axi_gmem_WUSER,
	qsort_6_m_axi_gmem_BREADY,
	qsort_6_m_axi_gmem_BVALID,
	qsort_6_m_axi_gmem_BID,
	qsort_6_m_axi_gmem_BRESP,
	qsort_6_m_axi_gmem_BUSER,
	qsort_6_s_axi_control_ARREADY,
	qsort_6_s_axi_control_ARVALID,
	qsort_6_s_axi_control_ARADDR,
	qsort_6_s_axi_control_RREADY,
	qsort_6_s_axi_control_RVALID,
	qsort_6_s_axi_control_RDATA,
	qsort_6_s_axi_control_RRESP,
	qsort_6_s_axi_control_AWREADY,
	qsort_6_s_axi_control_AWVALID,
	qsort_6_s_axi_control_AWADDR,
	qsort_6_s_axi_control_WREADY,
	qsort_6_s_axi_control_WVALID,
	qsort_6_s_axi_control_WDATA,
	qsort_6_s_axi_control_WSTRB,
	qsort_6_s_axi_control_BREADY,
	qsort_6_s_axi_control_BVALID,
	qsort_6_s_axi_control_BRESP,
	qsort_7_m_axi_gmem_ARREADY,
	qsort_7_m_axi_gmem_ARVALID,
	qsort_7_m_axi_gmem_ARID,
	qsort_7_m_axi_gmem_ARADDR,
	qsort_7_m_axi_gmem_ARLEN,
	qsort_7_m_axi_gmem_ARSIZE,
	qsort_7_m_axi_gmem_ARBURST,
	qsort_7_m_axi_gmem_ARLOCK,
	qsort_7_m_axi_gmem_ARCACHE,
	qsort_7_m_axi_gmem_ARPROT,
	qsort_7_m_axi_gmem_ARQOS,
	qsort_7_m_axi_gmem_ARREGION,
	qsort_7_m_axi_gmem_ARUSER,
	qsort_7_m_axi_gmem_RREADY,
	qsort_7_m_axi_gmem_RVALID,
	qsort_7_m_axi_gmem_RID,
	qsort_7_m_axi_gmem_RDATA,
	qsort_7_m_axi_gmem_RRESP,
	qsort_7_m_axi_gmem_RLAST,
	qsort_7_m_axi_gmem_RUSER,
	qsort_7_m_axi_gmem_AWREADY,
	qsort_7_m_axi_gmem_AWVALID,
	qsort_7_m_axi_gmem_AWID,
	qsort_7_m_axi_gmem_AWADDR,
	qsort_7_m_axi_gmem_AWLEN,
	qsort_7_m_axi_gmem_AWSIZE,
	qsort_7_m_axi_gmem_AWBURST,
	qsort_7_m_axi_gmem_AWLOCK,
	qsort_7_m_axi_gmem_AWCACHE,
	qsort_7_m_axi_gmem_AWPROT,
	qsort_7_m_axi_gmem_AWQOS,
	qsort_7_m_axi_gmem_AWREGION,
	qsort_7_m_axi_gmem_AWUSER,
	qsort_7_m_axi_gmem_WREADY,
	qsort_7_m_axi_gmem_WVALID,
	qsort_7_m_axi_gmem_WDATA,
	qsort_7_m_axi_gmem_WSTRB,
	qsort_7_m_axi_gmem_WLAST,
	qsort_7_m_axi_gmem_WUSER,
	qsort_7_m_axi_gmem_BREADY,
	qsort_7_m_axi_gmem_BVALID,
	qsort_7_m_axi_gmem_BID,
	qsort_7_m_axi_gmem_BRESP,
	qsort_7_m_axi_gmem_BUSER,
	qsort_7_s_axi_control_ARREADY,
	qsort_7_s_axi_control_ARVALID,
	qsort_7_s_axi_control_ARADDR,
	qsort_7_s_axi_control_RREADY,
	qsort_7_s_axi_control_RVALID,
	qsort_7_s_axi_control_RDATA,
	qsort_7_s_axi_control_RRESP,
	qsort_7_s_axi_control_AWREADY,
	qsort_7_s_axi_control_AWVALID,
	qsort_7_s_axi_control_AWADDR,
	qsort_7_s_axi_control_WREADY,
	qsort_7_s_axi_control_WVALID,
	qsort_7_s_axi_control_WDATA,
	qsort_7_s_axi_control_WSTRB,
	qsort_7_s_axi_control_BREADY,
	qsort_7_s_axi_control_BVALID,
	qsort_7_s_axi_control_BRESP,
	qsort_8_m_axi_gmem_ARREADY,
	qsort_8_m_axi_gmem_ARVALID,
	qsort_8_m_axi_gmem_ARID,
	qsort_8_m_axi_gmem_ARADDR,
	qsort_8_m_axi_gmem_ARLEN,
	qsort_8_m_axi_gmem_ARSIZE,
	qsort_8_m_axi_gmem_ARBURST,
	qsort_8_m_axi_gmem_ARLOCK,
	qsort_8_m_axi_gmem_ARCACHE,
	qsort_8_m_axi_gmem_ARPROT,
	qsort_8_m_axi_gmem_ARQOS,
	qsort_8_m_axi_gmem_ARREGION,
	qsort_8_m_axi_gmem_ARUSER,
	qsort_8_m_axi_gmem_RREADY,
	qsort_8_m_axi_gmem_RVALID,
	qsort_8_m_axi_gmem_RID,
	qsort_8_m_axi_gmem_RDATA,
	qsort_8_m_axi_gmem_RRESP,
	qsort_8_m_axi_gmem_RLAST,
	qsort_8_m_axi_gmem_RUSER,
	qsort_8_m_axi_gmem_AWREADY,
	qsort_8_m_axi_gmem_AWVALID,
	qsort_8_m_axi_gmem_AWID,
	qsort_8_m_axi_gmem_AWADDR,
	qsort_8_m_axi_gmem_AWLEN,
	qsort_8_m_axi_gmem_AWSIZE,
	qsort_8_m_axi_gmem_AWBURST,
	qsort_8_m_axi_gmem_AWLOCK,
	qsort_8_m_axi_gmem_AWCACHE,
	qsort_8_m_axi_gmem_AWPROT,
	qsort_8_m_axi_gmem_AWQOS,
	qsort_8_m_axi_gmem_AWREGION,
	qsort_8_m_axi_gmem_AWUSER,
	qsort_8_m_axi_gmem_WREADY,
	qsort_8_m_axi_gmem_WVALID,
	qsort_8_m_axi_gmem_WDATA,
	qsort_8_m_axi_gmem_WSTRB,
	qsort_8_m_axi_gmem_WLAST,
	qsort_8_m_axi_gmem_WUSER,
	qsort_8_m_axi_gmem_BREADY,
	qsort_8_m_axi_gmem_BVALID,
	qsort_8_m_axi_gmem_BID,
	qsort_8_m_axi_gmem_BRESP,
	qsort_8_m_axi_gmem_BUSER,
	qsort_8_s_axi_control_ARREADY,
	qsort_8_s_axi_control_ARVALID,
	qsort_8_s_axi_control_ARADDR,
	qsort_8_s_axi_control_RREADY,
	qsort_8_s_axi_control_RVALID,
	qsort_8_s_axi_control_RDATA,
	qsort_8_s_axi_control_RRESP,
	qsort_8_s_axi_control_AWREADY,
	qsort_8_s_axi_control_AWVALID,
	qsort_8_s_axi_control_AWADDR,
	qsort_8_s_axi_control_WREADY,
	qsort_8_s_axi_control_WVALID,
	qsort_8_s_axi_control_WDATA,
	qsort_8_s_axi_control_WSTRB,
	qsort_8_s_axi_control_BREADY,
	qsort_8_s_axi_control_BVALID,
	qsort_8_s_axi_control_BRESP,
	qsort_9_m_axi_gmem_ARREADY,
	qsort_9_m_axi_gmem_ARVALID,
	qsort_9_m_axi_gmem_ARID,
	qsort_9_m_axi_gmem_ARADDR,
	qsort_9_m_axi_gmem_ARLEN,
	qsort_9_m_axi_gmem_ARSIZE,
	qsort_9_m_axi_gmem_ARBURST,
	qsort_9_m_axi_gmem_ARLOCK,
	qsort_9_m_axi_gmem_ARCACHE,
	qsort_9_m_axi_gmem_ARPROT,
	qsort_9_m_axi_gmem_ARQOS,
	qsort_9_m_axi_gmem_ARREGION,
	qsort_9_m_axi_gmem_ARUSER,
	qsort_9_m_axi_gmem_RREADY,
	qsort_9_m_axi_gmem_RVALID,
	qsort_9_m_axi_gmem_RID,
	qsort_9_m_axi_gmem_RDATA,
	qsort_9_m_axi_gmem_RRESP,
	qsort_9_m_axi_gmem_RLAST,
	qsort_9_m_axi_gmem_RUSER,
	qsort_9_m_axi_gmem_AWREADY,
	qsort_9_m_axi_gmem_AWVALID,
	qsort_9_m_axi_gmem_AWID,
	qsort_9_m_axi_gmem_AWADDR,
	qsort_9_m_axi_gmem_AWLEN,
	qsort_9_m_axi_gmem_AWSIZE,
	qsort_9_m_axi_gmem_AWBURST,
	qsort_9_m_axi_gmem_AWLOCK,
	qsort_9_m_axi_gmem_AWCACHE,
	qsort_9_m_axi_gmem_AWPROT,
	qsort_9_m_axi_gmem_AWQOS,
	qsort_9_m_axi_gmem_AWREGION,
	qsort_9_m_axi_gmem_AWUSER,
	qsort_9_m_axi_gmem_WREADY,
	qsort_9_m_axi_gmem_WVALID,
	qsort_9_m_axi_gmem_WDATA,
	qsort_9_m_axi_gmem_WSTRB,
	qsort_9_m_axi_gmem_WLAST,
	qsort_9_m_axi_gmem_WUSER,
	qsort_9_m_axi_gmem_BREADY,
	qsort_9_m_axi_gmem_BVALID,
	qsort_9_m_axi_gmem_BID,
	qsort_9_m_axi_gmem_BRESP,
	qsort_9_m_axi_gmem_BUSER,
	qsort_9_s_axi_control_ARREADY,
	qsort_9_s_axi_control_ARVALID,
	qsort_9_s_axi_control_ARADDR,
	qsort_9_s_axi_control_RREADY,
	qsort_9_s_axi_control_RVALID,
	qsort_9_s_axi_control_RDATA,
	qsort_9_s_axi_control_RRESP,
	qsort_9_s_axi_control_AWREADY,
	qsort_9_s_axi_control_AWVALID,
	qsort_9_s_axi_control_AWADDR,
	qsort_9_s_axi_control_WREADY,
	qsort_9_s_axi_control_WVALID,
	qsort_9_s_axi_control_WDATA,
	qsort_9_s_axi_control_WSTRB,
	qsort_9_s_axi_control_BREADY,
	qsort_9_s_axi_control_BVALID,
	qsort_9_s_axi_control_BRESP,
	qsort_10_m_axi_gmem_ARREADY,
	qsort_10_m_axi_gmem_ARVALID,
	qsort_10_m_axi_gmem_ARID,
	qsort_10_m_axi_gmem_ARADDR,
	qsort_10_m_axi_gmem_ARLEN,
	qsort_10_m_axi_gmem_ARSIZE,
	qsort_10_m_axi_gmem_ARBURST,
	qsort_10_m_axi_gmem_ARLOCK,
	qsort_10_m_axi_gmem_ARCACHE,
	qsort_10_m_axi_gmem_ARPROT,
	qsort_10_m_axi_gmem_ARQOS,
	qsort_10_m_axi_gmem_ARREGION,
	qsort_10_m_axi_gmem_ARUSER,
	qsort_10_m_axi_gmem_RREADY,
	qsort_10_m_axi_gmem_RVALID,
	qsort_10_m_axi_gmem_RID,
	qsort_10_m_axi_gmem_RDATA,
	qsort_10_m_axi_gmem_RRESP,
	qsort_10_m_axi_gmem_RLAST,
	qsort_10_m_axi_gmem_RUSER,
	qsort_10_m_axi_gmem_AWREADY,
	qsort_10_m_axi_gmem_AWVALID,
	qsort_10_m_axi_gmem_AWID,
	qsort_10_m_axi_gmem_AWADDR,
	qsort_10_m_axi_gmem_AWLEN,
	qsort_10_m_axi_gmem_AWSIZE,
	qsort_10_m_axi_gmem_AWBURST,
	qsort_10_m_axi_gmem_AWLOCK,
	qsort_10_m_axi_gmem_AWCACHE,
	qsort_10_m_axi_gmem_AWPROT,
	qsort_10_m_axi_gmem_AWQOS,
	qsort_10_m_axi_gmem_AWREGION,
	qsort_10_m_axi_gmem_AWUSER,
	qsort_10_m_axi_gmem_WREADY,
	qsort_10_m_axi_gmem_WVALID,
	qsort_10_m_axi_gmem_WDATA,
	qsort_10_m_axi_gmem_WSTRB,
	qsort_10_m_axi_gmem_WLAST,
	qsort_10_m_axi_gmem_WUSER,
	qsort_10_m_axi_gmem_BREADY,
	qsort_10_m_axi_gmem_BVALID,
	qsort_10_m_axi_gmem_BID,
	qsort_10_m_axi_gmem_BRESP,
	qsort_10_m_axi_gmem_BUSER,
	qsort_10_s_axi_control_ARREADY,
	qsort_10_s_axi_control_ARVALID,
	qsort_10_s_axi_control_ARADDR,
	qsort_10_s_axi_control_RREADY,
	qsort_10_s_axi_control_RVALID,
	qsort_10_s_axi_control_RDATA,
	qsort_10_s_axi_control_RRESP,
	qsort_10_s_axi_control_AWREADY,
	qsort_10_s_axi_control_AWVALID,
	qsort_10_s_axi_control_AWADDR,
	qsort_10_s_axi_control_WREADY,
	qsort_10_s_axi_control_WVALID,
	qsort_10_s_axi_control_WDATA,
	qsort_10_s_axi_control_WSTRB,
	qsort_10_s_axi_control_BREADY,
	qsort_10_s_axi_control_BVALID,
	qsort_10_s_axi_control_BRESP,
	qsort_11_m_axi_gmem_ARREADY,
	qsort_11_m_axi_gmem_ARVALID,
	qsort_11_m_axi_gmem_ARID,
	qsort_11_m_axi_gmem_ARADDR,
	qsort_11_m_axi_gmem_ARLEN,
	qsort_11_m_axi_gmem_ARSIZE,
	qsort_11_m_axi_gmem_ARBURST,
	qsort_11_m_axi_gmem_ARLOCK,
	qsort_11_m_axi_gmem_ARCACHE,
	qsort_11_m_axi_gmem_ARPROT,
	qsort_11_m_axi_gmem_ARQOS,
	qsort_11_m_axi_gmem_ARREGION,
	qsort_11_m_axi_gmem_ARUSER,
	qsort_11_m_axi_gmem_RREADY,
	qsort_11_m_axi_gmem_RVALID,
	qsort_11_m_axi_gmem_RID,
	qsort_11_m_axi_gmem_RDATA,
	qsort_11_m_axi_gmem_RRESP,
	qsort_11_m_axi_gmem_RLAST,
	qsort_11_m_axi_gmem_RUSER,
	qsort_11_m_axi_gmem_AWREADY,
	qsort_11_m_axi_gmem_AWVALID,
	qsort_11_m_axi_gmem_AWID,
	qsort_11_m_axi_gmem_AWADDR,
	qsort_11_m_axi_gmem_AWLEN,
	qsort_11_m_axi_gmem_AWSIZE,
	qsort_11_m_axi_gmem_AWBURST,
	qsort_11_m_axi_gmem_AWLOCK,
	qsort_11_m_axi_gmem_AWCACHE,
	qsort_11_m_axi_gmem_AWPROT,
	qsort_11_m_axi_gmem_AWQOS,
	qsort_11_m_axi_gmem_AWREGION,
	qsort_11_m_axi_gmem_AWUSER,
	qsort_11_m_axi_gmem_WREADY,
	qsort_11_m_axi_gmem_WVALID,
	qsort_11_m_axi_gmem_WDATA,
	qsort_11_m_axi_gmem_WSTRB,
	qsort_11_m_axi_gmem_WLAST,
	qsort_11_m_axi_gmem_WUSER,
	qsort_11_m_axi_gmem_BREADY,
	qsort_11_m_axi_gmem_BVALID,
	qsort_11_m_axi_gmem_BID,
	qsort_11_m_axi_gmem_BRESP,
	qsort_11_m_axi_gmem_BUSER,
	qsort_11_s_axi_control_ARREADY,
	qsort_11_s_axi_control_ARVALID,
	qsort_11_s_axi_control_ARADDR,
	qsort_11_s_axi_control_RREADY,
	qsort_11_s_axi_control_RVALID,
	qsort_11_s_axi_control_RDATA,
	qsort_11_s_axi_control_RRESP,
	qsort_11_s_axi_control_AWREADY,
	qsort_11_s_axi_control_AWVALID,
	qsort_11_s_axi_control_AWADDR,
	qsort_11_s_axi_control_WREADY,
	qsort_11_s_axi_control_WVALID,
	qsort_11_s_axi_control_WDATA,
	qsort_11_s_axi_control_WSTRB,
	qsort_11_s_axi_control_BREADY,
	qsort_11_s_axi_control_BVALID,
	qsort_11_s_axi_control_BRESP,
	qsort_12_m_axi_gmem_ARREADY,
	qsort_12_m_axi_gmem_ARVALID,
	qsort_12_m_axi_gmem_ARID,
	qsort_12_m_axi_gmem_ARADDR,
	qsort_12_m_axi_gmem_ARLEN,
	qsort_12_m_axi_gmem_ARSIZE,
	qsort_12_m_axi_gmem_ARBURST,
	qsort_12_m_axi_gmem_ARLOCK,
	qsort_12_m_axi_gmem_ARCACHE,
	qsort_12_m_axi_gmem_ARPROT,
	qsort_12_m_axi_gmem_ARQOS,
	qsort_12_m_axi_gmem_ARREGION,
	qsort_12_m_axi_gmem_ARUSER,
	qsort_12_m_axi_gmem_RREADY,
	qsort_12_m_axi_gmem_RVALID,
	qsort_12_m_axi_gmem_RID,
	qsort_12_m_axi_gmem_RDATA,
	qsort_12_m_axi_gmem_RRESP,
	qsort_12_m_axi_gmem_RLAST,
	qsort_12_m_axi_gmem_RUSER,
	qsort_12_m_axi_gmem_AWREADY,
	qsort_12_m_axi_gmem_AWVALID,
	qsort_12_m_axi_gmem_AWID,
	qsort_12_m_axi_gmem_AWADDR,
	qsort_12_m_axi_gmem_AWLEN,
	qsort_12_m_axi_gmem_AWSIZE,
	qsort_12_m_axi_gmem_AWBURST,
	qsort_12_m_axi_gmem_AWLOCK,
	qsort_12_m_axi_gmem_AWCACHE,
	qsort_12_m_axi_gmem_AWPROT,
	qsort_12_m_axi_gmem_AWQOS,
	qsort_12_m_axi_gmem_AWREGION,
	qsort_12_m_axi_gmem_AWUSER,
	qsort_12_m_axi_gmem_WREADY,
	qsort_12_m_axi_gmem_WVALID,
	qsort_12_m_axi_gmem_WDATA,
	qsort_12_m_axi_gmem_WSTRB,
	qsort_12_m_axi_gmem_WLAST,
	qsort_12_m_axi_gmem_WUSER,
	qsort_12_m_axi_gmem_BREADY,
	qsort_12_m_axi_gmem_BVALID,
	qsort_12_m_axi_gmem_BID,
	qsort_12_m_axi_gmem_BRESP,
	qsort_12_m_axi_gmem_BUSER,
	qsort_12_s_axi_control_ARREADY,
	qsort_12_s_axi_control_ARVALID,
	qsort_12_s_axi_control_ARADDR,
	qsort_12_s_axi_control_RREADY,
	qsort_12_s_axi_control_RVALID,
	qsort_12_s_axi_control_RDATA,
	qsort_12_s_axi_control_RRESP,
	qsort_12_s_axi_control_AWREADY,
	qsort_12_s_axi_control_AWVALID,
	qsort_12_s_axi_control_AWADDR,
	qsort_12_s_axi_control_WREADY,
	qsort_12_s_axi_control_WVALID,
	qsort_12_s_axi_control_WDATA,
	qsort_12_s_axi_control_WSTRB,
	qsort_12_s_axi_control_BREADY,
	qsort_12_s_axi_control_BVALID,
	qsort_12_s_axi_control_BRESP,
	qsort_13_m_axi_gmem_ARREADY,
	qsort_13_m_axi_gmem_ARVALID,
	qsort_13_m_axi_gmem_ARID,
	qsort_13_m_axi_gmem_ARADDR,
	qsort_13_m_axi_gmem_ARLEN,
	qsort_13_m_axi_gmem_ARSIZE,
	qsort_13_m_axi_gmem_ARBURST,
	qsort_13_m_axi_gmem_ARLOCK,
	qsort_13_m_axi_gmem_ARCACHE,
	qsort_13_m_axi_gmem_ARPROT,
	qsort_13_m_axi_gmem_ARQOS,
	qsort_13_m_axi_gmem_ARREGION,
	qsort_13_m_axi_gmem_ARUSER,
	qsort_13_m_axi_gmem_RREADY,
	qsort_13_m_axi_gmem_RVALID,
	qsort_13_m_axi_gmem_RID,
	qsort_13_m_axi_gmem_RDATA,
	qsort_13_m_axi_gmem_RRESP,
	qsort_13_m_axi_gmem_RLAST,
	qsort_13_m_axi_gmem_RUSER,
	qsort_13_m_axi_gmem_AWREADY,
	qsort_13_m_axi_gmem_AWVALID,
	qsort_13_m_axi_gmem_AWID,
	qsort_13_m_axi_gmem_AWADDR,
	qsort_13_m_axi_gmem_AWLEN,
	qsort_13_m_axi_gmem_AWSIZE,
	qsort_13_m_axi_gmem_AWBURST,
	qsort_13_m_axi_gmem_AWLOCK,
	qsort_13_m_axi_gmem_AWCACHE,
	qsort_13_m_axi_gmem_AWPROT,
	qsort_13_m_axi_gmem_AWQOS,
	qsort_13_m_axi_gmem_AWREGION,
	qsort_13_m_axi_gmem_AWUSER,
	qsort_13_m_axi_gmem_WREADY,
	qsort_13_m_axi_gmem_WVALID,
	qsort_13_m_axi_gmem_WDATA,
	qsort_13_m_axi_gmem_WSTRB,
	qsort_13_m_axi_gmem_WLAST,
	qsort_13_m_axi_gmem_WUSER,
	qsort_13_m_axi_gmem_BREADY,
	qsort_13_m_axi_gmem_BVALID,
	qsort_13_m_axi_gmem_BID,
	qsort_13_m_axi_gmem_BRESP,
	qsort_13_m_axi_gmem_BUSER,
	qsort_13_s_axi_control_ARREADY,
	qsort_13_s_axi_control_ARVALID,
	qsort_13_s_axi_control_ARADDR,
	qsort_13_s_axi_control_RREADY,
	qsort_13_s_axi_control_RVALID,
	qsort_13_s_axi_control_RDATA,
	qsort_13_s_axi_control_RRESP,
	qsort_13_s_axi_control_AWREADY,
	qsort_13_s_axi_control_AWVALID,
	qsort_13_s_axi_control_AWADDR,
	qsort_13_s_axi_control_WREADY,
	qsort_13_s_axi_control_WVALID,
	qsort_13_s_axi_control_WDATA,
	qsort_13_s_axi_control_WSTRB,
	qsort_13_s_axi_control_BREADY,
	qsort_13_s_axi_control_BVALID,
	qsort_13_s_axi_control_BRESP,
	qsort_14_m_axi_gmem_ARREADY,
	qsort_14_m_axi_gmem_ARVALID,
	qsort_14_m_axi_gmem_ARID,
	qsort_14_m_axi_gmem_ARADDR,
	qsort_14_m_axi_gmem_ARLEN,
	qsort_14_m_axi_gmem_ARSIZE,
	qsort_14_m_axi_gmem_ARBURST,
	qsort_14_m_axi_gmem_ARLOCK,
	qsort_14_m_axi_gmem_ARCACHE,
	qsort_14_m_axi_gmem_ARPROT,
	qsort_14_m_axi_gmem_ARQOS,
	qsort_14_m_axi_gmem_ARREGION,
	qsort_14_m_axi_gmem_ARUSER,
	qsort_14_m_axi_gmem_RREADY,
	qsort_14_m_axi_gmem_RVALID,
	qsort_14_m_axi_gmem_RID,
	qsort_14_m_axi_gmem_RDATA,
	qsort_14_m_axi_gmem_RRESP,
	qsort_14_m_axi_gmem_RLAST,
	qsort_14_m_axi_gmem_RUSER,
	qsort_14_m_axi_gmem_AWREADY,
	qsort_14_m_axi_gmem_AWVALID,
	qsort_14_m_axi_gmem_AWID,
	qsort_14_m_axi_gmem_AWADDR,
	qsort_14_m_axi_gmem_AWLEN,
	qsort_14_m_axi_gmem_AWSIZE,
	qsort_14_m_axi_gmem_AWBURST,
	qsort_14_m_axi_gmem_AWLOCK,
	qsort_14_m_axi_gmem_AWCACHE,
	qsort_14_m_axi_gmem_AWPROT,
	qsort_14_m_axi_gmem_AWQOS,
	qsort_14_m_axi_gmem_AWREGION,
	qsort_14_m_axi_gmem_AWUSER,
	qsort_14_m_axi_gmem_WREADY,
	qsort_14_m_axi_gmem_WVALID,
	qsort_14_m_axi_gmem_WDATA,
	qsort_14_m_axi_gmem_WSTRB,
	qsort_14_m_axi_gmem_WLAST,
	qsort_14_m_axi_gmem_WUSER,
	qsort_14_m_axi_gmem_BREADY,
	qsort_14_m_axi_gmem_BVALID,
	qsort_14_m_axi_gmem_BID,
	qsort_14_m_axi_gmem_BRESP,
	qsort_14_m_axi_gmem_BUSER,
	qsort_14_s_axi_control_ARREADY,
	qsort_14_s_axi_control_ARVALID,
	qsort_14_s_axi_control_ARADDR,
	qsort_14_s_axi_control_RREADY,
	qsort_14_s_axi_control_RVALID,
	qsort_14_s_axi_control_RDATA,
	qsort_14_s_axi_control_RRESP,
	qsort_14_s_axi_control_AWREADY,
	qsort_14_s_axi_control_AWVALID,
	qsort_14_s_axi_control_AWADDR,
	qsort_14_s_axi_control_WREADY,
	qsort_14_s_axi_control_WVALID,
	qsort_14_s_axi_control_WDATA,
	qsort_14_s_axi_control_WSTRB,
	qsort_14_s_axi_control_BREADY,
	qsort_14_s_axi_control_BVALID,
	qsort_14_s_axi_control_BRESP,
	qsort_15_m_axi_gmem_ARREADY,
	qsort_15_m_axi_gmem_ARVALID,
	qsort_15_m_axi_gmem_ARID,
	qsort_15_m_axi_gmem_ARADDR,
	qsort_15_m_axi_gmem_ARLEN,
	qsort_15_m_axi_gmem_ARSIZE,
	qsort_15_m_axi_gmem_ARBURST,
	qsort_15_m_axi_gmem_ARLOCK,
	qsort_15_m_axi_gmem_ARCACHE,
	qsort_15_m_axi_gmem_ARPROT,
	qsort_15_m_axi_gmem_ARQOS,
	qsort_15_m_axi_gmem_ARREGION,
	qsort_15_m_axi_gmem_ARUSER,
	qsort_15_m_axi_gmem_RREADY,
	qsort_15_m_axi_gmem_RVALID,
	qsort_15_m_axi_gmem_RID,
	qsort_15_m_axi_gmem_RDATA,
	qsort_15_m_axi_gmem_RRESP,
	qsort_15_m_axi_gmem_RLAST,
	qsort_15_m_axi_gmem_RUSER,
	qsort_15_m_axi_gmem_AWREADY,
	qsort_15_m_axi_gmem_AWVALID,
	qsort_15_m_axi_gmem_AWID,
	qsort_15_m_axi_gmem_AWADDR,
	qsort_15_m_axi_gmem_AWLEN,
	qsort_15_m_axi_gmem_AWSIZE,
	qsort_15_m_axi_gmem_AWBURST,
	qsort_15_m_axi_gmem_AWLOCK,
	qsort_15_m_axi_gmem_AWCACHE,
	qsort_15_m_axi_gmem_AWPROT,
	qsort_15_m_axi_gmem_AWQOS,
	qsort_15_m_axi_gmem_AWREGION,
	qsort_15_m_axi_gmem_AWUSER,
	qsort_15_m_axi_gmem_WREADY,
	qsort_15_m_axi_gmem_WVALID,
	qsort_15_m_axi_gmem_WDATA,
	qsort_15_m_axi_gmem_WSTRB,
	qsort_15_m_axi_gmem_WLAST,
	qsort_15_m_axi_gmem_WUSER,
	qsort_15_m_axi_gmem_BREADY,
	qsort_15_m_axi_gmem_BVALID,
	qsort_15_m_axi_gmem_BID,
	qsort_15_m_axi_gmem_BRESP,
	qsort_15_m_axi_gmem_BUSER,
	qsort_15_s_axi_control_ARREADY,
	qsort_15_s_axi_control_ARVALID,
	qsort_15_s_axi_control_ARADDR,
	qsort_15_s_axi_control_RREADY,
	qsort_15_s_axi_control_RVALID,
	qsort_15_s_axi_control_RDATA,
	qsort_15_s_axi_control_RRESP,
	qsort_15_s_axi_control_AWREADY,
	qsort_15_s_axi_control_AWVALID,
	qsort_15_s_axi_control_AWADDR,
	qsort_15_s_axi_control_WREADY,
	qsort_15_s_axi_control_WVALID,
	qsort_15_s_axi_control_WDATA,
	qsort_15_s_axi_control_WSTRB,
	qsort_15_s_axi_control_BREADY,
	qsort_15_s_axi_control_BVALID,
	qsort_15_s_axi_control_BRESP,
	qsort_16_m_axi_gmem_ARREADY,
	qsort_16_m_axi_gmem_ARVALID,
	qsort_16_m_axi_gmem_ARID,
	qsort_16_m_axi_gmem_ARADDR,
	qsort_16_m_axi_gmem_ARLEN,
	qsort_16_m_axi_gmem_ARSIZE,
	qsort_16_m_axi_gmem_ARBURST,
	qsort_16_m_axi_gmem_ARLOCK,
	qsort_16_m_axi_gmem_ARCACHE,
	qsort_16_m_axi_gmem_ARPROT,
	qsort_16_m_axi_gmem_ARQOS,
	qsort_16_m_axi_gmem_ARREGION,
	qsort_16_m_axi_gmem_ARUSER,
	qsort_16_m_axi_gmem_RREADY,
	qsort_16_m_axi_gmem_RVALID,
	qsort_16_m_axi_gmem_RID,
	qsort_16_m_axi_gmem_RDATA,
	qsort_16_m_axi_gmem_RRESP,
	qsort_16_m_axi_gmem_RLAST,
	qsort_16_m_axi_gmem_RUSER,
	qsort_16_m_axi_gmem_AWREADY,
	qsort_16_m_axi_gmem_AWVALID,
	qsort_16_m_axi_gmem_AWID,
	qsort_16_m_axi_gmem_AWADDR,
	qsort_16_m_axi_gmem_AWLEN,
	qsort_16_m_axi_gmem_AWSIZE,
	qsort_16_m_axi_gmem_AWBURST,
	qsort_16_m_axi_gmem_AWLOCK,
	qsort_16_m_axi_gmem_AWCACHE,
	qsort_16_m_axi_gmem_AWPROT,
	qsort_16_m_axi_gmem_AWQOS,
	qsort_16_m_axi_gmem_AWREGION,
	qsort_16_m_axi_gmem_AWUSER,
	qsort_16_m_axi_gmem_WREADY,
	qsort_16_m_axi_gmem_WVALID,
	qsort_16_m_axi_gmem_WDATA,
	qsort_16_m_axi_gmem_WSTRB,
	qsort_16_m_axi_gmem_WLAST,
	qsort_16_m_axi_gmem_WUSER,
	qsort_16_m_axi_gmem_BREADY,
	qsort_16_m_axi_gmem_BVALID,
	qsort_16_m_axi_gmem_BID,
	qsort_16_m_axi_gmem_BRESP,
	qsort_16_m_axi_gmem_BUSER,
	qsort_16_s_axi_control_ARREADY,
	qsort_16_s_axi_control_ARVALID,
	qsort_16_s_axi_control_ARADDR,
	qsort_16_s_axi_control_RREADY,
	qsort_16_s_axi_control_RVALID,
	qsort_16_s_axi_control_RDATA,
	qsort_16_s_axi_control_RRESP,
	qsort_16_s_axi_control_AWREADY,
	qsort_16_s_axi_control_AWVALID,
	qsort_16_s_axi_control_AWADDR,
	qsort_16_s_axi_control_WREADY,
	qsort_16_s_axi_control_WVALID,
	qsort_16_s_axi_control_WDATA,
	qsort_16_s_axi_control_WSTRB,
	qsort_16_s_axi_control_BREADY,
	qsort_16_s_axi_control_BVALID,
	qsort_16_s_axi_control_BRESP,
	qsort_17_m_axi_gmem_ARREADY,
	qsort_17_m_axi_gmem_ARVALID,
	qsort_17_m_axi_gmem_ARID,
	qsort_17_m_axi_gmem_ARADDR,
	qsort_17_m_axi_gmem_ARLEN,
	qsort_17_m_axi_gmem_ARSIZE,
	qsort_17_m_axi_gmem_ARBURST,
	qsort_17_m_axi_gmem_ARLOCK,
	qsort_17_m_axi_gmem_ARCACHE,
	qsort_17_m_axi_gmem_ARPROT,
	qsort_17_m_axi_gmem_ARQOS,
	qsort_17_m_axi_gmem_ARREGION,
	qsort_17_m_axi_gmem_ARUSER,
	qsort_17_m_axi_gmem_RREADY,
	qsort_17_m_axi_gmem_RVALID,
	qsort_17_m_axi_gmem_RID,
	qsort_17_m_axi_gmem_RDATA,
	qsort_17_m_axi_gmem_RRESP,
	qsort_17_m_axi_gmem_RLAST,
	qsort_17_m_axi_gmem_RUSER,
	qsort_17_m_axi_gmem_AWREADY,
	qsort_17_m_axi_gmem_AWVALID,
	qsort_17_m_axi_gmem_AWID,
	qsort_17_m_axi_gmem_AWADDR,
	qsort_17_m_axi_gmem_AWLEN,
	qsort_17_m_axi_gmem_AWSIZE,
	qsort_17_m_axi_gmem_AWBURST,
	qsort_17_m_axi_gmem_AWLOCK,
	qsort_17_m_axi_gmem_AWCACHE,
	qsort_17_m_axi_gmem_AWPROT,
	qsort_17_m_axi_gmem_AWQOS,
	qsort_17_m_axi_gmem_AWREGION,
	qsort_17_m_axi_gmem_AWUSER,
	qsort_17_m_axi_gmem_WREADY,
	qsort_17_m_axi_gmem_WVALID,
	qsort_17_m_axi_gmem_WDATA,
	qsort_17_m_axi_gmem_WSTRB,
	qsort_17_m_axi_gmem_WLAST,
	qsort_17_m_axi_gmem_WUSER,
	qsort_17_m_axi_gmem_BREADY,
	qsort_17_m_axi_gmem_BVALID,
	qsort_17_m_axi_gmem_BID,
	qsort_17_m_axi_gmem_BRESP,
	qsort_17_m_axi_gmem_BUSER,
	qsort_17_s_axi_control_ARREADY,
	qsort_17_s_axi_control_ARVALID,
	qsort_17_s_axi_control_ARADDR,
	qsort_17_s_axi_control_RREADY,
	qsort_17_s_axi_control_RVALID,
	qsort_17_s_axi_control_RDATA,
	qsort_17_s_axi_control_RRESP,
	qsort_17_s_axi_control_AWREADY,
	qsort_17_s_axi_control_AWVALID,
	qsort_17_s_axi_control_AWADDR,
	qsort_17_s_axi_control_WREADY,
	qsort_17_s_axi_control_WVALID,
	qsort_17_s_axi_control_WDATA,
	qsort_17_s_axi_control_WSTRB,
	qsort_17_s_axi_control_BREADY,
	qsort_17_s_axi_control_BVALID,
	qsort_17_s_axi_control_BRESP,
	qsort_18_m_axi_gmem_ARREADY,
	qsort_18_m_axi_gmem_ARVALID,
	qsort_18_m_axi_gmem_ARID,
	qsort_18_m_axi_gmem_ARADDR,
	qsort_18_m_axi_gmem_ARLEN,
	qsort_18_m_axi_gmem_ARSIZE,
	qsort_18_m_axi_gmem_ARBURST,
	qsort_18_m_axi_gmem_ARLOCK,
	qsort_18_m_axi_gmem_ARCACHE,
	qsort_18_m_axi_gmem_ARPROT,
	qsort_18_m_axi_gmem_ARQOS,
	qsort_18_m_axi_gmem_ARREGION,
	qsort_18_m_axi_gmem_ARUSER,
	qsort_18_m_axi_gmem_RREADY,
	qsort_18_m_axi_gmem_RVALID,
	qsort_18_m_axi_gmem_RID,
	qsort_18_m_axi_gmem_RDATA,
	qsort_18_m_axi_gmem_RRESP,
	qsort_18_m_axi_gmem_RLAST,
	qsort_18_m_axi_gmem_RUSER,
	qsort_18_m_axi_gmem_AWREADY,
	qsort_18_m_axi_gmem_AWVALID,
	qsort_18_m_axi_gmem_AWID,
	qsort_18_m_axi_gmem_AWADDR,
	qsort_18_m_axi_gmem_AWLEN,
	qsort_18_m_axi_gmem_AWSIZE,
	qsort_18_m_axi_gmem_AWBURST,
	qsort_18_m_axi_gmem_AWLOCK,
	qsort_18_m_axi_gmem_AWCACHE,
	qsort_18_m_axi_gmem_AWPROT,
	qsort_18_m_axi_gmem_AWQOS,
	qsort_18_m_axi_gmem_AWREGION,
	qsort_18_m_axi_gmem_AWUSER,
	qsort_18_m_axi_gmem_WREADY,
	qsort_18_m_axi_gmem_WVALID,
	qsort_18_m_axi_gmem_WDATA,
	qsort_18_m_axi_gmem_WSTRB,
	qsort_18_m_axi_gmem_WLAST,
	qsort_18_m_axi_gmem_WUSER,
	qsort_18_m_axi_gmem_BREADY,
	qsort_18_m_axi_gmem_BVALID,
	qsort_18_m_axi_gmem_BID,
	qsort_18_m_axi_gmem_BRESP,
	qsort_18_m_axi_gmem_BUSER,
	qsort_18_s_axi_control_ARREADY,
	qsort_18_s_axi_control_ARVALID,
	qsort_18_s_axi_control_ARADDR,
	qsort_18_s_axi_control_RREADY,
	qsort_18_s_axi_control_RVALID,
	qsort_18_s_axi_control_RDATA,
	qsort_18_s_axi_control_RRESP,
	qsort_18_s_axi_control_AWREADY,
	qsort_18_s_axi_control_AWVALID,
	qsort_18_s_axi_control_AWADDR,
	qsort_18_s_axi_control_WREADY,
	qsort_18_s_axi_control_WVALID,
	qsort_18_s_axi_control_WDATA,
	qsort_18_s_axi_control_WSTRB,
	qsort_18_s_axi_control_BREADY,
	qsort_18_s_axi_control_BVALID,
	qsort_18_s_axi_control_BRESP,
	qsort_19_m_axi_gmem_ARREADY,
	qsort_19_m_axi_gmem_ARVALID,
	qsort_19_m_axi_gmem_ARID,
	qsort_19_m_axi_gmem_ARADDR,
	qsort_19_m_axi_gmem_ARLEN,
	qsort_19_m_axi_gmem_ARSIZE,
	qsort_19_m_axi_gmem_ARBURST,
	qsort_19_m_axi_gmem_ARLOCK,
	qsort_19_m_axi_gmem_ARCACHE,
	qsort_19_m_axi_gmem_ARPROT,
	qsort_19_m_axi_gmem_ARQOS,
	qsort_19_m_axi_gmem_ARREGION,
	qsort_19_m_axi_gmem_ARUSER,
	qsort_19_m_axi_gmem_RREADY,
	qsort_19_m_axi_gmem_RVALID,
	qsort_19_m_axi_gmem_RID,
	qsort_19_m_axi_gmem_RDATA,
	qsort_19_m_axi_gmem_RRESP,
	qsort_19_m_axi_gmem_RLAST,
	qsort_19_m_axi_gmem_RUSER,
	qsort_19_m_axi_gmem_AWREADY,
	qsort_19_m_axi_gmem_AWVALID,
	qsort_19_m_axi_gmem_AWID,
	qsort_19_m_axi_gmem_AWADDR,
	qsort_19_m_axi_gmem_AWLEN,
	qsort_19_m_axi_gmem_AWSIZE,
	qsort_19_m_axi_gmem_AWBURST,
	qsort_19_m_axi_gmem_AWLOCK,
	qsort_19_m_axi_gmem_AWCACHE,
	qsort_19_m_axi_gmem_AWPROT,
	qsort_19_m_axi_gmem_AWQOS,
	qsort_19_m_axi_gmem_AWREGION,
	qsort_19_m_axi_gmem_AWUSER,
	qsort_19_m_axi_gmem_WREADY,
	qsort_19_m_axi_gmem_WVALID,
	qsort_19_m_axi_gmem_WDATA,
	qsort_19_m_axi_gmem_WSTRB,
	qsort_19_m_axi_gmem_WLAST,
	qsort_19_m_axi_gmem_WUSER,
	qsort_19_m_axi_gmem_BREADY,
	qsort_19_m_axi_gmem_BVALID,
	qsort_19_m_axi_gmem_BID,
	qsort_19_m_axi_gmem_BRESP,
	qsort_19_m_axi_gmem_BUSER,
	qsort_19_s_axi_control_ARREADY,
	qsort_19_s_axi_control_ARVALID,
	qsort_19_s_axi_control_ARADDR,
	qsort_19_s_axi_control_RREADY,
	qsort_19_s_axi_control_RVALID,
	qsort_19_s_axi_control_RDATA,
	qsort_19_s_axi_control_RRESP,
	qsort_19_s_axi_control_AWREADY,
	qsort_19_s_axi_control_AWVALID,
	qsort_19_s_axi_control_AWADDR,
	qsort_19_s_axi_control_WREADY,
	qsort_19_s_axi_control_WVALID,
	qsort_19_s_axi_control_WDATA,
	qsort_19_s_axi_control_WSTRB,
	qsort_19_s_axi_control_BREADY,
	qsort_19_s_axi_control_BVALID,
	qsort_19_s_axi_control_BRESP,
	qsort_20_m_axi_gmem_ARREADY,
	qsort_20_m_axi_gmem_ARVALID,
	qsort_20_m_axi_gmem_ARID,
	qsort_20_m_axi_gmem_ARADDR,
	qsort_20_m_axi_gmem_ARLEN,
	qsort_20_m_axi_gmem_ARSIZE,
	qsort_20_m_axi_gmem_ARBURST,
	qsort_20_m_axi_gmem_ARLOCK,
	qsort_20_m_axi_gmem_ARCACHE,
	qsort_20_m_axi_gmem_ARPROT,
	qsort_20_m_axi_gmem_ARQOS,
	qsort_20_m_axi_gmem_ARREGION,
	qsort_20_m_axi_gmem_ARUSER,
	qsort_20_m_axi_gmem_RREADY,
	qsort_20_m_axi_gmem_RVALID,
	qsort_20_m_axi_gmem_RID,
	qsort_20_m_axi_gmem_RDATA,
	qsort_20_m_axi_gmem_RRESP,
	qsort_20_m_axi_gmem_RLAST,
	qsort_20_m_axi_gmem_RUSER,
	qsort_20_m_axi_gmem_AWREADY,
	qsort_20_m_axi_gmem_AWVALID,
	qsort_20_m_axi_gmem_AWID,
	qsort_20_m_axi_gmem_AWADDR,
	qsort_20_m_axi_gmem_AWLEN,
	qsort_20_m_axi_gmem_AWSIZE,
	qsort_20_m_axi_gmem_AWBURST,
	qsort_20_m_axi_gmem_AWLOCK,
	qsort_20_m_axi_gmem_AWCACHE,
	qsort_20_m_axi_gmem_AWPROT,
	qsort_20_m_axi_gmem_AWQOS,
	qsort_20_m_axi_gmem_AWREGION,
	qsort_20_m_axi_gmem_AWUSER,
	qsort_20_m_axi_gmem_WREADY,
	qsort_20_m_axi_gmem_WVALID,
	qsort_20_m_axi_gmem_WDATA,
	qsort_20_m_axi_gmem_WSTRB,
	qsort_20_m_axi_gmem_WLAST,
	qsort_20_m_axi_gmem_WUSER,
	qsort_20_m_axi_gmem_BREADY,
	qsort_20_m_axi_gmem_BVALID,
	qsort_20_m_axi_gmem_BID,
	qsort_20_m_axi_gmem_BRESP,
	qsort_20_m_axi_gmem_BUSER,
	qsort_20_s_axi_control_ARREADY,
	qsort_20_s_axi_control_ARVALID,
	qsort_20_s_axi_control_ARADDR,
	qsort_20_s_axi_control_RREADY,
	qsort_20_s_axi_control_RVALID,
	qsort_20_s_axi_control_RDATA,
	qsort_20_s_axi_control_RRESP,
	qsort_20_s_axi_control_AWREADY,
	qsort_20_s_axi_control_AWVALID,
	qsort_20_s_axi_control_AWADDR,
	qsort_20_s_axi_control_WREADY,
	qsort_20_s_axi_control_WVALID,
	qsort_20_s_axi_control_WDATA,
	qsort_20_s_axi_control_WSTRB,
	qsort_20_s_axi_control_BREADY,
	qsort_20_s_axi_control_BVALID,
	qsort_20_s_axi_control_BRESP,
	qsort_21_m_axi_gmem_ARREADY,
	qsort_21_m_axi_gmem_ARVALID,
	qsort_21_m_axi_gmem_ARID,
	qsort_21_m_axi_gmem_ARADDR,
	qsort_21_m_axi_gmem_ARLEN,
	qsort_21_m_axi_gmem_ARSIZE,
	qsort_21_m_axi_gmem_ARBURST,
	qsort_21_m_axi_gmem_ARLOCK,
	qsort_21_m_axi_gmem_ARCACHE,
	qsort_21_m_axi_gmem_ARPROT,
	qsort_21_m_axi_gmem_ARQOS,
	qsort_21_m_axi_gmem_ARREGION,
	qsort_21_m_axi_gmem_ARUSER,
	qsort_21_m_axi_gmem_RREADY,
	qsort_21_m_axi_gmem_RVALID,
	qsort_21_m_axi_gmem_RID,
	qsort_21_m_axi_gmem_RDATA,
	qsort_21_m_axi_gmem_RRESP,
	qsort_21_m_axi_gmem_RLAST,
	qsort_21_m_axi_gmem_RUSER,
	qsort_21_m_axi_gmem_AWREADY,
	qsort_21_m_axi_gmem_AWVALID,
	qsort_21_m_axi_gmem_AWID,
	qsort_21_m_axi_gmem_AWADDR,
	qsort_21_m_axi_gmem_AWLEN,
	qsort_21_m_axi_gmem_AWSIZE,
	qsort_21_m_axi_gmem_AWBURST,
	qsort_21_m_axi_gmem_AWLOCK,
	qsort_21_m_axi_gmem_AWCACHE,
	qsort_21_m_axi_gmem_AWPROT,
	qsort_21_m_axi_gmem_AWQOS,
	qsort_21_m_axi_gmem_AWREGION,
	qsort_21_m_axi_gmem_AWUSER,
	qsort_21_m_axi_gmem_WREADY,
	qsort_21_m_axi_gmem_WVALID,
	qsort_21_m_axi_gmem_WDATA,
	qsort_21_m_axi_gmem_WSTRB,
	qsort_21_m_axi_gmem_WLAST,
	qsort_21_m_axi_gmem_WUSER,
	qsort_21_m_axi_gmem_BREADY,
	qsort_21_m_axi_gmem_BVALID,
	qsort_21_m_axi_gmem_BID,
	qsort_21_m_axi_gmem_BRESP,
	qsort_21_m_axi_gmem_BUSER,
	qsort_21_s_axi_control_ARREADY,
	qsort_21_s_axi_control_ARVALID,
	qsort_21_s_axi_control_ARADDR,
	qsort_21_s_axi_control_RREADY,
	qsort_21_s_axi_control_RVALID,
	qsort_21_s_axi_control_RDATA,
	qsort_21_s_axi_control_RRESP,
	qsort_21_s_axi_control_AWREADY,
	qsort_21_s_axi_control_AWVALID,
	qsort_21_s_axi_control_AWADDR,
	qsort_21_s_axi_control_WREADY,
	qsort_21_s_axi_control_WVALID,
	qsort_21_s_axi_control_WDATA,
	qsort_21_s_axi_control_WSTRB,
	qsort_21_s_axi_control_BREADY,
	qsort_21_s_axi_control_BVALID,
	qsort_21_s_axi_control_BRESP,
	qsort_22_m_axi_gmem_ARREADY,
	qsort_22_m_axi_gmem_ARVALID,
	qsort_22_m_axi_gmem_ARID,
	qsort_22_m_axi_gmem_ARADDR,
	qsort_22_m_axi_gmem_ARLEN,
	qsort_22_m_axi_gmem_ARSIZE,
	qsort_22_m_axi_gmem_ARBURST,
	qsort_22_m_axi_gmem_ARLOCK,
	qsort_22_m_axi_gmem_ARCACHE,
	qsort_22_m_axi_gmem_ARPROT,
	qsort_22_m_axi_gmem_ARQOS,
	qsort_22_m_axi_gmem_ARREGION,
	qsort_22_m_axi_gmem_ARUSER,
	qsort_22_m_axi_gmem_RREADY,
	qsort_22_m_axi_gmem_RVALID,
	qsort_22_m_axi_gmem_RID,
	qsort_22_m_axi_gmem_RDATA,
	qsort_22_m_axi_gmem_RRESP,
	qsort_22_m_axi_gmem_RLAST,
	qsort_22_m_axi_gmem_RUSER,
	qsort_22_m_axi_gmem_AWREADY,
	qsort_22_m_axi_gmem_AWVALID,
	qsort_22_m_axi_gmem_AWID,
	qsort_22_m_axi_gmem_AWADDR,
	qsort_22_m_axi_gmem_AWLEN,
	qsort_22_m_axi_gmem_AWSIZE,
	qsort_22_m_axi_gmem_AWBURST,
	qsort_22_m_axi_gmem_AWLOCK,
	qsort_22_m_axi_gmem_AWCACHE,
	qsort_22_m_axi_gmem_AWPROT,
	qsort_22_m_axi_gmem_AWQOS,
	qsort_22_m_axi_gmem_AWREGION,
	qsort_22_m_axi_gmem_AWUSER,
	qsort_22_m_axi_gmem_WREADY,
	qsort_22_m_axi_gmem_WVALID,
	qsort_22_m_axi_gmem_WDATA,
	qsort_22_m_axi_gmem_WSTRB,
	qsort_22_m_axi_gmem_WLAST,
	qsort_22_m_axi_gmem_WUSER,
	qsort_22_m_axi_gmem_BREADY,
	qsort_22_m_axi_gmem_BVALID,
	qsort_22_m_axi_gmem_BID,
	qsort_22_m_axi_gmem_BRESP,
	qsort_22_m_axi_gmem_BUSER,
	qsort_22_s_axi_control_ARREADY,
	qsort_22_s_axi_control_ARVALID,
	qsort_22_s_axi_control_ARADDR,
	qsort_22_s_axi_control_RREADY,
	qsort_22_s_axi_control_RVALID,
	qsort_22_s_axi_control_RDATA,
	qsort_22_s_axi_control_RRESP,
	qsort_22_s_axi_control_AWREADY,
	qsort_22_s_axi_control_AWVALID,
	qsort_22_s_axi_control_AWADDR,
	qsort_22_s_axi_control_WREADY,
	qsort_22_s_axi_control_WVALID,
	qsort_22_s_axi_control_WDATA,
	qsort_22_s_axi_control_WSTRB,
	qsort_22_s_axi_control_BREADY,
	qsort_22_s_axi_control_BVALID,
	qsort_22_s_axi_control_BRESP,
	qsort_23_m_axi_gmem_ARREADY,
	qsort_23_m_axi_gmem_ARVALID,
	qsort_23_m_axi_gmem_ARID,
	qsort_23_m_axi_gmem_ARADDR,
	qsort_23_m_axi_gmem_ARLEN,
	qsort_23_m_axi_gmem_ARSIZE,
	qsort_23_m_axi_gmem_ARBURST,
	qsort_23_m_axi_gmem_ARLOCK,
	qsort_23_m_axi_gmem_ARCACHE,
	qsort_23_m_axi_gmem_ARPROT,
	qsort_23_m_axi_gmem_ARQOS,
	qsort_23_m_axi_gmem_ARREGION,
	qsort_23_m_axi_gmem_ARUSER,
	qsort_23_m_axi_gmem_RREADY,
	qsort_23_m_axi_gmem_RVALID,
	qsort_23_m_axi_gmem_RID,
	qsort_23_m_axi_gmem_RDATA,
	qsort_23_m_axi_gmem_RRESP,
	qsort_23_m_axi_gmem_RLAST,
	qsort_23_m_axi_gmem_RUSER,
	qsort_23_m_axi_gmem_AWREADY,
	qsort_23_m_axi_gmem_AWVALID,
	qsort_23_m_axi_gmem_AWID,
	qsort_23_m_axi_gmem_AWADDR,
	qsort_23_m_axi_gmem_AWLEN,
	qsort_23_m_axi_gmem_AWSIZE,
	qsort_23_m_axi_gmem_AWBURST,
	qsort_23_m_axi_gmem_AWLOCK,
	qsort_23_m_axi_gmem_AWCACHE,
	qsort_23_m_axi_gmem_AWPROT,
	qsort_23_m_axi_gmem_AWQOS,
	qsort_23_m_axi_gmem_AWREGION,
	qsort_23_m_axi_gmem_AWUSER,
	qsort_23_m_axi_gmem_WREADY,
	qsort_23_m_axi_gmem_WVALID,
	qsort_23_m_axi_gmem_WDATA,
	qsort_23_m_axi_gmem_WSTRB,
	qsort_23_m_axi_gmem_WLAST,
	qsort_23_m_axi_gmem_WUSER,
	qsort_23_m_axi_gmem_BREADY,
	qsort_23_m_axi_gmem_BVALID,
	qsort_23_m_axi_gmem_BID,
	qsort_23_m_axi_gmem_BRESP,
	qsort_23_m_axi_gmem_BUSER,
	qsort_23_s_axi_control_ARREADY,
	qsort_23_s_axi_control_ARVALID,
	qsort_23_s_axi_control_ARADDR,
	qsort_23_s_axi_control_RREADY,
	qsort_23_s_axi_control_RVALID,
	qsort_23_s_axi_control_RDATA,
	qsort_23_s_axi_control_RRESP,
	qsort_23_s_axi_control_AWREADY,
	qsort_23_s_axi_control_AWVALID,
	qsort_23_s_axi_control_AWADDR,
	qsort_23_s_axi_control_WREADY,
	qsort_23_s_axi_control_WVALID,
	qsort_23_s_axi_control_WDATA,
	qsort_23_s_axi_control_WSTRB,
	qsort_23_s_axi_control_BREADY,
	qsort_23_s_axi_control_BVALID,
	qsort_23_s_axi_control_BRESP,
	qsort_24_m_axi_gmem_ARREADY,
	qsort_24_m_axi_gmem_ARVALID,
	qsort_24_m_axi_gmem_ARID,
	qsort_24_m_axi_gmem_ARADDR,
	qsort_24_m_axi_gmem_ARLEN,
	qsort_24_m_axi_gmem_ARSIZE,
	qsort_24_m_axi_gmem_ARBURST,
	qsort_24_m_axi_gmem_ARLOCK,
	qsort_24_m_axi_gmem_ARCACHE,
	qsort_24_m_axi_gmem_ARPROT,
	qsort_24_m_axi_gmem_ARQOS,
	qsort_24_m_axi_gmem_ARREGION,
	qsort_24_m_axi_gmem_ARUSER,
	qsort_24_m_axi_gmem_RREADY,
	qsort_24_m_axi_gmem_RVALID,
	qsort_24_m_axi_gmem_RID,
	qsort_24_m_axi_gmem_RDATA,
	qsort_24_m_axi_gmem_RRESP,
	qsort_24_m_axi_gmem_RLAST,
	qsort_24_m_axi_gmem_RUSER,
	qsort_24_m_axi_gmem_AWREADY,
	qsort_24_m_axi_gmem_AWVALID,
	qsort_24_m_axi_gmem_AWID,
	qsort_24_m_axi_gmem_AWADDR,
	qsort_24_m_axi_gmem_AWLEN,
	qsort_24_m_axi_gmem_AWSIZE,
	qsort_24_m_axi_gmem_AWBURST,
	qsort_24_m_axi_gmem_AWLOCK,
	qsort_24_m_axi_gmem_AWCACHE,
	qsort_24_m_axi_gmem_AWPROT,
	qsort_24_m_axi_gmem_AWQOS,
	qsort_24_m_axi_gmem_AWREGION,
	qsort_24_m_axi_gmem_AWUSER,
	qsort_24_m_axi_gmem_WREADY,
	qsort_24_m_axi_gmem_WVALID,
	qsort_24_m_axi_gmem_WDATA,
	qsort_24_m_axi_gmem_WSTRB,
	qsort_24_m_axi_gmem_WLAST,
	qsort_24_m_axi_gmem_WUSER,
	qsort_24_m_axi_gmem_BREADY,
	qsort_24_m_axi_gmem_BVALID,
	qsort_24_m_axi_gmem_BID,
	qsort_24_m_axi_gmem_BRESP,
	qsort_24_m_axi_gmem_BUSER,
	qsort_24_s_axi_control_ARREADY,
	qsort_24_s_axi_control_ARVALID,
	qsort_24_s_axi_control_ARADDR,
	qsort_24_s_axi_control_RREADY,
	qsort_24_s_axi_control_RVALID,
	qsort_24_s_axi_control_RDATA,
	qsort_24_s_axi_control_RRESP,
	qsort_24_s_axi_control_AWREADY,
	qsort_24_s_axi_control_AWVALID,
	qsort_24_s_axi_control_AWADDR,
	qsort_24_s_axi_control_WREADY,
	qsort_24_s_axi_control_WVALID,
	qsort_24_s_axi_control_WDATA,
	qsort_24_s_axi_control_WSTRB,
	qsort_24_s_axi_control_BREADY,
	qsort_24_s_axi_control_BVALID,
	qsort_24_s_axi_control_BRESP,
	qsort_25_m_axi_gmem_ARREADY,
	qsort_25_m_axi_gmem_ARVALID,
	qsort_25_m_axi_gmem_ARID,
	qsort_25_m_axi_gmem_ARADDR,
	qsort_25_m_axi_gmem_ARLEN,
	qsort_25_m_axi_gmem_ARSIZE,
	qsort_25_m_axi_gmem_ARBURST,
	qsort_25_m_axi_gmem_ARLOCK,
	qsort_25_m_axi_gmem_ARCACHE,
	qsort_25_m_axi_gmem_ARPROT,
	qsort_25_m_axi_gmem_ARQOS,
	qsort_25_m_axi_gmem_ARREGION,
	qsort_25_m_axi_gmem_ARUSER,
	qsort_25_m_axi_gmem_RREADY,
	qsort_25_m_axi_gmem_RVALID,
	qsort_25_m_axi_gmem_RID,
	qsort_25_m_axi_gmem_RDATA,
	qsort_25_m_axi_gmem_RRESP,
	qsort_25_m_axi_gmem_RLAST,
	qsort_25_m_axi_gmem_RUSER,
	qsort_25_m_axi_gmem_AWREADY,
	qsort_25_m_axi_gmem_AWVALID,
	qsort_25_m_axi_gmem_AWID,
	qsort_25_m_axi_gmem_AWADDR,
	qsort_25_m_axi_gmem_AWLEN,
	qsort_25_m_axi_gmem_AWSIZE,
	qsort_25_m_axi_gmem_AWBURST,
	qsort_25_m_axi_gmem_AWLOCK,
	qsort_25_m_axi_gmem_AWCACHE,
	qsort_25_m_axi_gmem_AWPROT,
	qsort_25_m_axi_gmem_AWQOS,
	qsort_25_m_axi_gmem_AWREGION,
	qsort_25_m_axi_gmem_AWUSER,
	qsort_25_m_axi_gmem_WREADY,
	qsort_25_m_axi_gmem_WVALID,
	qsort_25_m_axi_gmem_WDATA,
	qsort_25_m_axi_gmem_WSTRB,
	qsort_25_m_axi_gmem_WLAST,
	qsort_25_m_axi_gmem_WUSER,
	qsort_25_m_axi_gmem_BREADY,
	qsort_25_m_axi_gmem_BVALID,
	qsort_25_m_axi_gmem_BID,
	qsort_25_m_axi_gmem_BRESP,
	qsort_25_m_axi_gmem_BUSER,
	qsort_25_s_axi_control_ARREADY,
	qsort_25_s_axi_control_ARVALID,
	qsort_25_s_axi_control_ARADDR,
	qsort_25_s_axi_control_RREADY,
	qsort_25_s_axi_control_RVALID,
	qsort_25_s_axi_control_RDATA,
	qsort_25_s_axi_control_RRESP,
	qsort_25_s_axi_control_AWREADY,
	qsort_25_s_axi_control_AWVALID,
	qsort_25_s_axi_control_AWADDR,
	qsort_25_s_axi_control_WREADY,
	qsort_25_s_axi_control_WVALID,
	qsort_25_s_axi_control_WDATA,
	qsort_25_s_axi_control_WSTRB,
	qsort_25_s_axi_control_BREADY,
	qsort_25_s_axi_control_BVALID,
	qsort_25_s_axi_control_BRESP,
	qsort_26_m_axi_gmem_ARREADY,
	qsort_26_m_axi_gmem_ARVALID,
	qsort_26_m_axi_gmem_ARID,
	qsort_26_m_axi_gmem_ARADDR,
	qsort_26_m_axi_gmem_ARLEN,
	qsort_26_m_axi_gmem_ARSIZE,
	qsort_26_m_axi_gmem_ARBURST,
	qsort_26_m_axi_gmem_ARLOCK,
	qsort_26_m_axi_gmem_ARCACHE,
	qsort_26_m_axi_gmem_ARPROT,
	qsort_26_m_axi_gmem_ARQOS,
	qsort_26_m_axi_gmem_ARREGION,
	qsort_26_m_axi_gmem_ARUSER,
	qsort_26_m_axi_gmem_RREADY,
	qsort_26_m_axi_gmem_RVALID,
	qsort_26_m_axi_gmem_RID,
	qsort_26_m_axi_gmem_RDATA,
	qsort_26_m_axi_gmem_RRESP,
	qsort_26_m_axi_gmem_RLAST,
	qsort_26_m_axi_gmem_RUSER,
	qsort_26_m_axi_gmem_AWREADY,
	qsort_26_m_axi_gmem_AWVALID,
	qsort_26_m_axi_gmem_AWID,
	qsort_26_m_axi_gmem_AWADDR,
	qsort_26_m_axi_gmem_AWLEN,
	qsort_26_m_axi_gmem_AWSIZE,
	qsort_26_m_axi_gmem_AWBURST,
	qsort_26_m_axi_gmem_AWLOCK,
	qsort_26_m_axi_gmem_AWCACHE,
	qsort_26_m_axi_gmem_AWPROT,
	qsort_26_m_axi_gmem_AWQOS,
	qsort_26_m_axi_gmem_AWREGION,
	qsort_26_m_axi_gmem_AWUSER,
	qsort_26_m_axi_gmem_WREADY,
	qsort_26_m_axi_gmem_WVALID,
	qsort_26_m_axi_gmem_WDATA,
	qsort_26_m_axi_gmem_WSTRB,
	qsort_26_m_axi_gmem_WLAST,
	qsort_26_m_axi_gmem_WUSER,
	qsort_26_m_axi_gmem_BREADY,
	qsort_26_m_axi_gmem_BVALID,
	qsort_26_m_axi_gmem_BID,
	qsort_26_m_axi_gmem_BRESP,
	qsort_26_m_axi_gmem_BUSER,
	qsort_26_s_axi_control_ARREADY,
	qsort_26_s_axi_control_ARVALID,
	qsort_26_s_axi_control_ARADDR,
	qsort_26_s_axi_control_RREADY,
	qsort_26_s_axi_control_RVALID,
	qsort_26_s_axi_control_RDATA,
	qsort_26_s_axi_control_RRESP,
	qsort_26_s_axi_control_AWREADY,
	qsort_26_s_axi_control_AWVALID,
	qsort_26_s_axi_control_AWADDR,
	qsort_26_s_axi_control_WREADY,
	qsort_26_s_axi_control_WVALID,
	qsort_26_s_axi_control_WDATA,
	qsort_26_s_axi_control_WSTRB,
	qsort_26_s_axi_control_BREADY,
	qsort_26_s_axi_control_BVALID,
	qsort_26_s_axi_control_BRESP,
	qsort_27_m_axi_gmem_ARREADY,
	qsort_27_m_axi_gmem_ARVALID,
	qsort_27_m_axi_gmem_ARID,
	qsort_27_m_axi_gmem_ARADDR,
	qsort_27_m_axi_gmem_ARLEN,
	qsort_27_m_axi_gmem_ARSIZE,
	qsort_27_m_axi_gmem_ARBURST,
	qsort_27_m_axi_gmem_ARLOCK,
	qsort_27_m_axi_gmem_ARCACHE,
	qsort_27_m_axi_gmem_ARPROT,
	qsort_27_m_axi_gmem_ARQOS,
	qsort_27_m_axi_gmem_ARREGION,
	qsort_27_m_axi_gmem_ARUSER,
	qsort_27_m_axi_gmem_RREADY,
	qsort_27_m_axi_gmem_RVALID,
	qsort_27_m_axi_gmem_RID,
	qsort_27_m_axi_gmem_RDATA,
	qsort_27_m_axi_gmem_RRESP,
	qsort_27_m_axi_gmem_RLAST,
	qsort_27_m_axi_gmem_RUSER,
	qsort_27_m_axi_gmem_AWREADY,
	qsort_27_m_axi_gmem_AWVALID,
	qsort_27_m_axi_gmem_AWID,
	qsort_27_m_axi_gmem_AWADDR,
	qsort_27_m_axi_gmem_AWLEN,
	qsort_27_m_axi_gmem_AWSIZE,
	qsort_27_m_axi_gmem_AWBURST,
	qsort_27_m_axi_gmem_AWLOCK,
	qsort_27_m_axi_gmem_AWCACHE,
	qsort_27_m_axi_gmem_AWPROT,
	qsort_27_m_axi_gmem_AWQOS,
	qsort_27_m_axi_gmem_AWREGION,
	qsort_27_m_axi_gmem_AWUSER,
	qsort_27_m_axi_gmem_WREADY,
	qsort_27_m_axi_gmem_WVALID,
	qsort_27_m_axi_gmem_WDATA,
	qsort_27_m_axi_gmem_WSTRB,
	qsort_27_m_axi_gmem_WLAST,
	qsort_27_m_axi_gmem_WUSER,
	qsort_27_m_axi_gmem_BREADY,
	qsort_27_m_axi_gmem_BVALID,
	qsort_27_m_axi_gmem_BID,
	qsort_27_m_axi_gmem_BRESP,
	qsort_27_m_axi_gmem_BUSER,
	qsort_27_s_axi_control_ARREADY,
	qsort_27_s_axi_control_ARVALID,
	qsort_27_s_axi_control_ARADDR,
	qsort_27_s_axi_control_RREADY,
	qsort_27_s_axi_control_RVALID,
	qsort_27_s_axi_control_RDATA,
	qsort_27_s_axi_control_RRESP,
	qsort_27_s_axi_control_AWREADY,
	qsort_27_s_axi_control_AWVALID,
	qsort_27_s_axi_control_AWADDR,
	qsort_27_s_axi_control_WREADY,
	qsort_27_s_axi_control_WVALID,
	qsort_27_s_axi_control_WDATA,
	qsort_27_s_axi_control_WSTRB,
	qsort_27_s_axi_control_BREADY,
	qsort_27_s_axi_control_BVALID,
	qsort_27_s_axi_control_BRESP,
	qsort_28_m_axi_gmem_ARREADY,
	qsort_28_m_axi_gmem_ARVALID,
	qsort_28_m_axi_gmem_ARID,
	qsort_28_m_axi_gmem_ARADDR,
	qsort_28_m_axi_gmem_ARLEN,
	qsort_28_m_axi_gmem_ARSIZE,
	qsort_28_m_axi_gmem_ARBURST,
	qsort_28_m_axi_gmem_ARLOCK,
	qsort_28_m_axi_gmem_ARCACHE,
	qsort_28_m_axi_gmem_ARPROT,
	qsort_28_m_axi_gmem_ARQOS,
	qsort_28_m_axi_gmem_ARREGION,
	qsort_28_m_axi_gmem_ARUSER,
	qsort_28_m_axi_gmem_RREADY,
	qsort_28_m_axi_gmem_RVALID,
	qsort_28_m_axi_gmem_RID,
	qsort_28_m_axi_gmem_RDATA,
	qsort_28_m_axi_gmem_RRESP,
	qsort_28_m_axi_gmem_RLAST,
	qsort_28_m_axi_gmem_RUSER,
	qsort_28_m_axi_gmem_AWREADY,
	qsort_28_m_axi_gmem_AWVALID,
	qsort_28_m_axi_gmem_AWID,
	qsort_28_m_axi_gmem_AWADDR,
	qsort_28_m_axi_gmem_AWLEN,
	qsort_28_m_axi_gmem_AWSIZE,
	qsort_28_m_axi_gmem_AWBURST,
	qsort_28_m_axi_gmem_AWLOCK,
	qsort_28_m_axi_gmem_AWCACHE,
	qsort_28_m_axi_gmem_AWPROT,
	qsort_28_m_axi_gmem_AWQOS,
	qsort_28_m_axi_gmem_AWREGION,
	qsort_28_m_axi_gmem_AWUSER,
	qsort_28_m_axi_gmem_WREADY,
	qsort_28_m_axi_gmem_WVALID,
	qsort_28_m_axi_gmem_WDATA,
	qsort_28_m_axi_gmem_WSTRB,
	qsort_28_m_axi_gmem_WLAST,
	qsort_28_m_axi_gmem_WUSER,
	qsort_28_m_axi_gmem_BREADY,
	qsort_28_m_axi_gmem_BVALID,
	qsort_28_m_axi_gmem_BID,
	qsort_28_m_axi_gmem_BRESP,
	qsort_28_m_axi_gmem_BUSER,
	qsort_28_s_axi_control_ARREADY,
	qsort_28_s_axi_control_ARVALID,
	qsort_28_s_axi_control_ARADDR,
	qsort_28_s_axi_control_RREADY,
	qsort_28_s_axi_control_RVALID,
	qsort_28_s_axi_control_RDATA,
	qsort_28_s_axi_control_RRESP,
	qsort_28_s_axi_control_AWREADY,
	qsort_28_s_axi_control_AWVALID,
	qsort_28_s_axi_control_AWADDR,
	qsort_28_s_axi_control_WREADY,
	qsort_28_s_axi_control_WVALID,
	qsort_28_s_axi_control_WDATA,
	qsort_28_s_axi_control_WSTRB,
	qsort_28_s_axi_control_BREADY,
	qsort_28_s_axi_control_BVALID,
	qsort_28_s_axi_control_BRESP,
	qsort_29_m_axi_gmem_ARREADY,
	qsort_29_m_axi_gmem_ARVALID,
	qsort_29_m_axi_gmem_ARID,
	qsort_29_m_axi_gmem_ARADDR,
	qsort_29_m_axi_gmem_ARLEN,
	qsort_29_m_axi_gmem_ARSIZE,
	qsort_29_m_axi_gmem_ARBURST,
	qsort_29_m_axi_gmem_ARLOCK,
	qsort_29_m_axi_gmem_ARCACHE,
	qsort_29_m_axi_gmem_ARPROT,
	qsort_29_m_axi_gmem_ARQOS,
	qsort_29_m_axi_gmem_ARREGION,
	qsort_29_m_axi_gmem_ARUSER,
	qsort_29_m_axi_gmem_RREADY,
	qsort_29_m_axi_gmem_RVALID,
	qsort_29_m_axi_gmem_RID,
	qsort_29_m_axi_gmem_RDATA,
	qsort_29_m_axi_gmem_RRESP,
	qsort_29_m_axi_gmem_RLAST,
	qsort_29_m_axi_gmem_RUSER,
	qsort_29_m_axi_gmem_AWREADY,
	qsort_29_m_axi_gmem_AWVALID,
	qsort_29_m_axi_gmem_AWID,
	qsort_29_m_axi_gmem_AWADDR,
	qsort_29_m_axi_gmem_AWLEN,
	qsort_29_m_axi_gmem_AWSIZE,
	qsort_29_m_axi_gmem_AWBURST,
	qsort_29_m_axi_gmem_AWLOCK,
	qsort_29_m_axi_gmem_AWCACHE,
	qsort_29_m_axi_gmem_AWPROT,
	qsort_29_m_axi_gmem_AWQOS,
	qsort_29_m_axi_gmem_AWREGION,
	qsort_29_m_axi_gmem_AWUSER,
	qsort_29_m_axi_gmem_WREADY,
	qsort_29_m_axi_gmem_WVALID,
	qsort_29_m_axi_gmem_WDATA,
	qsort_29_m_axi_gmem_WSTRB,
	qsort_29_m_axi_gmem_WLAST,
	qsort_29_m_axi_gmem_WUSER,
	qsort_29_m_axi_gmem_BREADY,
	qsort_29_m_axi_gmem_BVALID,
	qsort_29_m_axi_gmem_BID,
	qsort_29_m_axi_gmem_BRESP,
	qsort_29_m_axi_gmem_BUSER,
	qsort_29_s_axi_control_ARREADY,
	qsort_29_s_axi_control_ARVALID,
	qsort_29_s_axi_control_ARADDR,
	qsort_29_s_axi_control_RREADY,
	qsort_29_s_axi_control_RVALID,
	qsort_29_s_axi_control_RDATA,
	qsort_29_s_axi_control_RRESP,
	qsort_29_s_axi_control_AWREADY,
	qsort_29_s_axi_control_AWVALID,
	qsort_29_s_axi_control_AWADDR,
	qsort_29_s_axi_control_WREADY,
	qsort_29_s_axi_control_WVALID,
	qsort_29_s_axi_control_WDATA,
	qsort_29_s_axi_control_WSTRB,
	qsort_29_s_axi_control_BREADY,
	qsort_29_s_axi_control_BVALID,
	qsort_29_s_axi_control_BRESP,
	qsort_30_m_axi_gmem_ARREADY,
	qsort_30_m_axi_gmem_ARVALID,
	qsort_30_m_axi_gmem_ARID,
	qsort_30_m_axi_gmem_ARADDR,
	qsort_30_m_axi_gmem_ARLEN,
	qsort_30_m_axi_gmem_ARSIZE,
	qsort_30_m_axi_gmem_ARBURST,
	qsort_30_m_axi_gmem_ARLOCK,
	qsort_30_m_axi_gmem_ARCACHE,
	qsort_30_m_axi_gmem_ARPROT,
	qsort_30_m_axi_gmem_ARQOS,
	qsort_30_m_axi_gmem_ARREGION,
	qsort_30_m_axi_gmem_ARUSER,
	qsort_30_m_axi_gmem_RREADY,
	qsort_30_m_axi_gmem_RVALID,
	qsort_30_m_axi_gmem_RID,
	qsort_30_m_axi_gmem_RDATA,
	qsort_30_m_axi_gmem_RRESP,
	qsort_30_m_axi_gmem_RLAST,
	qsort_30_m_axi_gmem_RUSER,
	qsort_30_m_axi_gmem_AWREADY,
	qsort_30_m_axi_gmem_AWVALID,
	qsort_30_m_axi_gmem_AWID,
	qsort_30_m_axi_gmem_AWADDR,
	qsort_30_m_axi_gmem_AWLEN,
	qsort_30_m_axi_gmem_AWSIZE,
	qsort_30_m_axi_gmem_AWBURST,
	qsort_30_m_axi_gmem_AWLOCK,
	qsort_30_m_axi_gmem_AWCACHE,
	qsort_30_m_axi_gmem_AWPROT,
	qsort_30_m_axi_gmem_AWQOS,
	qsort_30_m_axi_gmem_AWREGION,
	qsort_30_m_axi_gmem_AWUSER,
	qsort_30_m_axi_gmem_WREADY,
	qsort_30_m_axi_gmem_WVALID,
	qsort_30_m_axi_gmem_WDATA,
	qsort_30_m_axi_gmem_WSTRB,
	qsort_30_m_axi_gmem_WLAST,
	qsort_30_m_axi_gmem_WUSER,
	qsort_30_m_axi_gmem_BREADY,
	qsort_30_m_axi_gmem_BVALID,
	qsort_30_m_axi_gmem_BID,
	qsort_30_m_axi_gmem_BRESP,
	qsort_30_m_axi_gmem_BUSER,
	qsort_30_s_axi_control_ARREADY,
	qsort_30_s_axi_control_ARVALID,
	qsort_30_s_axi_control_ARADDR,
	qsort_30_s_axi_control_RREADY,
	qsort_30_s_axi_control_RVALID,
	qsort_30_s_axi_control_RDATA,
	qsort_30_s_axi_control_RRESP,
	qsort_30_s_axi_control_AWREADY,
	qsort_30_s_axi_control_AWVALID,
	qsort_30_s_axi_control_AWADDR,
	qsort_30_s_axi_control_WREADY,
	qsort_30_s_axi_control_WVALID,
	qsort_30_s_axi_control_WDATA,
	qsort_30_s_axi_control_WSTRB,
	qsort_30_s_axi_control_BREADY,
	qsort_30_s_axi_control_BVALID,
	qsort_30_s_axi_control_BRESP,
	qsort_31_m_axi_gmem_ARREADY,
	qsort_31_m_axi_gmem_ARVALID,
	qsort_31_m_axi_gmem_ARID,
	qsort_31_m_axi_gmem_ARADDR,
	qsort_31_m_axi_gmem_ARLEN,
	qsort_31_m_axi_gmem_ARSIZE,
	qsort_31_m_axi_gmem_ARBURST,
	qsort_31_m_axi_gmem_ARLOCK,
	qsort_31_m_axi_gmem_ARCACHE,
	qsort_31_m_axi_gmem_ARPROT,
	qsort_31_m_axi_gmem_ARQOS,
	qsort_31_m_axi_gmem_ARREGION,
	qsort_31_m_axi_gmem_ARUSER,
	qsort_31_m_axi_gmem_RREADY,
	qsort_31_m_axi_gmem_RVALID,
	qsort_31_m_axi_gmem_RID,
	qsort_31_m_axi_gmem_RDATA,
	qsort_31_m_axi_gmem_RRESP,
	qsort_31_m_axi_gmem_RLAST,
	qsort_31_m_axi_gmem_RUSER,
	qsort_31_m_axi_gmem_AWREADY,
	qsort_31_m_axi_gmem_AWVALID,
	qsort_31_m_axi_gmem_AWID,
	qsort_31_m_axi_gmem_AWADDR,
	qsort_31_m_axi_gmem_AWLEN,
	qsort_31_m_axi_gmem_AWSIZE,
	qsort_31_m_axi_gmem_AWBURST,
	qsort_31_m_axi_gmem_AWLOCK,
	qsort_31_m_axi_gmem_AWCACHE,
	qsort_31_m_axi_gmem_AWPROT,
	qsort_31_m_axi_gmem_AWQOS,
	qsort_31_m_axi_gmem_AWREGION,
	qsort_31_m_axi_gmem_AWUSER,
	qsort_31_m_axi_gmem_WREADY,
	qsort_31_m_axi_gmem_WVALID,
	qsort_31_m_axi_gmem_WDATA,
	qsort_31_m_axi_gmem_WSTRB,
	qsort_31_m_axi_gmem_WLAST,
	qsort_31_m_axi_gmem_WUSER,
	qsort_31_m_axi_gmem_BREADY,
	qsort_31_m_axi_gmem_BVALID,
	qsort_31_m_axi_gmem_BID,
	qsort_31_m_axi_gmem_BRESP,
	qsort_31_m_axi_gmem_BUSER,
	qsort_31_s_axi_control_ARREADY,
	qsort_31_s_axi_control_ARVALID,
	qsort_31_s_axi_control_ARADDR,
	qsort_31_s_axi_control_RREADY,
	qsort_31_s_axi_control_RVALID,
	qsort_31_s_axi_control_RDATA,
	qsort_31_s_axi_control_RRESP,
	qsort_31_s_axi_control_AWREADY,
	qsort_31_s_axi_control_AWVALID,
	qsort_31_s_axi_control_AWADDR,
	qsort_31_s_axi_control_WREADY,
	qsort_31_s_axi_control_WVALID,
	qsort_31_s_axi_control_WDATA,
	qsort_31_s_axi_control_WSTRB,
	qsort_31_s_axi_control_BREADY,
	qsort_31_s_axi_control_BVALID,
	qsort_31_s_axi_control_BRESP,
	qsort_32_m_axi_gmem_ARREADY,
	qsort_32_m_axi_gmem_ARVALID,
	qsort_32_m_axi_gmem_ARID,
	qsort_32_m_axi_gmem_ARADDR,
	qsort_32_m_axi_gmem_ARLEN,
	qsort_32_m_axi_gmem_ARSIZE,
	qsort_32_m_axi_gmem_ARBURST,
	qsort_32_m_axi_gmem_ARLOCK,
	qsort_32_m_axi_gmem_ARCACHE,
	qsort_32_m_axi_gmem_ARPROT,
	qsort_32_m_axi_gmem_ARQOS,
	qsort_32_m_axi_gmem_ARREGION,
	qsort_32_m_axi_gmem_ARUSER,
	qsort_32_m_axi_gmem_RREADY,
	qsort_32_m_axi_gmem_RVALID,
	qsort_32_m_axi_gmem_RID,
	qsort_32_m_axi_gmem_RDATA,
	qsort_32_m_axi_gmem_RRESP,
	qsort_32_m_axi_gmem_RLAST,
	qsort_32_m_axi_gmem_RUSER,
	qsort_32_m_axi_gmem_AWREADY,
	qsort_32_m_axi_gmem_AWVALID,
	qsort_32_m_axi_gmem_AWID,
	qsort_32_m_axi_gmem_AWADDR,
	qsort_32_m_axi_gmem_AWLEN,
	qsort_32_m_axi_gmem_AWSIZE,
	qsort_32_m_axi_gmem_AWBURST,
	qsort_32_m_axi_gmem_AWLOCK,
	qsort_32_m_axi_gmem_AWCACHE,
	qsort_32_m_axi_gmem_AWPROT,
	qsort_32_m_axi_gmem_AWQOS,
	qsort_32_m_axi_gmem_AWREGION,
	qsort_32_m_axi_gmem_AWUSER,
	qsort_32_m_axi_gmem_WREADY,
	qsort_32_m_axi_gmem_WVALID,
	qsort_32_m_axi_gmem_WDATA,
	qsort_32_m_axi_gmem_WSTRB,
	qsort_32_m_axi_gmem_WLAST,
	qsort_32_m_axi_gmem_WUSER,
	qsort_32_m_axi_gmem_BREADY,
	qsort_32_m_axi_gmem_BVALID,
	qsort_32_m_axi_gmem_BID,
	qsort_32_m_axi_gmem_BRESP,
	qsort_32_m_axi_gmem_BUSER,
	qsort_32_s_axi_control_ARREADY,
	qsort_32_s_axi_control_ARVALID,
	qsort_32_s_axi_control_ARADDR,
	qsort_32_s_axi_control_RREADY,
	qsort_32_s_axi_control_RVALID,
	qsort_32_s_axi_control_RDATA,
	qsort_32_s_axi_control_RRESP,
	qsort_32_s_axi_control_AWREADY,
	qsort_32_s_axi_control_AWVALID,
	qsort_32_s_axi_control_AWADDR,
	qsort_32_s_axi_control_WREADY,
	qsort_32_s_axi_control_WVALID,
	qsort_32_s_axi_control_WDATA,
	qsort_32_s_axi_control_WSTRB,
	qsort_32_s_axi_control_BREADY,
	qsort_32_s_axi_control_BVALID,
	qsort_32_s_axi_control_BRESP,
	qsort_33_m_axi_gmem_ARREADY,
	qsort_33_m_axi_gmem_ARVALID,
	qsort_33_m_axi_gmem_ARID,
	qsort_33_m_axi_gmem_ARADDR,
	qsort_33_m_axi_gmem_ARLEN,
	qsort_33_m_axi_gmem_ARSIZE,
	qsort_33_m_axi_gmem_ARBURST,
	qsort_33_m_axi_gmem_ARLOCK,
	qsort_33_m_axi_gmem_ARCACHE,
	qsort_33_m_axi_gmem_ARPROT,
	qsort_33_m_axi_gmem_ARQOS,
	qsort_33_m_axi_gmem_ARREGION,
	qsort_33_m_axi_gmem_ARUSER,
	qsort_33_m_axi_gmem_RREADY,
	qsort_33_m_axi_gmem_RVALID,
	qsort_33_m_axi_gmem_RID,
	qsort_33_m_axi_gmem_RDATA,
	qsort_33_m_axi_gmem_RRESP,
	qsort_33_m_axi_gmem_RLAST,
	qsort_33_m_axi_gmem_RUSER,
	qsort_33_m_axi_gmem_AWREADY,
	qsort_33_m_axi_gmem_AWVALID,
	qsort_33_m_axi_gmem_AWID,
	qsort_33_m_axi_gmem_AWADDR,
	qsort_33_m_axi_gmem_AWLEN,
	qsort_33_m_axi_gmem_AWSIZE,
	qsort_33_m_axi_gmem_AWBURST,
	qsort_33_m_axi_gmem_AWLOCK,
	qsort_33_m_axi_gmem_AWCACHE,
	qsort_33_m_axi_gmem_AWPROT,
	qsort_33_m_axi_gmem_AWQOS,
	qsort_33_m_axi_gmem_AWREGION,
	qsort_33_m_axi_gmem_AWUSER,
	qsort_33_m_axi_gmem_WREADY,
	qsort_33_m_axi_gmem_WVALID,
	qsort_33_m_axi_gmem_WDATA,
	qsort_33_m_axi_gmem_WSTRB,
	qsort_33_m_axi_gmem_WLAST,
	qsort_33_m_axi_gmem_WUSER,
	qsort_33_m_axi_gmem_BREADY,
	qsort_33_m_axi_gmem_BVALID,
	qsort_33_m_axi_gmem_BID,
	qsort_33_m_axi_gmem_BRESP,
	qsort_33_m_axi_gmem_BUSER,
	qsort_33_s_axi_control_ARREADY,
	qsort_33_s_axi_control_ARVALID,
	qsort_33_s_axi_control_ARADDR,
	qsort_33_s_axi_control_RREADY,
	qsort_33_s_axi_control_RVALID,
	qsort_33_s_axi_control_RDATA,
	qsort_33_s_axi_control_RRESP,
	qsort_33_s_axi_control_AWREADY,
	qsort_33_s_axi_control_AWVALID,
	qsort_33_s_axi_control_AWADDR,
	qsort_33_s_axi_control_WREADY,
	qsort_33_s_axi_control_WVALID,
	qsort_33_s_axi_control_WDATA,
	qsort_33_s_axi_control_WSTRB,
	qsort_33_s_axi_control_BREADY,
	qsort_33_s_axi_control_BVALID,
	qsort_33_s_axi_control_BRESP,
	qsort_34_m_axi_gmem_ARREADY,
	qsort_34_m_axi_gmem_ARVALID,
	qsort_34_m_axi_gmem_ARID,
	qsort_34_m_axi_gmem_ARADDR,
	qsort_34_m_axi_gmem_ARLEN,
	qsort_34_m_axi_gmem_ARSIZE,
	qsort_34_m_axi_gmem_ARBURST,
	qsort_34_m_axi_gmem_ARLOCK,
	qsort_34_m_axi_gmem_ARCACHE,
	qsort_34_m_axi_gmem_ARPROT,
	qsort_34_m_axi_gmem_ARQOS,
	qsort_34_m_axi_gmem_ARREGION,
	qsort_34_m_axi_gmem_ARUSER,
	qsort_34_m_axi_gmem_RREADY,
	qsort_34_m_axi_gmem_RVALID,
	qsort_34_m_axi_gmem_RID,
	qsort_34_m_axi_gmem_RDATA,
	qsort_34_m_axi_gmem_RRESP,
	qsort_34_m_axi_gmem_RLAST,
	qsort_34_m_axi_gmem_RUSER,
	qsort_34_m_axi_gmem_AWREADY,
	qsort_34_m_axi_gmem_AWVALID,
	qsort_34_m_axi_gmem_AWID,
	qsort_34_m_axi_gmem_AWADDR,
	qsort_34_m_axi_gmem_AWLEN,
	qsort_34_m_axi_gmem_AWSIZE,
	qsort_34_m_axi_gmem_AWBURST,
	qsort_34_m_axi_gmem_AWLOCK,
	qsort_34_m_axi_gmem_AWCACHE,
	qsort_34_m_axi_gmem_AWPROT,
	qsort_34_m_axi_gmem_AWQOS,
	qsort_34_m_axi_gmem_AWREGION,
	qsort_34_m_axi_gmem_AWUSER,
	qsort_34_m_axi_gmem_WREADY,
	qsort_34_m_axi_gmem_WVALID,
	qsort_34_m_axi_gmem_WDATA,
	qsort_34_m_axi_gmem_WSTRB,
	qsort_34_m_axi_gmem_WLAST,
	qsort_34_m_axi_gmem_WUSER,
	qsort_34_m_axi_gmem_BREADY,
	qsort_34_m_axi_gmem_BVALID,
	qsort_34_m_axi_gmem_BID,
	qsort_34_m_axi_gmem_BRESP,
	qsort_34_m_axi_gmem_BUSER,
	qsort_34_s_axi_control_ARREADY,
	qsort_34_s_axi_control_ARVALID,
	qsort_34_s_axi_control_ARADDR,
	qsort_34_s_axi_control_RREADY,
	qsort_34_s_axi_control_RVALID,
	qsort_34_s_axi_control_RDATA,
	qsort_34_s_axi_control_RRESP,
	qsort_34_s_axi_control_AWREADY,
	qsort_34_s_axi_control_AWVALID,
	qsort_34_s_axi_control_AWADDR,
	qsort_34_s_axi_control_WREADY,
	qsort_34_s_axi_control_WVALID,
	qsort_34_s_axi_control_WDATA,
	qsort_34_s_axi_control_WSTRB,
	qsort_34_s_axi_control_BREADY,
	qsort_34_s_axi_control_BVALID,
	qsort_34_s_axi_control_BRESP,
	qsort_35_m_axi_gmem_ARREADY,
	qsort_35_m_axi_gmem_ARVALID,
	qsort_35_m_axi_gmem_ARID,
	qsort_35_m_axi_gmem_ARADDR,
	qsort_35_m_axi_gmem_ARLEN,
	qsort_35_m_axi_gmem_ARSIZE,
	qsort_35_m_axi_gmem_ARBURST,
	qsort_35_m_axi_gmem_ARLOCK,
	qsort_35_m_axi_gmem_ARCACHE,
	qsort_35_m_axi_gmem_ARPROT,
	qsort_35_m_axi_gmem_ARQOS,
	qsort_35_m_axi_gmem_ARREGION,
	qsort_35_m_axi_gmem_ARUSER,
	qsort_35_m_axi_gmem_RREADY,
	qsort_35_m_axi_gmem_RVALID,
	qsort_35_m_axi_gmem_RID,
	qsort_35_m_axi_gmem_RDATA,
	qsort_35_m_axi_gmem_RRESP,
	qsort_35_m_axi_gmem_RLAST,
	qsort_35_m_axi_gmem_RUSER,
	qsort_35_m_axi_gmem_AWREADY,
	qsort_35_m_axi_gmem_AWVALID,
	qsort_35_m_axi_gmem_AWID,
	qsort_35_m_axi_gmem_AWADDR,
	qsort_35_m_axi_gmem_AWLEN,
	qsort_35_m_axi_gmem_AWSIZE,
	qsort_35_m_axi_gmem_AWBURST,
	qsort_35_m_axi_gmem_AWLOCK,
	qsort_35_m_axi_gmem_AWCACHE,
	qsort_35_m_axi_gmem_AWPROT,
	qsort_35_m_axi_gmem_AWQOS,
	qsort_35_m_axi_gmem_AWREGION,
	qsort_35_m_axi_gmem_AWUSER,
	qsort_35_m_axi_gmem_WREADY,
	qsort_35_m_axi_gmem_WVALID,
	qsort_35_m_axi_gmem_WDATA,
	qsort_35_m_axi_gmem_WSTRB,
	qsort_35_m_axi_gmem_WLAST,
	qsort_35_m_axi_gmem_WUSER,
	qsort_35_m_axi_gmem_BREADY,
	qsort_35_m_axi_gmem_BVALID,
	qsort_35_m_axi_gmem_BID,
	qsort_35_m_axi_gmem_BRESP,
	qsort_35_m_axi_gmem_BUSER,
	qsort_35_s_axi_control_ARREADY,
	qsort_35_s_axi_control_ARVALID,
	qsort_35_s_axi_control_ARADDR,
	qsort_35_s_axi_control_RREADY,
	qsort_35_s_axi_control_RVALID,
	qsort_35_s_axi_control_RDATA,
	qsort_35_s_axi_control_RRESP,
	qsort_35_s_axi_control_AWREADY,
	qsort_35_s_axi_control_AWVALID,
	qsort_35_s_axi_control_AWADDR,
	qsort_35_s_axi_control_WREADY,
	qsort_35_s_axi_control_WVALID,
	qsort_35_s_axi_control_WDATA,
	qsort_35_s_axi_control_WSTRB,
	qsort_35_s_axi_control_BREADY,
	qsort_35_s_axi_control_BVALID,
	qsort_35_s_axi_control_BRESP,
	qsort_36_m_axi_gmem_ARREADY,
	qsort_36_m_axi_gmem_ARVALID,
	qsort_36_m_axi_gmem_ARID,
	qsort_36_m_axi_gmem_ARADDR,
	qsort_36_m_axi_gmem_ARLEN,
	qsort_36_m_axi_gmem_ARSIZE,
	qsort_36_m_axi_gmem_ARBURST,
	qsort_36_m_axi_gmem_ARLOCK,
	qsort_36_m_axi_gmem_ARCACHE,
	qsort_36_m_axi_gmem_ARPROT,
	qsort_36_m_axi_gmem_ARQOS,
	qsort_36_m_axi_gmem_ARREGION,
	qsort_36_m_axi_gmem_ARUSER,
	qsort_36_m_axi_gmem_RREADY,
	qsort_36_m_axi_gmem_RVALID,
	qsort_36_m_axi_gmem_RID,
	qsort_36_m_axi_gmem_RDATA,
	qsort_36_m_axi_gmem_RRESP,
	qsort_36_m_axi_gmem_RLAST,
	qsort_36_m_axi_gmem_RUSER,
	qsort_36_m_axi_gmem_AWREADY,
	qsort_36_m_axi_gmem_AWVALID,
	qsort_36_m_axi_gmem_AWID,
	qsort_36_m_axi_gmem_AWADDR,
	qsort_36_m_axi_gmem_AWLEN,
	qsort_36_m_axi_gmem_AWSIZE,
	qsort_36_m_axi_gmem_AWBURST,
	qsort_36_m_axi_gmem_AWLOCK,
	qsort_36_m_axi_gmem_AWCACHE,
	qsort_36_m_axi_gmem_AWPROT,
	qsort_36_m_axi_gmem_AWQOS,
	qsort_36_m_axi_gmem_AWREGION,
	qsort_36_m_axi_gmem_AWUSER,
	qsort_36_m_axi_gmem_WREADY,
	qsort_36_m_axi_gmem_WVALID,
	qsort_36_m_axi_gmem_WDATA,
	qsort_36_m_axi_gmem_WSTRB,
	qsort_36_m_axi_gmem_WLAST,
	qsort_36_m_axi_gmem_WUSER,
	qsort_36_m_axi_gmem_BREADY,
	qsort_36_m_axi_gmem_BVALID,
	qsort_36_m_axi_gmem_BID,
	qsort_36_m_axi_gmem_BRESP,
	qsort_36_m_axi_gmem_BUSER,
	qsort_36_s_axi_control_ARREADY,
	qsort_36_s_axi_control_ARVALID,
	qsort_36_s_axi_control_ARADDR,
	qsort_36_s_axi_control_RREADY,
	qsort_36_s_axi_control_RVALID,
	qsort_36_s_axi_control_RDATA,
	qsort_36_s_axi_control_RRESP,
	qsort_36_s_axi_control_AWREADY,
	qsort_36_s_axi_control_AWVALID,
	qsort_36_s_axi_control_AWADDR,
	qsort_36_s_axi_control_WREADY,
	qsort_36_s_axi_control_WVALID,
	qsort_36_s_axi_control_WDATA,
	qsort_36_s_axi_control_WSTRB,
	qsort_36_s_axi_control_BREADY,
	qsort_36_s_axi_control_BVALID,
	qsort_36_s_axi_control_BRESP,
	qsort_37_m_axi_gmem_ARREADY,
	qsort_37_m_axi_gmem_ARVALID,
	qsort_37_m_axi_gmem_ARID,
	qsort_37_m_axi_gmem_ARADDR,
	qsort_37_m_axi_gmem_ARLEN,
	qsort_37_m_axi_gmem_ARSIZE,
	qsort_37_m_axi_gmem_ARBURST,
	qsort_37_m_axi_gmem_ARLOCK,
	qsort_37_m_axi_gmem_ARCACHE,
	qsort_37_m_axi_gmem_ARPROT,
	qsort_37_m_axi_gmem_ARQOS,
	qsort_37_m_axi_gmem_ARREGION,
	qsort_37_m_axi_gmem_ARUSER,
	qsort_37_m_axi_gmem_RREADY,
	qsort_37_m_axi_gmem_RVALID,
	qsort_37_m_axi_gmem_RID,
	qsort_37_m_axi_gmem_RDATA,
	qsort_37_m_axi_gmem_RRESP,
	qsort_37_m_axi_gmem_RLAST,
	qsort_37_m_axi_gmem_RUSER,
	qsort_37_m_axi_gmem_AWREADY,
	qsort_37_m_axi_gmem_AWVALID,
	qsort_37_m_axi_gmem_AWID,
	qsort_37_m_axi_gmem_AWADDR,
	qsort_37_m_axi_gmem_AWLEN,
	qsort_37_m_axi_gmem_AWSIZE,
	qsort_37_m_axi_gmem_AWBURST,
	qsort_37_m_axi_gmem_AWLOCK,
	qsort_37_m_axi_gmem_AWCACHE,
	qsort_37_m_axi_gmem_AWPROT,
	qsort_37_m_axi_gmem_AWQOS,
	qsort_37_m_axi_gmem_AWREGION,
	qsort_37_m_axi_gmem_AWUSER,
	qsort_37_m_axi_gmem_WREADY,
	qsort_37_m_axi_gmem_WVALID,
	qsort_37_m_axi_gmem_WDATA,
	qsort_37_m_axi_gmem_WSTRB,
	qsort_37_m_axi_gmem_WLAST,
	qsort_37_m_axi_gmem_WUSER,
	qsort_37_m_axi_gmem_BREADY,
	qsort_37_m_axi_gmem_BVALID,
	qsort_37_m_axi_gmem_BID,
	qsort_37_m_axi_gmem_BRESP,
	qsort_37_m_axi_gmem_BUSER,
	qsort_37_s_axi_control_ARREADY,
	qsort_37_s_axi_control_ARVALID,
	qsort_37_s_axi_control_ARADDR,
	qsort_37_s_axi_control_RREADY,
	qsort_37_s_axi_control_RVALID,
	qsort_37_s_axi_control_RDATA,
	qsort_37_s_axi_control_RRESP,
	qsort_37_s_axi_control_AWREADY,
	qsort_37_s_axi_control_AWVALID,
	qsort_37_s_axi_control_AWADDR,
	qsort_37_s_axi_control_WREADY,
	qsort_37_s_axi_control_WVALID,
	qsort_37_s_axi_control_WDATA,
	qsort_37_s_axi_control_WSTRB,
	qsort_37_s_axi_control_BREADY,
	qsort_37_s_axi_control_BVALID,
	qsort_37_s_axi_control_BRESP,
	qsort_38_m_axi_gmem_ARREADY,
	qsort_38_m_axi_gmem_ARVALID,
	qsort_38_m_axi_gmem_ARID,
	qsort_38_m_axi_gmem_ARADDR,
	qsort_38_m_axi_gmem_ARLEN,
	qsort_38_m_axi_gmem_ARSIZE,
	qsort_38_m_axi_gmem_ARBURST,
	qsort_38_m_axi_gmem_ARLOCK,
	qsort_38_m_axi_gmem_ARCACHE,
	qsort_38_m_axi_gmem_ARPROT,
	qsort_38_m_axi_gmem_ARQOS,
	qsort_38_m_axi_gmem_ARREGION,
	qsort_38_m_axi_gmem_ARUSER,
	qsort_38_m_axi_gmem_RREADY,
	qsort_38_m_axi_gmem_RVALID,
	qsort_38_m_axi_gmem_RID,
	qsort_38_m_axi_gmem_RDATA,
	qsort_38_m_axi_gmem_RRESP,
	qsort_38_m_axi_gmem_RLAST,
	qsort_38_m_axi_gmem_RUSER,
	qsort_38_m_axi_gmem_AWREADY,
	qsort_38_m_axi_gmem_AWVALID,
	qsort_38_m_axi_gmem_AWID,
	qsort_38_m_axi_gmem_AWADDR,
	qsort_38_m_axi_gmem_AWLEN,
	qsort_38_m_axi_gmem_AWSIZE,
	qsort_38_m_axi_gmem_AWBURST,
	qsort_38_m_axi_gmem_AWLOCK,
	qsort_38_m_axi_gmem_AWCACHE,
	qsort_38_m_axi_gmem_AWPROT,
	qsort_38_m_axi_gmem_AWQOS,
	qsort_38_m_axi_gmem_AWREGION,
	qsort_38_m_axi_gmem_AWUSER,
	qsort_38_m_axi_gmem_WREADY,
	qsort_38_m_axi_gmem_WVALID,
	qsort_38_m_axi_gmem_WDATA,
	qsort_38_m_axi_gmem_WSTRB,
	qsort_38_m_axi_gmem_WLAST,
	qsort_38_m_axi_gmem_WUSER,
	qsort_38_m_axi_gmem_BREADY,
	qsort_38_m_axi_gmem_BVALID,
	qsort_38_m_axi_gmem_BID,
	qsort_38_m_axi_gmem_BRESP,
	qsort_38_m_axi_gmem_BUSER,
	qsort_38_s_axi_control_ARREADY,
	qsort_38_s_axi_control_ARVALID,
	qsort_38_s_axi_control_ARADDR,
	qsort_38_s_axi_control_RREADY,
	qsort_38_s_axi_control_RVALID,
	qsort_38_s_axi_control_RDATA,
	qsort_38_s_axi_control_RRESP,
	qsort_38_s_axi_control_AWREADY,
	qsort_38_s_axi_control_AWVALID,
	qsort_38_s_axi_control_AWADDR,
	qsort_38_s_axi_control_WREADY,
	qsort_38_s_axi_control_WVALID,
	qsort_38_s_axi_control_WDATA,
	qsort_38_s_axi_control_WSTRB,
	qsort_38_s_axi_control_BREADY,
	qsort_38_s_axi_control_BVALID,
	qsort_38_s_axi_control_BRESP,
	qsort_39_m_axi_gmem_ARREADY,
	qsort_39_m_axi_gmem_ARVALID,
	qsort_39_m_axi_gmem_ARID,
	qsort_39_m_axi_gmem_ARADDR,
	qsort_39_m_axi_gmem_ARLEN,
	qsort_39_m_axi_gmem_ARSIZE,
	qsort_39_m_axi_gmem_ARBURST,
	qsort_39_m_axi_gmem_ARLOCK,
	qsort_39_m_axi_gmem_ARCACHE,
	qsort_39_m_axi_gmem_ARPROT,
	qsort_39_m_axi_gmem_ARQOS,
	qsort_39_m_axi_gmem_ARREGION,
	qsort_39_m_axi_gmem_ARUSER,
	qsort_39_m_axi_gmem_RREADY,
	qsort_39_m_axi_gmem_RVALID,
	qsort_39_m_axi_gmem_RID,
	qsort_39_m_axi_gmem_RDATA,
	qsort_39_m_axi_gmem_RRESP,
	qsort_39_m_axi_gmem_RLAST,
	qsort_39_m_axi_gmem_RUSER,
	qsort_39_m_axi_gmem_AWREADY,
	qsort_39_m_axi_gmem_AWVALID,
	qsort_39_m_axi_gmem_AWID,
	qsort_39_m_axi_gmem_AWADDR,
	qsort_39_m_axi_gmem_AWLEN,
	qsort_39_m_axi_gmem_AWSIZE,
	qsort_39_m_axi_gmem_AWBURST,
	qsort_39_m_axi_gmem_AWLOCK,
	qsort_39_m_axi_gmem_AWCACHE,
	qsort_39_m_axi_gmem_AWPROT,
	qsort_39_m_axi_gmem_AWQOS,
	qsort_39_m_axi_gmem_AWREGION,
	qsort_39_m_axi_gmem_AWUSER,
	qsort_39_m_axi_gmem_WREADY,
	qsort_39_m_axi_gmem_WVALID,
	qsort_39_m_axi_gmem_WDATA,
	qsort_39_m_axi_gmem_WSTRB,
	qsort_39_m_axi_gmem_WLAST,
	qsort_39_m_axi_gmem_WUSER,
	qsort_39_m_axi_gmem_BREADY,
	qsort_39_m_axi_gmem_BVALID,
	qsort_39_m_axi_gmem_BID,
	qsort_39_m_axi_gmem_BRESP,
	qsort_39_m_axi_gmem_BUSER,
	qsort_39_s_axi_control_ARREADY,
	qsort_39_s_axi_control_ARVALID,
	qsort_39_s_axi_control_ARADDR,
	qsort_39_s_axi_control_RREADY,
	qsort_39_s_axi_control_RVALID,
	qsort_39_s_axi_control_RDATA,
	qsort_39_s_axi_control_RRESP,
	qsort_39_s_axi_control_AWREADY,
	qsort_39_s_axi_control_AWVALID,
	qsort_39_s_axi_control_AWADDR,
	qsort_39_s_axi_control_WREADY,
	qsort_39_s_axi_control_WVALID,
	qsort_39_s_axi_control_WDATA,
	qsort_39_s_axi_control_WSTRB,
	qsort_39_s_axi_control_BREADY,
	qsort_39_s_axi_control_BVALID,
	qsort_39_s_axi_control_BRESP,
	qsort_40_m_axi_gmem_ARREADY,
	qsort_40_m_axi_gmem_ARVALID,
	qsort_40_m_axi_gmem_ARID,
	qsort_40_m_axi_gmem_ARADDR,
	qsort_40_m_axi_gmem_ARLEN,
	qsort_40_m_axi_gmem_ARSIZE,
	qsort_40_m_axi_gmem_ARBURST,
	qsort_40_m_axi_gmem_ARLOCK,
	qsort_40_m_axi_gmem_ARCACHE,
	qsort_40_m_axi_gmem_ARPROT,
	qsort_40_m_axi_gmem_ARQOS,
	qsort_40_m_axi_gmem_ARREGION,
	qsort_40_m_axi_gmem_ARUSER,
	qsort_40_m_axi_gmem_RREADY,
	qsort_40_m_axi_gmem_RVALID,
	qsort_40_m_axi_gmem_RID,
	qsort_40_m_axi_gmem_RDATA,
	qsort_40_m_axi_gmem_RRESP,
	qsort_40_m_axi_gmem_RLAST,
	qsort_40_m_axi_gmem_RUSER,
	qsort_40_m_axi_gmem_AWREADY,
	qsort_40_m_axi_gmem_AWVALID,
	qsort_40_m_axi_gmem_AWID,
	qsort_40_m_axi_gmem_AWADDR,
	qsort_40_m_axi_gmem_AWLEN,
	qsort_40_m_axi_gmem_AWSIZE,
	qsort_40_m_axi_gmem_AWBURST,
	qsort_40_m_axi_gmem_AWLOCK,
	qsort_40_m_axi_gmem_AWCACHE,
	qsort_40_m_axi_gmem_AWPROT,
	qsort_40_m_axi_gmem_AWQOS,
	qsort_40_m_axi_gmem_AWREGION,
	qsort_40_m_axi_gmem_AWUSER,
	qsort_40_m_axi_gmem_WREADY,
	qsort_40_m_axi_gmem_WVALID,
	qsort_40_m_axi_gmem_WDATA,
	qsort_40_m_axi_gmem_WSTRB,
	qsort_40_m_axi_gmem_WLAST,
	qsort_40_m_axi_gmem_WUSER,
	qsort_40_m_axi_gmem_BREADY,
	qsort_40_m_axi_gmem_BVALID,
	qsort_40_m_axi_gmem_BID,
	qsort_40_m_axi_gmem_BRESP,
	qsort_40_m_axi_gmem_BUSER,
	qsort_40_s_axi_control_ARREADY,
	qsort_40_s_axi_control_ARVALID,
	qsort_40_s_axi_control_ARADDR,
	qsort_40_s_axi_control_RREADY,
	qsort_40_s_axi_control_RVALID,
	qsort_40_s_axi_control_RDATA,
	qsort_40_s_axi_control_RRESP,
	qsort_40_s_axi_control_AWREADY,
	qsort_40_s_axi_control_AWVALID,
	qsort_40_s_axi_control_AWADDR,
	qsort_40_s_axi_control_WREADY,
	qsort_40_s_axi_control_WVALID,
	qsort_40_s_axi_control_WDATA,
	qsort_40_s_axi_control_WSTRB,
	qsort_40_s_axi_control_BREADY,
	qsort_40_s_axi_control_BVALID,
	qsort_40_s_axi_control_BRESP,
	qsort_41_m_axi_gmem_ARREADY,
	qsort_41_m_axi_gmem_ARVALID,
	qsort_41_m_axi_gmem_ARID,
	qsort_41_m_axi_gmem_ARADDR,
	qsort_41_m_axi_gmem_ARLEN,
	qsort_41_m_axi_gmem_ARSIZE,
	qsort_41_m_axi_gmem_ARBURST,
	qsort_41_m_axi_gmem_ARLOCK,
	qsort_41_m_axi_gmem_ARCACHE,
	qsort_41_m_axi_gmem_ARPROT,
	qsort_41_m_axi_gmem_ARQOS,
	qsort_41_m_axi_gmem_ARREGION,
	qsort_41_m_axi_gmem_ARUSER,
	qsort_41_m_axi_gmem_RREADY,
	qsort_41_m_axi_gmem_RVALID,
	qsort_41_m_axi_gmem_RID,
	qsort_41_m_axi_gmem_RDATA,
	qsort_41_m_axi_gmem_RRESP,
	qsort_41_m_axi_gmem_RLAST,
	qsort_41_m_axi_gmem_RUSER,
	qsort_41_m_axi_gmem_AWREADY,
	qsort_41_m_axi_gmem_AWVALID,
	qsort_41_m_axi_gmem_AWID,
	qsort_41_m_axi_gmem_AWADDR,
	qsort_41_m_axi_gmem_AWLEN,
	qsort_41_m_axi_gmem_AWSIZE,
	qsort_41_m_axi_gmem_AWBURST,
	qsort_41_m_axi_gmem_AWLOCK,
	qsort_41_m_axi_gmem_AWCACHE,
	qsort_41_m_axi_gmem_AWPROT,
	qsort_41_m_axi_gmem_AWQOS,
	qsort_41_m_axi_gmem_AWREGION,
	qsort_41_m_axi_gmem_AWUSER,
	qsort_41_m_axi_gmem_WREADY,
	qsort_41_m_axi_gmem_WVALID,
	qsort_41_m_axi_gmem_WDATA,
	qsort_41_m_axi_gmem_WSTRB,
	qsort_41_m_axi_gmem_WLAST,
	qsort_41_m_axi_gmem_WUSER,
	qsort_41_m_axi_gmem_BREADY,
	qsort_41_m_axi_gmem_BVALID,
	qsort_41_m_axi_gmem_BID,
	qsort_41_m_axi_gmem_BRESP,
	qsort_41_m_axi_gmem_BUSER,
	qsort_41_s_axi_control_ARREADY,
	qsort_41_s_axi_control_ARVALID,
	qsort_41_s_axi_control_ARADDR,
	qsort_41_s_axi_control_RREADY,
	qsort_41_s_axi_control_RVALID,
	qsort_41_s_axi_control_RDATA,
	qsort_41_s_axi_control_RRESP,
	qsort_41_s_axi_control_AWREADY,
	qsort_41_s_axi_control_AWVALID,
	qsort_41_s_axi_control_AWADDR,
	qsort_41_s_axi_control_WREADY,
	qsort_41_s_axi_control_WVALID,
	qsort_41_s_axi_control_WDATA,
	qsort_41_s_axi_control_WSTRB,
	qsort_41_s_axi_control_BREADY,
	qsort_41_s_axi_control_BVALID,
	qsort_41_s_axi_control_BRESP,
	qsort_42_m_axi_gmem_ARREADY,
	qsort_42_m_axi_gmem_ARVALID,
	qsort_42_m_axi_gmem_ARID,
	qsort_42_m_axi_gmem_ARADDR,
	qsort_42_m_axi_gmem_ARLEN,
	qsort_42_m_axi_gmem_ARSIZE,
	qsort_42_m_axi_gmem_ARBURST,
	qsort_42_m_axi_gmem_ARLOCK,
	qsort_42_m_axi_gmem_ARCACHE,
	qsort_42_m_axi_gmem_ARPROT,
	qsort_42_m_axi_gmem_ARQOS,
	qsort_42_m_axi_gmem_ARREGION,
	qsort_42_m_axi_gmem_ARUSER,
	qsort_42_m_axi_gmem_RREADY,
	qsort_42_m_axi_gmem_RVALID,
	qsort_42_m_axi_gmem_RID,
	qsort_42_m_axi_gmem_RDATA,
	qsort_42_m_axi_gmem_RRESP,
	qsort_42_m_axi_gmem_RLAST,
	qsort_42_m_axi_gmem_RUSER,
	qsort_42_m_axi_gmem_AWREADY,
	qsort_42_m_axi_gmem_AWVALID,
	qsort_42_m_axi_gmem_AWID,
	qsort_42_m_axi_gmem_AWADDR,
	qsort_42_m_axi_gmem_AWLEN,
	qsort_42_m_axi_gmem_AWSIZE,
	qsort_42_m_axi_gmem_AWBURST,
	qsort_42_m_axi_gmem_AWLOCK,
	qsort_42_m_axi_gmem_AWCACHE,
	qsort_42_m_axi_gmem_AWPROT,
	qsort_42_m_axi_gmem_AWQOS,
	qsort_42_m_axi_gmem_AWREGION,
	qsort_42_m_axi_gmem_AWUSER,
	qsort_42_m_axi_gmem_WREADY,
	qsort_42_m_axi_gmem_WVALID,
	qsort_42_m_axi_gmem_WDATA,
	qsort_42_m_axi_gmem_WSTRB,
	qsort_42_m_axi_gmem_WLAST,
	qsort_42_m_axi_gmem_WUSER,
	qsort_42_m_axi_gmem_BREADY,
	qsort_42_m_axi_gmem_BVALID,
	qsort_42_m_axi_gmem_BID,
	qsort_42_m_axi_gmem_BRESP,
	qsort_42_m_axi_gmem_BUSER,
	qsort_42_s_axi_control_ARREADY,
	qsort_42_s_axi_control_ARVALID,
	qsort_42_s_axi_control_ARADDR,
	qsort_42_s_axi_control_RREADY,
	qsort_42_s_axi_control_RVALID,
	qsort_42_s_axi_control_RDATA,
	qsort_42_s_axi_control_RRESP,
	qsort_42_s_axi_control_AWREADY,
	qsort_42_s_axi_control_AWVALID,
	qsort_42_s_axi_control_AWADDR,
	qsort_42_s_axi_control_WREADY,
	qsort_42_s_axi_control_WVALID,
	qsort_42_s_axi_control_WDATA,
	qsort_42_s_axi_control_WSTRB,
	qsort_42_s_axi_control_BREADY,
	qsort_42_s_axi_control_BVALID,
	qsort_42_s_axi_control_BRESP,
	qsort_43_m_axi_gmem_ARREADY,
	qsort_43_m_axi_gmem_ARVALID,
	qsort_43_m_axi_gmem_ARID,
	qsort_43_m_axi_gmem_ARADDR,
	qsort_43_m_axi_gmem_ARLEN,
	qsort_43_m_axi_gmem_ARSIZE,
	qsort_43_m_axi_gmem_ARBURST,
	qsort_43_m_axi_gmem_ARLOCK,
	qsort_43_m_axi_gmem_ARCACHE,
	qsort_43_m_axi_gmem_ARPROT,
	qsort_43_m_axi_gmem_ARQOS,
	qsort_43_m_axi_gmem_ARREGION,
	qsort_43_m_axi_gmem_ARUSER,
	qsort_43_m_axi_gmem_RREADY,
	qsort_43_m_axi_gmem_RVALID,
	qsort_43_m_axi_gmem_RID,
	qsort_43_m_axi_gmem_RDATA,
	qsort_43_m_axi_gmem_RRESP,
	qsort_43_m_axi_gmem_RLAST,
	qsort_43_m_axi_gmem_RUSER,
	qsort_43_m_axi_gmem_AWREADY,
	qsort_43_m_axi_gmem_AWVALID,
	qsort_43_m_axi_gmem_AWID,
	qsort_43_m_axi_gmem_AWADDR,
	qsort_43_m_axi_gmem_AWLEN,
	qsort_43_m_axi_gmem_AWSIZE,
	qsort_43_m_axi_gmem_AWBURST,
	qsort_43_m_axi_gmem_AWLOCK,
	qsort_43_m_axi_gmem_AWCACHE,
	qsort_43_m_axi_gmem_AWPROT,
	qsort_43_m_axi_gmem_AWQOS,
	qsort_43_m_axi_gmem_AWREGION,
	qsort_43_m_axi_gmem_AWUSER,
	qsort_43_m_axi_gmem_WREADY,
	qsort_43_m_axi_gmem_WVALID,
	qsort_43_m_axi_gmem_WDATA,
	qsort_43_m_axi_gmem_WSTRB,
	qsort_43_m_axi_gmem_WLAST,
	qsort_43_m_axi_gmem_WUSER,
	qsort_43_m_axi_gmem_BREADY,
	qsort_43_m_axi_gmem_BVALID,
	qsort_43_m_axi_gmem_BID,
	qsort_43_m_axi_gmem_BRESP,
	qsort_43_m_axi_gmem_BUSER,
	qsort_43_s_axi_control_ARREADY,
	qsort_43_s_axi_control_ARVALID,
	qsort_43_s_axi_control_ARADDR,
	qsort_43_s_axi_control_RREADY,
	qsort_43_s_axi_control_RVALID,
	qsort_43_s_axi_control_RDATA,
	qsort_43_s_axi_control_RRESP,
	qsort_43_s_axi_control_AWREADY,
	qsort_43_s_axi_control_AWVALID,
	qsort_43_s_axi_control_AWADDR,
	qsort_43_s_axi_control_WREADY,
	qsort_43_s_axi_control_WVALID,
	qsort_43_s_axi_control_WDATA,
	qsort_43_s_axi_control_WSTRB,
	qsort_43_s_axi_control_BREADY,
	qsort_43_s_axi_control_BVALID,
	qsort_43_s_axi_control_BRESP,
	qsort_44_m_axi_gmem_ARREADY,
	qsort_44_m_axi_gmem_ARVALID,
	qsort_44_m_axi_gmem_ARID,
	qsort_44_m_axi_gmem_ARADDR,
	qsort_44_m_axi_gmem_ARLEN,
	qsort_44_m_axi_gmem_ARSIZE,
	qsort_44_m_axi_gmem_ARBURST,
	qsort_44_m_axi_gmem_ARLOCK,
	qsort_44_m_axi_gmem_ARCACHE,
	qsort_44_m_axi_gmem_ARPROT,
	qsort_44_m_axi_gmem_ARQOS,
	qsort_44_m_axi_gmem_ARREGION,
	qsort_44_m_axi_gmem_ARUSER,
	qsort_44_m_axi_gmem_RREADY,
	qsort_44_m_axi_gmem_RVALID,
	qsort_44_m_axi_gmem_RID,
	qsort_44_m_axi_gmem_RDATA,
	qsort_44_m_axi_gmem_RRESP,
	qsort_44_m_axi_gmem_RLAST,
	qsort_44_m_axi_gmem_RUSER,
	qsort_44_m_axi_gmem_AWREADY,
	qsort_44_m_axi_gmem_AWVALID,
	qsort_44_m_axi_gmem_AWID,
	qsort_44_m_axi_gmem_AWADDR,
	qsort_44_m_axi_gmem_AWLEN,
	qsort_44_m_axi_gmem_AWSIZE,
	qsort_44_m_axi_gmem_AWBURST,
	qsort_44_m_axi_gmem_AWLOCK,
	qsort_44_m_axi_gmem_AWCACHE,
	qsort_44_m_axi_gmem_AWPROT,
	qsort_44_m_axi_gmem_AWQOS,
	qsort_44_m_axi_gmem_AWREGION,
	qsort_44_m_axi_gmem_AWUSER,
	qsort_44_m_axi_gmem_WREADY,
	qsort_44_m_axi_gmem_WVALID,
	qsort_44_m_axi_gmem_WDATA,
	qsort_44_m_axi_gmem_WSTRB,
	qsort_44_m_axi_gmem_WLAST,
	qsort_44_m_axi_gmem_WUSER,
	qsort_44_m_axi_gmem_BREADY,
	qsort_44_m_axi_gmem_BVALID,
	qsort_44_m_axi_gmem_BID,
	qsort_44_m_axi_gmem_BRESP,
	qsort_44_m_axi_gmem_BUSER,
	qsort_44_s_axi_control_ARREADY,
	qsort_44_s_axi_control_ARVALID,
	qsort_44_s_axi_control_ARADDR,
	qsort_44_s_axi_control_RREADY,
	qsort_44_s_axi_control_RVALID,
	qsort_44_s_axi_control_RDATA,
	qsort_44_s_axi_control_RRESP,
	qsort_44_s_axi_control_AWREADY,
	qsort_44_s_axi_control_AWVALID,
	qsort_44_s_axi_control_AWADDR,
	qsort_44_s_axi_control_WREADY,
	qsort_44_s_axi_control_WVALID,
	qsort_44_s_axi_control_WDATA,
	qsort_44_s_axi_control_WSTRB,
	qsort_44_s_axi_control_BREADY,
	qsort_44_s_axi_control_BVALID,
	qsort_44_s_axi_control_BRESP,
	qsort_45_m_axi_gmem_ARREADY,
	qsort_45_m_axi_gmem_ARVALID,
	qsort_45_m_axi_gmem_ARID,
	qsort_45_m_axi_gmem_ARADDR,
	qsort_45_m_axi_gmem_ARLEN,
	qsort_45_m_axi_gmem_ARSIZE,
	qsort_45_m_axi_gmem_ARBURST,
	qsort_45_m_axi_gmem_ARLOCK,
	qsort_45_m_axi_gmem_ARCACHE,
	qsort_45_m_axi_gmem_ARPROT,
	qsort_45_m_axi_gmem_ARQOS,
	qsort_45_m_axi_gmem_ARREGION,
	qsort_45_m_axi_gmem_ARUSER,
	qsort_45_m_axi_gmem_RREADY,
	qsort_45_m_axi_gmem_RVALID,
	qsort_45_m_axi_gmem_RID,
	qsort_45_m_axi_gmem_RDATA,
	qsort_45_m_axi_gmem_RRESP,
	qsort_45_m_axi_gmem_RLAST,
	qsort_45_m_axi_gmem_RUSER,
	qsort_45_m_axi_gmem_AWREADY,
	qsort_45_m_axi_gmem_AWVALID,
	qsort_45_m_axi_gmem_AWID,
	qsort_45_m_axi_gmem_AWADDR,
	qsort_45_m_axi_gmem_AWLEN,
	qsort_45_m_axi_gmem_AWSIZE,
	qsort_45_m_axi_gmem_AWBURST,
	qsort_45_m_axi_gmem_AWLOCK,
	qsort_45_m_axi_gmem_AWCACHE,
	qsort_45_m_axi_gmem_AWPROT,
	qsort_45_m_axi_gmem_AWQOS,
	qsort_45_m_axi_gmem_AWREGION,
	qsort_45_m_axi_gmem_AWUSER,
	qsort_45_m_axi_gmem_WREADY,
	qsort_45_m_axi_gmem_WVALID,
	qsort_45_m_axi_gmem_WDATA,
	qsort_45_m_axi_gmem_WSTRB,
	qsort_45_m_axi_gmem_WLAST,
	qsort_45_m_axi_gmem_WUSER,
	qsort_45_m_axi_gmem_BREADY,
	qsort_45_m_axi_gmem_BVALID,
	qsort_45_m_axi_gmem_BID,
	qsort_45_m_axi_gmem_BRESP,
	qsort_45_m_axi_gmem_BUSER,
	qsort_45_s_axi_control_ARREADY,
	qsort_45_s_axi_control_ARVALID,
	qsort_45_s_axi_control_ARADDR,
	qsort_45_s_axi_control_RREADY,
	qsort_45_s_axi_control_RVALID,
	qsort_45_s_axi_control_RDATA,
	qsort_45_s_axi_control_RRESP,
	qsort_45_s_axi_control_AWREADY,
	qsort_45_s_axi_control_AWVALID,
	qsort_45_s_axi_control_AWADDR,
	qsort_45_s_axi_control_WREADY,
	qsort_45_s_axi_control_WVALID,
	qsort_45_s_axi_control_WDATA,
	qsort_45_s_axi_control_WSTRB,
	qsort_45_s_axi_control_BREADY,
	qsort_45_s_axi_control_BVALID,
	qsort_45_s_axi_control_BRESP,
	qsort_46_m_axi_gmem_ARREADY,
	qsort_46_m_axi_gmem_ARVALID,
	qsort_46_m_axi_gmem_ARID,
	qsort_46_m_axi_gmem_ARADDR,
	qsort_46_m_axi_gmem_ARLEN,
	qsort_46_m_axi_gmem_ARSIZE,
	qsort_46_m_axi_gmem_ARBURST,
	qsort_46_m_axi_gmem_ARLOCK,
	qsort_46_m_axi_gmem_ARCACHE,
	qsort_46_m_axi_gmem_ARPROT,
	qsort_46_m_axi_gmem_ARQOS,
	qsort_46_m_axi_gmem_ARREGION,
	qsort_46_m_axi_gmem_ARUSER,
	qsort_46_m_axi_gmem_RREADY,
	qsort_46_m_axi_gmem_RVALID,
	qsort_46_m_axi_gmem_RID,
	qsort_46_m_axi_gmem_RDATA,
	qsort_46_m_axi_gmem_RRESP,
	qsort_46_m_axi_gmem_RLAST,
	qsort_46_m_axi_gmem_RUSER,
	qsort_46_m_axi_gmem_AWREADY,
	qsort_46_m_axi_gmem_AWVALID,
	qsort_46_m_axi_gmem_AWID,
	qsort_46_m_axi_gmem_AWADDR,
	qsort_46_m_axi_gmem_AWLEN,
	qsort_46_m_axi_gmem_AWSIZE,
	qsort_46_m_axi_gmem_AWBURST,
	qsort_46_m_axi_gmem_AWLOCK,
	qsort_46_m_axi_gmem_AWCACHE,
	qsort_46_m_axi_gmem_AWPROT,
	qsort_46_m_axi_gmem_AWQOS,
	qsort_46_m_axi_gmem_AWREGION,
	qsort_46_m_axi_gmem_AWUSER,
	qsort_46_m_axi_gmem_WREADY,
	qsort_46_m_axi_gmem_WVALID,
	qsort_46_m_axi_gmem_WDATA,
	qsort_46_m_axi_gmem_WSTRB,
	qsort_46_m_axi_gmem_WLAST,
	qsort_46_m_axi_gmem_WUSER,
	qsort_46_m_axi_gmem_BREADY,
	qsort_46_m_axi_gmem_BVALID,
	qsort_46_m_axi_gmem_BID,
	qsort_46_m_axi_gmem_BRESP,
	qsort_46_m_axi_gmem_BUSER,
	qsort_46_s_axi_control_ARREADY,
	qsort_46_s_axi_control_ARVALID,
	qsort_46_s_axi_control_ARADDR,
	qsort_46_s_axi_control_RREADY,
	qsort_46_s_axi_control_RVALID,
	qsort_46_s_axi_control_RDATA,
	qsort_46_s_axi_control_RRESP,
	qsort_46_s_axi_control_AWREADY,
	qsort_46_s_axi_control_AWVALID,
	qsort_46_s_axi_control_AWADDR,
	qsort_46_s_axi_control_WREADY,
	qsort_46_s_axi_control_WVALID,
	qsort_46_s_axi_control_WDATA,
	qsort_46_s_axi_control_WSTRB,
	qsort_46_s_axi_control_BREADY,
	qsort_46_s_axi_control_BVALID,
	qsort_46_s_axi_control_BRESP,
	qsort_47_m_axi_gmem_ARREADY,
	qsort_47_m_axi_gmem_ARVALID,
	qsort_47_m_axi_gmem_ARID,
	qsort_47_m_axi_gmem_ARADDR,
	qsort_47_m_axi_gmem_ARLEN,
	qsort_47_m_axi_gmem_ARSIZE,
	qsort_47_m_axi_gmem_ARBURST,
	qsort_47_m_axi_gmem_ARLOCK,
	qsort_47_m_axi_gmem_ARCACHE,
	qsort_47_m_axi_gmem_ARPROT,
	qsort_47_m_axi_gmem_ARQOS,
	qsort_47_m_axi_gmem_ARREGION,
	qsort_47_m_axi_gmem_ARUSER,
	qsort_47_m_axi_gmem_RREADY,
	qsort_47_m_axi_gmem_RVALID,
	qsort_47_m_axi_gmem_RID,
	qsort_47_m_axi_gmem_RDATA,
	qsort_47_m_axi_gmem_RRESP,
	qsort_47_m_axi_gmem_RLAST,
	qsort_47_m_axi_gmem_RUSER,
	qsort_47_m_axi_gmem_AWREADY,
	qsort_47_m_axi_gmem_AWVALID,
	qsort_47_m_axi_gmem_AWID,
	qsort_47_m_axi_gmem_AWADDR,
	qsort_47_m_axi_gmem_AWLEN,
	qsort_47_m_axi_gmem_AWSIZE,
	qsort_47_m_axi_gmem_AWBURST,
	qsort_47_m_axi_gmem_AWLOCK,
	qsort_47_m_axi_gmem_AWCACHE,
	qsort_47_m_axi_gmem_AWPROT,
	qsort_47_m_axi_gmem_AWQOS,
	qsort_47_m_axi_gmem_AWREGION,
	qsort_47_m_axi_gmem_AWUSER,
	qsort_47_m_axi_gmem_WREADY,
	qsort_47_m_axi_gmem_WVALID,
	qsort_47_m_axi_gmem_WDATA,
	qsort_47_m_axi_gmem_WSTRB,
	qsort_47_m_axi_gmem_WLAST,
	qsort_47_m_axi_gmem_WUSER,
	qsort_47_m_axi_gmem_BREADY,
	qsort_47_m_axi_gmem_BVALID,
	qsort_47_m_axi_gmem_BID,
	qsort_47_m_axi_gmem_BRESP,
	qsort_47_m_axi_gmem_BUSER,
	qsort_47_s_axi_control_ARREADY,
	qsort_47_s_axi_control_ARVALID,
	qsort_47_s_axi_control_ARADDR,
	qsort_47_s_axi_control_RREADY,
	qsort_47_s_axi_control_RVALID,
	qsort_47_s_axi_control_RDATA,
	qsort_47_s_axi_control_RRESP,
	qsort_47_s_axi_control_AWREADY,
	qsort_47_s_axi_control_AWVALID,
	qsort_47_s_axi_control_AWADDR,
	qsort_47_s_axi_control_WREADY,
	qsort_47_s_axi_control_WVALID,
	qsort_47_s_axi_control_WDATA,
	qsort_47_s_axi_control_WSTRB,
	qsort_47_s_axi_control_BREADY,
	qsort_47_s_axi_control_BVALID,
	qsort_47_s_axi_control_BRESP,
	qsort_48_m_axi_gmem_ARREADY,
	qsort_48_m_axi_gmem_ARVALID,
	qsort_48_m_axi_gmem_ARID,
	qsort_48_m_axi_gmem_ARADDR,
	qsort_48_m_axi_gmem_ARLEN,
	qsort_48_m_axi_gmem_ARSIZE,
	qsort_48_m_axi_gmem_ARBURST,
	qsort_48_m_axi_gmem_ARLOCK,
	qsort_48_m_axi_gmem_ARCACHE,
	qsort_48_m_axi_gmem_ARPROT,
	qsort_48_m_axi_gmem_ARQOS,
	qsort_48_m_axi_gmem_ARREGION,
	qsort_48_m_axi_gmem_ARUSER,
	qsort_48_m_axi_gmem_RREADY,
	qsort_48_m_axi_gmem_RVALID,
	qsort_48_m_axi_gmem_RID,
	qsort_48_m_axi_gmem_RDATA,
	qsort_48_m_axi_gmem_RRESP,
	qsort_48_m_axi_gmem_RLAST,
	qsort_48_m_axi_gmem_RUSER,
	qsort_48_m_axi_gmem_AWREADY,
	qsort_48_m_axi_gmem_AWVALID,
	qsort_48_m_axi_gmem_AWID,
	qsort_48_m_axi_gmem_AWADDR,
	qsort_48_m_axi_gmem_AWLEN,
	qsort_48_m_axi_gmem_AWSIZE,
	qsort_48_m_axi_gmem_AWBURST,
	qsort_48_m_axi_gmem_AWLOCK,
	qsort_48_m_axi_gmem_AWCACHE,
	qsort_48_m_axi_gmem_AWPROT,
	qsort_48_m_axi_gmem_AWQOS,
	qsort_48_m_axi_gmem_AWREGION,
	qsort_48_m_axi_gmem_AWUSER,
	qsort_48_m_axi_gmem_WREADY,
	qsort_48_m_axi_gmem_WVALID,
	qsort_48_m_axi_gmem_WDATA,
	qsort_48_m_axi_gmem_WSTRB,
	qsort_48_m_axi_gmem_WLAST,
	qsort_48_m_axi_gmem_WUSER,
	qsort_48_m_axi_gmem_BREADY,
	qsort_48_m_axi_gmem_BVALID,
	qsort_48_m_axi_gmem_BID,
	qsort_48_m_axi_gmem_BRESP,
	qsort_48_m_axi_gmem_BUSER,
	qsort_48_s_axi_control_ARREADY,
	qsort_48_s_axi_control_ARVALID,
	qsort_48_s_axi_control_ARADDR,
	qsort_48_s_axi_control_RREADY,
	qsort_48_s_axi_control_RVALID,
	qsort_48_s_axi_control_RDATA,
	qsort_48_s_axi_control_RRESP,
	qsort_48_s_axi_control_AWREADY,
	qsort_48_s_axi_control_AWVALID,
	qsort_48_s_axi_control_AWADDR,
	qsort_48_s_axi_control_WREADY,
	qsort_48_s_axi_control_WVALID,
	qsort_48_s_axi_control_WDATA,
	qsort_48_s_axi_control_WSTRB,
	qsort_48_s_axi_control_BREADY,
	qsort_48_s_axi_control_BVALID,
	qsort_48_s_axi_control_BRESP,
	qsort_49_m_axi_gmem_ARREADY,
	qsort_49_m_axi_gmem_ARVALID,
	qsort_49_m_axi_gmem_ARID,
	qsort_49_m_axi_gmem_ARADDR,
	qsort_49_m_axi_gmem_ARLEN,
	qsort_49_m_axi_gmem_ARSIZE,
	qsort_49_m_axi_gmem_ARBURST,
	qsort_49_m_axi_gmem_ARLOCK,
	qsort_49_m_axi_gmem_ARCACHE,
	qsort_49_m_axi_gmem_ARPROT,
	qsort_49_m_axi_gmem_ARQOS,
	qsort_49_m_axi_gmem_ARREGION,
	qsort_49_m_axi_gmem_ARUSER,
	qsort_49_m_axi_gmem_RREADY,
	qsort_49_m_axi_gmem_RVALID,
	qsort_49_m_axi_gmem_RID,
	qsort_49_m_axi_gmem_RDATA,
	qsort_49_m_axi_gmem_RRESP,
	qsort_49_m_axi_gmem_RLAST,
	qsort_49_m_axi_gmem_RUSER,
	qsort_49_m_axi_gmem_AWREADY,
	qsort_49_m_axi_gmem_AWVALID,
	qsort_49_m_axi_gmem_AWID,
	qsort_49_m_axi_gmem_AWADDR,
	qsort_49_m_axi_gmem_AWLEN,
	qsort_49_m_axi_gmem_AWSIZE,
	qsort_49_m_axi_gmem_AWBURST,
	qsort_49_m_axi_gmem_AWLOCK,
	qsort_49_m_axi_gmem_AWCACHE,
	qsort_49_m_axi_gmem_AWPROT,
	qsort_49_m_axi_gmem_AWQOS,
	qsort_49_m_axi_gmem_AWREGION,
	qsort_49_m_axi_gmem_AWUSER,
	qsort_49_m_axi_gmem_WREADY,
	qsort_49_m_axi_gmem_WVALID,
	qsort_49_m_axi_gmem_WDATA,
	qsort_49_m_axi_gmem_WSTRB,
	qsort_49_m_axi_gmem_WLAST,
	qsort_49_m_axi_gmem_WUSER,
	qsort_49_m_axi_gmem_BREADY,
	qsort_49_m_axi_gmem_BVALID,
	qsort_49_m_axi_gmem_BID,
	qsort_49_m_axi_gmem_BRESP,
	qsort_49_m_axi_gmem_BUSER,
	qsort_49_s_axi_control_ARREADY,
	qsort_49_s_axi_control_ARVALID,
	qsort_49_s_axi_control_ARADDR,
	qsort_49_s_axi_control_RREADY,
	qsort_49_s_axi_control_RVALID,
	qsort_49_s_axi_control_RDATA,
	qsort_49_s_axi_control_RRESP,
	qsort_49_s_axi_control_AWREADY,
	qsort_49_s_axi_control_AWVALID,
	qsort_49_s_axi_control_AWADDR,
	qsort_49_s_axi_control_WREADY,
	qsort_49_s_axi_control_WVALID,
	qsort_49_s_axi_control_WDATA,
	qsort_49_s_axi_control_WSTRB,
	qsort_49_s_axi_control_BREADY,
	qsort_49_s_axi_control_BVALID,
	qsort_49_s_axi_control_BRESP,
	qsort_50_m_axi_gmem_ARREADY,
	qsort_50_m_axi_gmem_ARVALID,
	qsort_50_m_axi_gmem_ARID,
	qsort_50_m_axi_gmem_ARADDR,
	qsort_50_m_axi_gmem_ARLEN,
	qsort_50_m_axi_gmem_ARSIZE,
	qsort_50_m_axi_gmem_ARBURST,
	qsort_50_m_axi_gmem_ARLOCK,
	qsort_50_m_axi_gmem_ARCACHE,
	qsort_50_m_axi_gmem_ARPROT,
	qsort_50_m_axi_gmem_ARQOS,
	qsort_50_m_axi_gmem_ARREGION,
	qsort_50_m_axi_gmem_ARUSER,
	qsort_50_m_axi_gmem_RREADY,
	qsort_50_m_axi_gmem_RVALID,
	qsort_50_m_axi_gmem_RID,
	qsort_50_m_axi_gmem_RDATA,
	qsort_50_m_axi_gmem_RRESP,
	qsort_50_m_axi_gmem_RLAST,
	qsort_50_m_axi_gmem_RUSER,
	qsort_50_m_axi_gmem_AWREADY,
	qsort_50_m_axi_gmem_AWVALID,
	qsort_50_m_axi_gmem_AWID,
	qsort_50_m_axi_gmem_AWADDR,
	qsort_50_m_axi_gmem_AWLEN,
	qsort_50_m_axi_gmem_AWSIZE,
	qsort_50_m_axi_gmem_AWBURST,
	qsort_50_m_axi_gmem_AWLOCK,
	qsort_50_m_axi_gmem_AWCACHE,
	qsort_50_m_axi_gmem_AWPROT,
	qsort_50_m_axi_gmem_AWQOS,
	qsort_50_m_axi_gmem_AWREGION,
	qsort_50_m_axi_gmem_AWUSER,
	qsort_50_m_axi_gmem_WREADY,
	qsort_50_m_axi_gmem_WVALID,
	qsort_50_m_axi_gmem_WDATA,
	qsort_50_m_axi_gmem_WSTRB,
	qsort_50_m_axi_gmem_WLAST,
	qsort_50_m_axi_gmem_WUSER,
	qsort_50_m_axi_gmem_BREADY,
	qsort_50_m_axi_gmem_BVALID,
	qsort_50_m_axi_gmem_BID,
	qsort_50_m_axi_gmem_BRESP,
	qsort_50_m_axi_gmem_BUSER,
	qsort_50_s_axi_control_ARREADY,
	qsort_50_s_axi_control_ARVALID,
	qsort_50_s_axi_control_ARADDR,
	qsort_50_s_axi_control_RREADY,
	qsort_50_s_axi_control_RVALID,
	qsort_50_s_axi_control_RDATA,
	qsort_50_s_axi_control_RRESP,
	qsort_50_s_axi_control_AWREADY,
	qsort_50_s_axi_control_AWVALID,
	qsort_50_s_axi_control_AWADDR,
	qsort_50_s_axi_control_WREADY,
	qsort_50_s_axi_control_WVALID,
	qsort_50_s_axi_control_WDATA,
	qsort_50_s_axi_control_WSTRB,
	qsort_50_s_axi_control_BREADY,
	qsort_50_s_axi_control_BVALID,
	qsort_50_s_axi_control_BRESP,
	qsort_51_m_axi_gmem_ARREADY,
	qsort_51_m_axi_gmem_ARVALID,
	qsort_51_m_axi_gmem_ARID,
	qsort_51_m_axi_gmem_ARADDR,
	qsort_51_m_axi_gmem_ARLEN,
	qsort_51_m_axi_gmem_ARSIZE,
	qsort_51_m_axi_gmem_ARBURST,
	qsort_51_m_axi_gmem_ARLOCK,
	qsort_51_m_axi_gmem_ARCACHE,
	qsort_51_m_axi_gmem_ARPROT,
	qsort_51_m_axi_gmem_ARQOS,
	qsort_51_m_axi_gmem_ARREGION,
	qsort_51_m_axi_gmem_ARUSER,
	qsort_51_m_axi_gmem_RREADY,
	qsort_51_m_axi_gmem_RVALID,
	qsort_51_m_axi_gmem_RID,
	qsort_51_m_axi_gmem_RDATA,
	qsort_51_m_axi_gmem_RRESP,
	qsort_51_m_axi_gmem_RLAST,
	qsort_51_m_axi_gmem_RUSER,
	qsort_51_m_axi_gmem_AWREADY,
	qsort_51_m_axi_gmem_AWVALID,
	qsort_51_m_axi_gmem_AWID,
	qsort_51_m_axi_gmem_AWADDR,
	qsort_51_m_axi_gmem_AWLEN,
	qsort_51_m_axi_gmem_AWSIZE,
	qsort_51_m_axi_gmem_AWBURST,
	qsort_51_m_axi_gmem_AWLOCK,
	qsort_51_m_axi_gmem_AWCACHE,
	qsort_51_m_axi_gmem_AWPROT,
	qsort_51_m_axi_gmem_AWQOS,
	qsort_51_m_axi_gmem_AWREGION,
	qsort_51_m_axi_gmem_AWUSER,
	qsort_51_m_axi_gmem_WREADY,
	qsort_51_m_axi_gmem_WVALID,
	qsort_51_m_axi_gmem_WDATA,
	qsort_51_m_axi_gmem_WSTRB,
	qsort_51_m_axi_gmem_WLAST,
	qsort_51_m_axi_gmem_WUSER,
	qsort_51_m_axi_gmem_BREADY,
	qsort_51_m_axi_gmem_BVALID,
	qsort_51_m_axi_gmem_BID,
	qsort_51_m_axi_gmem_BRESP,
	qsort_51_m_axi_gmem_BUSER,
	qsort_51_s_axi_control_ARREADY,
	qsort_51_s_axi_control_ARVALID,
	qsort_51_s_axi_control_ARADDR,
	qsort_51_s_axi_control_RREADY,
	qsort_51_s_axi_control_RVALID,
	qsort_51_s_axi_control_RDATA,
	qsort_51_s_axi_control_RRESP,
	qsort_51_s_axi_control_AWREADY,
	qsort_51_s_axi_control_AWVALID,
	qsort_51_s_axi_control_AWADDR,
	qsort_51_s_axi_control_WREADY,
	qsort_51_s_axi_control_WVALID,
	qsort_51_s_axi_control_WDATA,
	qsort_51_s_axi_control_WSTRB,
	qsort_51_s_axi_control_BREADY,
	qsort_51_s_axi_control_BVALID,
	qsort_51_s_axi_control_BRESP,
	qsort_52_m_axi_gmem_ARREADY,
	qsort_52_m_axi_gmem_ARVALID,
	qsort_52_m_axi_gmem_ARID,
	qsort_52_m_axi_gmem_ARADDR,
	qsort_52_m_axi_gmem_ARLEN,
	qsort_52_m_axi_gmem_ARSIZE,
	qsort_52_m_axi_gmem_ARBURST,
	qsort_52_m_axi_gmem_ARLOCK,
	qsort_52_m_axi_gmem_ARCACHE,
	qsort_52_m_axi_gmem_ARPROT,
	qsort_52_m_axi_gmem_ARQOS,
	qsort_52_m_axi_gmem_ARREGION,
	qsort_52_m_axi_gmem_ARUSER,
	qsort_52_m_axi_gmem_RREADY,
	qsort_52_m_axi_gmem_RVALID,
	qsort_52_m_axi_gmem_RID,
	qsort_52_m_axi_gmem_RDATA,
	qsort_52_m_axi_gmem_RRESP,
	qsort_52_m_axi_gmem_RLAST,
	qsort_52_m_axi_gmem_RUSER,
	qsort_52_m_axi_gmem_AWREADY,
	qsort_52_m_axi_gmem_AWVALID,
	qsort_52_m_axi_gmem_AWID,
	qsort_52_m_axi_gmem_AWADDR,
	qsort_52_m_axi_gmem_AWLEN,
	qsort_52_m_axi_gmem_AWSIZE,
	qsort_52_m_axi_gmem_AWBURST,
	qsort_52_m_axi_gmem_AWLOCK,
	qsort_52_m_axi_gmem_AWCACHE,
	qsort_52_m_axi_gmem_AWPROT,
	qsort_52_m_axi_gmem_AWQOS,
	qsort_52_m_axi_gmem_AWREGION,
	qsort_52_m_axi_gmem_AWUSER,
	qsort_52_m_axi_gmem_WREADY,
	qsort_52_m_axi_gmem_WVALID,
	qsort_52_m_axi_gmem_WDATA,
	qsort_52_m_axi_gmem_WSTRB,
	qsort_52_m_axi_gmem_WLAST,
	qsort_52_m_axi_gmem_WUSER,
	qsort_52_m_axi_gmem_BREADY,
	qsort_52_m_axi_gmem_BVALID,
	qsort_52_m_axi_gmem_BID,
	qsort_52_m_axi_gmem_BRESP,
	qsort_52_m_axi_gmem_BUSER,
	qsort_52_s_axi_control_ARREADY,
	qsort_52_s_axi_control_ARVALID,
	qsort_52_s_axi_control_ARADDR,
	qsort_52_s_axi_control_RREADY,
	qsort_52_s_axi_control_RVALID,
	qsort_52_s_axi_control_RDATA,
	qsort_52_s_axi_control_RRESP,
	qsort_52_s_axi_control_AWREADY,
	qsort_52_s_axi_control_AWVALID,
	qsort_52_s_axi_control_AWADDR,
	qsort_52_s_axi_control_WREADY,
	qsort_52_s_axi_control_WVALID,
	qsort_52_s_axi_control_WDATA,
	qsort_52_s_axi_control_WSTRB,
	qsort_52_s_axi_control_BREADY,
	qsort_52_s_axi_control_BVALID,
	qsort_52_s_axi_control_BRESP,
	qsort_53_m_axi_gmem_ARREADY,
	qsort_53_m_axi_gmem_ARVALID,
	qsort_53_m_axi_gmem_ARID,
	qsort_53_m_axi_gmem_ARADDR,
	qsort_53_m_axi_gmem_ARLEN,
	qsort_53_m_axi_gmem_ARSIZE,
	qsort_53_m_axi_gmem_ARBURST,
	qsort_53_m_axi_gmem_ARLOCK,
	qsort_53_m_axi_gmem_ARCACHE,
	qsort_53_m_axi_gmem_ARPROT,
	qsort_53_m_axi_gmem_ARQOS,
	qsort_53_m_axi_gmem_ARREGION,
	qsort_53_m_axi_gmem_ARUSER,
	qsort_53_m_axi_gmem_RREADY,
	qsort_53_m_axi_gmem_RVALID,
	qsort_53_m_axi_gmem_RID,
	qsort_53_m_axi_gmem_RDATA,
	qsort_53_m_axi_gmem_RRESP,
	qsort_53_m_axi_gmem_RLAST,
	qsort_53_m_axi_gmem_RUSER,
	qsort_53_m_axi_gmem_AWREADY,
	qsort_53_m_axi_gmem_AWVALID,
	qsort_53_m_axi_gmem_AWID,
	qsort_53_m_axi_gmem_AWADDR,
	qsort_53_m_axi_gmem_AWLEN,
	qsort_53_m_axi_gmem_AWSIZE,
	qsort_53_m_axi_gmem_AWBURST,
	qsort_53_m_axi_gmem_AWLOCK,
	qsort_53_m_axi_gmem_AWCACHE,
	qsort_53_m_axi_gmem_AWPROT,
	qsort_53_m_axi_gmem_AWQOS,
	qsort_53_m_axi_gmem_AWREGION,
	qsort_53_m_axi_gmem_AWUSER,
	qsort_53_m_axi_gmem_WREADY,
	qsort_53_m_axi_gmem_WVALID,
	qsort_53_m_axi_gmem_WDATA,
	qsort_53_m_axi_gmem_WSTRB,
	qsort_53_m_axi_gmem_WLAST,
	qsort_53_m_axi_gmem_WUSER,
	qsort_53_m_axi_gmem_BREADY,
	qsort_53_m_axi_gmem_BVALID,
	qsort_53_m_axi_gmem_BID,
	qsort_53_m_axi_gmem_BRESP,
	qsort_53_m_axi_gmem_BUSER,
	qsort_53_s_axi_control_ARREADY,
	qsort_53_s_axi_control_ARVALID,
	qsort_53_s_axi_control_ARADDR,
	qsort_53_s_axi_control_RREADY,
	qsort_53_s_axi_control_RVALID,
	qsort_53_s_axi_control_RDATA,
	qsort_53_s_axi_control_RRESP,
	qsort_53_s_axi_control_AWREADY,
	qsort_53_s_axi_control_AWVALID,
	qsort_53_s_axi_control_AWADDR,
	qsort_53_s_axi_control_WREADY,
	qsort_53_s_axi_control_WVALID,
	qsort_53_s_axi_control_WDATA,
	qsort_53_s_axi_control_WSTRB,
	qsort_53_s_axi_control_BREADY,
	qsort_53_s_axi_control_BVALID,
	qsort_53_s_axi_control_BRESP,
	qsort_54_m_axi_gmem_ARREADY,
	qsort_54_m_axi_gmem_ARVALID,
	qsort_54_m_axi_gmem_ARID,
	qsort_54_m_axi_gmem_ARADDR,
	qsort_54_m_axi_gmem_ARLEN,
	qsort_54_m_axi_gmem_ARSIZE,
	qsort_54_m_axi_gmem_ARBURST,
	qsort_54_m_axi_gmem_ARLOCK,
	qsort_54_m_axi_gmem_ARCACHE,
	qsort_54_m_axi_gmem_ARPROT,
	qsort_54_m_axi_gmem_ARQOS,
	qsort_54_m_axi_gmem_ARREGION,
	qsort_54_m_axi_gmem_ARUSER,
	qsort_54_m_axi_gmem_RREADY,
	qsort_54_m_axi_gmem_RVALID,
	qsort_54_m_axi_gmem_RID,
	qsort_54_m_axi_gmem_RDATA,
	qsort_54_m_axi_gmem_RRESP,
	qsort_54_m_axi_gmem_RLAST,
	qsort_54_m_axi_gmem_RUSER,
	qsort_54_m_axi_gmem_AWREADY,
	qsort_54_m_axi_gmem_AWVALID,
	qsort_54_m_axi_gmem_AWID,
	qsort_54_m_axi_gmem_AWADDR,
	qsort_54_m_axi_gmem_AWLEN,
	qsort_54_m_axi_gmem_AWSIZE,
	qsort_54_m_axi_gmem_AWBURST,
	qsort_54_m_axi_gmem_AWLOCK,
	qsort_54_m_axi_gmem_AWCACHE,
	qsort_54_m_axi_gmem_AWPROT,
	qsort_54_m_axi_gmem_AWQOS,
	qsort_54_m_axi_gmem_AWREGION,
	qsort_54_m_axi_gmem_AWUSER,
	qsort_54_m_axi_gmem_WREADY,
	qsort_54_m_axi_gmem_WVALID,
	qsort_54_m_axi_gmem_WDATA,
	qsort_54_m_axi_gmem_WSTRB,
	qsort_54_m_axi_gmem_WLAST,
	qsort_54_m_axi_gmem_WUSER,
	qsort_54_m_axi_gmem_BREADY,
	qsort_54_m_axi_gmem_BVALID,
	qsort_54_m_axi_gmem_BID,
	qsort_54_m_axi_gmem_BRESP,
	qsort_54_m_axi_gmem_BUSER,
	qsort_54_s_axi_control_ARREADY,
	qsort_54_s_axi_control_ARVALID,
	qsort_54_s_axi_control_ARADDR,
	qsort_54_s_axi_control_RREADY,
	qsort_54_s_axi_control_RVALID,
	qsort_54_s_axi_control_RDATA,
	qsort_54_s_axi_control_RRESP,
	qsort_54_s_axi_control_AWREADY,
	qsort_54_s_axi_control_AWVALID,
	qsort_54_s_axi_control_AWADDR,
	qsort_54_s_axi_control_WREADY,
	qsort_54_s_axi_control_WVALID,
	qsort_54_s_axi_control_WDATA,
	qsort_54_s_axi_control_WSTRB,
	qsort_54_s_axi_control_BREADY,
	qsort_54_s_axi_control_BVALID,
	qsort_54_s_axi_control_BRESP,
	qsort_55_m_axi_gmem_ARREADY,
	qsort_55_m_axi_gmem_ARVALID,
	qsort_55_m_axi_gmem_ARID,
	qsort_55_m_axi_gmem_ARADDR,
	qsort_55_m_axi_gmem_ARLEN,
	qsort_55_m_axi_gmem_ARSIZE,
	qsort_55_m_axi_gmem_ARBURST,
	qsort_55_m_axi_gmem_ARLOCK,
	qsort_55_m_axi_gmem_ARCACHE,
	qsort_55_m_axi_gmem_ARPROT,
	qsort_55_m_axi_gmem_ARQOS,
	qsort_55_m_axi_gmem_ARREGION,
	qsort_55_m_axi_gmem_ARUSER,
	qsort_55_m_axi_gmem_RREADY,
	qsort_55_m_axi_gmem_RVALID,
	qsort_55_m_axi_gmem_RID,
	qsort_55_m_axi_gmem_RDATA,
	qsort_55_m_axi_gmem_RRESP,
	qsort_55_m_axi_gmem_RLAST,
	qsort_55_m_axi_gmem_RUSER,
	qsort_55_m_axi_gmem_AWREADY,
	qsort_55_m_axi_gmem_AWVALID,
	qsort_55_m_axi_gmem_AWID,
	qsort_55_m_axi_gmem_AWADDR,
	qsort_55_m_axi_gmem_AWLEN,
	qsort_55_m_axi_gmem_AWSIZE,
	qsort_55_m_axi_gmem_AWBURST,
	qsort_55_m_axi_gmem_AWLOCK,
	qsort_55_m_axi_gmem_AWCACHE,
	qsort_55_m_axi_gmem_AWPROT,
	qsort_55_m_axi_gmem_AWQOS,
	qsort_55_m_axi_gmem_AWREGION,
	qsort_55_m_axi_gmem_AWUSER,
	qsort_55_m_axi_gmem_WREADY,
	qsort_55_m_axi_gmem_WVALID,
	qsort_55_m_axi_gmem_WDATA,
	qsort_55_m_axi_gmem_WSTRB,
	qsort_55_m_axi_gmem_WLAST,
	qsort_55_m_axi_gmem_WUSER,
	qsort_55_m_axi_gmem_BREADY,
	qsort_55_m_axi_gmem_BVALID,
	qsort_55_m_axi_gmem_BID,
	qsort_55_m_axi_gmem_BRESP,
	qsort_55_m_axi_gmem_BUSER,
	qsort_55_s_axi_control_ARREADY,
	qsort_55_s_axi_control_ARVALID,
	qsort_55_s_axi_control_ARADDR,
	qsort_55_s_axi_control_RREADY,
	qsort_55_s_axi_control_RVALID,
	qsort_55_s_axi_control_RDATA,
	qsort_55_s_axi_control_RRESP,
	qsort_55_s_axi_control_AWREADY,
	qsort_55_s_axi_control_AWVALID,
	qsort_55_s_axi_control_AWADDR,
	qsort_55_s_axi_control_WREADY,
	qsort_55_s_axi_control_WVALID,
	qsort_55_s_axi_control_WDATA,
	qsort_55_s_axi_control_WSTRB,
	qsort_55_s_axi_control_BREADY,
	qsort_55_s_axi_control_BVALID,
	qsort_55_s_axi_control_BRESP,
	qsort_56_m_axi_gmem_ARREADY,
	qsort_56_m_axi_gmem_ARVALID,
	qsort_56_m_axi_gmem_ARID,
	qsort_56_m_axi_gmem_ARADDR,
	qsort_56_m_axi_gmem_ARLEN,
	qsort_56_m_axi_gmem_ARSIZE,
	qsort_56_m_axi_gmem_ARBURST,
	qsort_56_m_axi_gmem_ARLOCK,
	qsort_56_m_axi_gmem_ARCACHE,
	qsort_56_m_axi_gmem_ARPROT,
	qsort_56_m_axi_gmem_ARQOS,
	qsort_56_m_axi_gmem_ARREGION,
	qsort_56_m_axi_gmem_ARUSER,
	qsort_56_m_axi_gmem_RREADY,
	qsort_56_m_axi_gmem_RVALID,
	qsort_56_m_axi_gmem_RID,
	qsort_56_m_axi_gmem_RDATA,
	qsort_56_m_axi_gmem_RRESP,
	qsort_56_m_axi_gmem_RLAST,
	qsort_56_m_axi_gmem_RUSER,
	qsort_56_m_axi_gmem_AWREADY,
	qsort_56_m_axi_gmem_AWVALID,
	qsort_56_m_axi_gmem_AWID,
	qsort_56_m_axi_gmem_AWADDR,
	qsort_56_m_axi_gmem_AWLEN,
	qsort_56_m_axi_gmem_AWSIZE,
	qsort_56_m_axi_gmem_AWBURST,
	qsort_56_m_axi_gmem_AWLOCK,
	qsort_56_m_axi_gmem_AWCACHE,
	qsort_56_m_axi_gmem_AWPROT,
	qsort_56_m_axi_gmem_AWQOS,
	qsort_56_m_axi_gmem_AWREGION,
	qsort_56_m_axi_gmem_AWUSER,
	qsort_56_m_axi_gmem_WREADY,
	qsort_56_m_axi_gmem_WVALID,
	qsort_56_m_axi_gmem_WDATA,
	qsort_56_m_axi_gmem_WSTRB,
	qsort_56_m_axi_gmem_WLAST,
	qsort_56_m_axi_gmem_WUSER,
	qsort_56_m_axi_gmem_BREADY,
	qsort_56_m_axi_gmem_BVALID,
	qsort_56_m_axi_gmem_BID,
	qsort_56_m_axi_gmem_BRESP,
	qsort_56_m_axi_gmem_BUSER,
	qsort_56_s_axi_control_ARREADY,
	qsort_56_s_axi_control_ARVALID,
	qsort_56_s_axi_control_ARADDR,
	qsort_56_s_axi_control_RREADY,
	qsort_56_s_axi_control_RVALID,
	qsort_56_s_axi_control_RDATA,
	qsort_56_s_axi_control_RRESP,
	qsort_56_s_axi_control_AWREADY,
	qsort_56_s_axi_control_AWVALID,
	qsort_56_s_axi_control_AWADDR,
	qsort_56_s_axi_control_WREADY,
	qsort_56_s_axi_control_WVALID,
	qsort_56_s_axi_control_WDATA,
	qsort_56_s_axi_control_WSTRB,
	qsort_56_s_axi_control_BREADY,
	qsort_56_s_axi_control_BVALID,
	qsort_56_s_axi_control_BRESP,
	qsort_57_m_axi_gmem_ARREADY,
	qsort_57_m_axi_gmem_ARVALID,
	qsort_57_m_axi_gmem_ARID,
	qsort_57_m_axi_gmem_ARADDR,
	qsort_57_m_axi_gmem_ARLEN,
	qsort_57_m_axi_gmem_ARSIZE,
	qsort_57_m_axi_gmem_ARBURST,
	qsort_57_m_axi_gmem_ARLOCK,
	qsort_57_m_axi_gmem_ARCACHE,
	qsort_57_m_axi_gmem_ARPROT,
	qsort_57_m_axi_gmem_ARQOS,
	qsort_57_m_axi_gmem_ARREGION,
	qsort_57_m_axi_gmem_ARUSER,
	qsort_57_m_axi_gmem_RREADY,
	qsort_57_m_axi_gmem_RVALID,
	qsort_57_m_axi_gmem_RID,
	qsort_57_m_axi_gmem_RDATA,
	qsort_57_m_axi_gmem_RRESP,
	qsort_57_m_axi_gmem_RLAST,
	qsort_57_m_axi_gmem_RUSER,
	qsort_57_m_axi_gmem_AWREADY,
	qsort_57_m_axi_gmem_AWVALID,
	qsort_57_m_axi_gmem_AWID,
	qsort_57_m_axi_gmem_AWADDR,
	qsort_57_m_axi_gmem_AWLEN,
	qsort_57_m_axi_gmem_AWSIZE,
	qsort_57_m_axi_gmem_AWBURST,
	qsort_57_m_axi_gmem_AWLOCK,
	qsort_57_m_axi_gmem_AWCACHE,
	qsort_57_m_axi_gmem_AWPROT,
	qsort_57_m_axi_gmem_AWQOS,
	qsort_57_m_axi_gmem_AWREGION,
	qsort_57_m_axi_gmem_AWUSER,
	qsort_57_m_axi_gmem_WREADY,
	qsort_57_m_axi_gmem_WVALID,
	qsort_57_m_axi_gmem_WDATA,
	qsort_57_m_axi_gmem_WSTRB,
	qsort_57_m_axi_gmem_WLAST,
	qsort_57_m_axi_gmem_WUSER,
	qsort_57_m_axi_gmem_BREADY,
	qsort_57_m_axi_gmem_BVALID,
	qsort_57_m_axi_gmem_BID,
	qsort_57_m_axi_gmem_BRESP,
	qsort_57_m_axi_gmem_BUSER,
	qsort_57_s_axi_control_ARREADY,
	qsort_57_s_axi_control_ARVALID,
	qsort_57_s_axi_control_ARADDR,
	qsort_57_s_axi_control_RREADY,
	qsort_57_s_axi_control_RVALID,
	qsort_57_s_axi_control_RDATA,
	qsort_57_s_axi_control_RRESP,
	qsort_57_s_axi_control_AWREADY,
	qsort_57_s_axi_control_AWVALID,
	qsort_57_s_axi_control_AWADDR,
	qsort_57_s_axi_control_WREADY,
	qsort_57_s_axi_control_WVALID,
	qsort_57_s_axi_control_WDATA,
	qsort_57_s_axi_control_WSTRB,
	qsort_57_s_axi_control_BREADY,
	qsort_57_s_axi_control_BVALID,
	qsort_57_s_axi_control_BRESP,
	qsort_58_m_axi_gmem_ARREADY,
	qsort_58_m_axi_gmem_ARVALID,
	qsort_58_m_axi_gmem_ARID,
	qsort_58_m_axi_gmem_ARADDR,
	qsort_58_m_axi_gmem_ARLEN,
	qsort_58_m_axi_gmem_ARSIZE,
	qsort_58_m_axi_gmem_ARBURST,
	qsort_58_m_axi_gmem_ARLOCK,
	qsort_58_m_axi_gmem_ARCACHE,
	qsort_58_m_axi_gmem_ARPROT,
	qsort_58_m_axi_gmem_ARQOS,
	qsort_58_m_axi_gmem_ARREGION,
	qsort_58_m_axi_gmem_ARUSER,
	qsort_58_m_axi_gmem_RREADY,
	qsort_58_m_axi_gmem_RVALID,
	qsort_58_m_axi_gmem_RID,
	qsort_58_m_axi_gmem_RDATA,
	qsort_58_m_axi_gmem_RRESP,
	qsort_58_m_axi_gmem_RLAST,
	qsort_58_m_axi_gmem_RUSER,
	qsort_58_m_axi_gmem_AWREADY,
	qsort_58_m_axi_gmem_AWVALID,
	qsort_58_m_axi_gmem_AWID,
	qsort_58_m_axi_gmem_AWADDR,
	qsort_58_m_axi_gmem_AWLEN,
	qsort_58_m_axi_gmem_AWSIZE,
	qsort_58_m_axi_gmem_AWBURST,
	qsort_58_m_axi_gmem_AWLOCK,
	qsort_58_m_axi_gmem_AWCACHE,
	qsort_58_m_axi_gmem_AWPROT,
	qsort_58_m_axi_gmem_AWQOS,
	qsort_58_m_axi_gmem_AWREGION,
	qsort_58_m_axi_gmem_AWUSER,
	qsort_58_m_axi_gmem_WREADY,
	qsort_58_m_axi_gmem_WVALID,
	qsort_58_m_axi_gmem_WDATA,
	qsort_58_m_axi_gmem_WSTRB,
	qsort_58_m_axi_gmem_WLAST,
	qsort_58_m_axi_gmem_WUSER,
	qsort_58_m_axi_gmem_BREADY,
	qsort_58_m_axi_gmem_BVALID,
	qsort_58_m_axi_gmem_BID,
	qsort_58_m_axi_gmem_BRESP,
	qsort_58_m_axi_gmem_BUSER,
	qsort_58_s_axi_control_ARREADY,
	qsort_58_s_axi_control_ARVALID,
	qsort_58_s_axi_control_ARADDR,
	qsort_58_s_axi_control_RREADY,
	qsort_58_s_axi_control_RVALID,
	qsort_58_s_axi_control_RDATA,
	qsort_58_s_axi_control_RRESP,
	qsort_58_s_axi_control_AWREADY,
	qsort_58_s_axi_control_AWVALID,
	qsort_58_s_axi_control_AWADDR,
	qsort_58_s_axi_control_WREADY,
	qsort_58_s_axi_control_WVALID,
	qsort_58_s_axi_control_WDATA,
	qsort_58_s_axi_control_WSTRB,
	qsort_58_s_axi_control_BREADY,
	qsort_58_s_axi_control_BVALID,
	qsort_58_s_axi_control_BRESP,
	qsort_59_m_axi_gmem_ARREADY,
	qsort_59_m_axi_gmem_ARVALID,
	qsort_59_m_axi_gmem_ARID,
	qsort_59_m_axi_gmem_ARADDR,
	qsort_59_m_axi_gmem_ARLEN,
	qsort_59_m_axi_gmem_ARSIZE,
	qsort_59_m_axi_gmem_ARBURST,
	qsort_59_m_axi_gmem_ARLOCK,
	qsort_59_m_axi_gmem_ARCACHE,
	qsort_59_m_axi_gmem_ARPROT,
	qsort_59_m_axi_gmem_ARQOS,
	qsort_59_m_axi_gmem_ARREGION,
	qsort_59_m_axi_gmem_ARUSER,
	qsort_59_m_axi_gmem_RREADY,
	qsort_59_m_axi_gmem_RVALID,
	qsort_59_m_axi_gmem_RID,
	qsort_59_m_axi_gmem_RDATA,
	qsort_59_m_axi_gmem_RRESP,
	qsort_59_m_axi_gmem_RLAST,
	qsort_59_m_axi_gmem_RUSER,
	qsort_59_m_axi_gmem_AWREADY,
	qsort_59_m_axi_gmem_AWVALID,
	qsort_59_m_axi_gmem_AWID,
	qsort_59_m_axi_gmem_AWADDR,
	qsort_59_m_axi_gmem_AWLEN,
	qsort_59_m_axi_gmem_AWSIZE,
	qsort_59_m_axi_gmem_AWBURST,
	qsort_59_m_axi_gmem_AWLOCK,
	qsort_59_m_axi_gmem_AWCACHE,
	qsort_59_m_axi_gmem_AWPROT,
	qsort_59_m_axi_gmem_AWQOS,
	qsort_59_m_axi_gmem_AWREGION,
	qsort_59_m_axi_gmem_AWUSER,
	qsort_59_m_axi_gmem_WREADY,
	qsort_59_m_axi_gmem_WVALID,
	qsort_59_m_axi_gmem_WDATA,
	qsort_59_m_axi_gmem_WSTRB,
	qsort_59_m_axi_gmem_WLAST,
	qsort_59_m_axi_gmem_WUSER,
	qsort_59_m_axi_gmem_BREADY,
	qsort_59_m_axi_gmem_BVALID,
	qsort_59_m_axi_gmem_BID,
	qsort_59_m_axi_gmem_BRESP,
	qsort_59_m_axi_gmem_BUSER,
	qsort_59_s_axi_control_ARREADY,
	qsort_59_s_axi_control_ARVALID,
	qsort_59_s_axi_control_ARADDR,
	qsort_59_s_axi_control_RREADY,
	qsort_59_s_axi_control_RVALID,
	qsort_59_s_axi_control_RDATA,
	qsort_59_s_axi_control_RRESP,
	qsort_59_s_axi_control_AWREADY,
	qsort_59_s_axi_control_AWVALID,
	qsort_59_s_axi_control_AWADDR,
	qsort_59_s_axi_control_WREADY,
	qsort_59_s_axi_control_WVALID,
	qsort_59_s_axi_control_WDATA,
	qsort_59_s_axi_control_WSTRB,
	qsort_59_s_axi_control_BREADY,
	qsort_59_s_axi_control_BVALID,
	qsort_59_s_axi_control_BRESP,
	qsort_60_m_axi_gmem_ARREADY,
	qsort_60_m_axi_gmem_ARVALID,
	qsort_60_m_axi_gmem_ARID,
	qsort_60_m_axi_gmem_ARADDR,
	qsort_60_m_axi_gmem_ARLEN,
	qsort_60_m_axi_gmem_ARSIZE,
	qsort_60_m_axi_gmem_ARBURST,
	qsort_60_m_axi_gmem_ARLOCK,
	qsort_60_m_axi_gmem_ARCACHE,
	qsort_60_m_axi_gmem_ARPROT,
	qsort_60_m_axi_gmem_ARQOS,
	qsort_60_m_axi_gmem_ARREGION,
	qsort_60_m_axi_gmem_ARUSER,
	qsort_60_m_axi_gmem_RREADY,
	qsort_60_m_axi_gmem_RVALID,
	qsort_60_m_axi_gmem_RID,
	qsort_60_m_axi_gmem_RDATA,
	qsort_60_m_axi_gmem_RRESP,
	qsort_60_m_axi_gmem_RLAST,
	qsort_60_m_axi_gmem_RUSER,
	qsort_60_m_axi_gmem_AWREADY,
	qsort_60_m_axi_gmem_AWVALID,
	qsort_60_m_axi_gmem_AWID,
	qsort_60_m_axi_gmem_AWADDR,
	qsort_60_m_axi_gmem_AWLEN,
	qsort_60_m_axi_gmem_AWSIZE,
	qsort_60_m_axi_gmem_AWBURST,
	qsort_60_m_axi_gmem_AWLOCK,
	qsort_60_m_axi_gmem_AWCACHE,
	qsort_60_m_axi_gmem_AWPROT,
	qsort_60_m_axi_gmem_AWQOS,
	qsort_60_m_axi_gmem_AWREGION,
	qsort_60_m_axi_gmem_AWUSER,
	qsort_60_m_axi_gmem_WREADY,
	qsort_60_m_axi_gmem_WVALID,
	qsort_60_m_axi_gmem_WDATA,
	qsort_60_m_axi_gmem_WSTRB,
	qsort_60_m_axi_gmem_WLAST,
	qsort_60_m_axi_gmem_WUSER,
	qsort_60_m_axi_gmem_BREADY,
	qsort_60_m_axi_gmem_BVALID,
	qsort_60_m_axi_gmem_BID,
	qsort_60_m_axi_gmem_BRESP,
	qsort_60_m_axi_gmem_BUSER,
	qsort_60_s_axi_control_ARREADY,
	qsort_60_s_axi_control_ARVALID,
	qsort_60_s_axi_control_ARADDR,
	qsort_60_s_axi_control_RREADY,
	qsort_60_s_axi_control_RVALID,
	qsort_60_s_axi_control_RDATA,
	qsort_60_s_axi_control_RRESP,
	qsort_60_s_axi_control_AWREADY,
	qsort_60_s_axi_control_AWVALID,
	qsort_60_s_axi_control_AWADDR,
	qsort_60_s_axi_control_WREADY,
	qsort_60_s_axi_control_WVALID,
	qsort_60_s_axi_control_WDATA,
	qsort_60_s_axi_control_WSTRB,
	qsort_60_s_axi_control_BREADY,
	qsort_60_s_axi_control_BVALID,
	qsort_60_s_axi_control_BRESP,
	qsort_61_m_axi_gmem_ARREADY,
	qsort_61_m_axi_gmem_ARVALID,
	qsort_61_m_axi_gmem_ARID,
	qsort_61_m_axi_gmem_ARADDR,
	qsort_61_m_axi_gmem_ARLEN,
	qsort_61_m_axi_gmem_ARSIZE,
	qsort_61_m_axi_gmem_ARBURST,
	qsort_61_m_axi_gmem_ARLOCK,
	qsort_61_m_axi_gmem_ARCACHE,
	qsort_61_m_axi_gmem_ARPROT,
	qsort_61_m_axi_gmem_ARQOS,
	qsort_61_m_axi_gmem_ARREGION,
	qsort_61_m_axi_gmem_ARUSER,
	qsort_61_m_axi_gmem_RREADY,
	qsort_61_m_axi_gmem_RVALID,
	qsort_61_m_axi_gmem_RID,
	qsort_61_m_axi_gmem_RDATA,
	qsort_61_m_axi_gmem_RRESP,
	qsort_61_m_axi_gmem_RLAST,
	qsort_61_m_axi_gmem_RUSER,
	qsort_61_m_axi_gmem_AWREADY,
	qsort_61_m_axi_gmem_AWVALID,
	qsort_61_m_axi_gmem_AWID,
	qsort_61_m_axi_gmem_AWADDR,
	qsort_61_m_axi_gmem_AWLEN,
	qsort_61_m_axi_gmem_AWSIZE,
	qsort_61_m_axi_gmem_AWBURST,
	qsort_61_m_axi_gmem_AWLOCK,
	qsort_61_m_axi_gmem_AWCACHE,
	qsort_61_m_axi_gmem_AWPROT,
	qsort_61_m_axi_gmem_AWQOS,
	qsort_61_m_axi_gmem_AWREGION,
	qsort_61_m_axi_gmem_AWUSER,
	qsort_61_m_axi_gmem_WREADY,
	qsort_61_m_axi_gmem_WVALID,
	qsort_61_m_axi_gmem_WDATA,
	qsort_61_m_axi_gmem_WSTRB,
	qsort_61_m_axi_gmem_WLAST,
	qsort_61_m_axi_gmem_WUSER,
	qsort_61_m_axi_gmem_BREADY,
	qsort_61_m_axi_gmem_BVALID,
	qsort_61_m_axi_gmem_BID,
	qsort_61_m_axi_gmem_BRESP,
	qsort_61_m_axi_gmem_BUSER,
	qsort_61_s_axi_control_ARREADY,
	qsort_61_s_axi_control_ARVALID,
	qsort_61_s_axi_control_ARADDR,
	qsort_61_s_axi_control_RREADY,
	qsort_61_s_axi_control_RVALID,
	qsort_61_s_axi_control_RDATA,
	qsort_61_s_axi_control_RRESP,
	qsort_61_s_axi_control_AWREADY,
	qsort_61_s_axi_control_AWVALID,
	qsort_61_s_axi_control_AWADDR,
	qsort_61_s_axi_control_WREADY,
	qsort_61_s_axi_control_WVALID,
	qsort_61_s_axi_control_WDATA,
	qsort_61_s_axi_control_WSTRB,
	qsort_61_s_axi_control_BREADY,
	qsort_61_s_axi_control_BVALID,
	qsort_61_s_axi_control_BRESP,
	qsort_62_m_axi_gmem_ARREADY,
	qsort_62_m_axi_gmem_ARVALID,
	qsort_62_m_axi_gmem_ARID,
	qsort_62_m_axi_gmem_ARADDR,
	qsort_62_m_axi_gmem_ARLEN,
	qsort_62_m_axi_gmem_ARSIZE,
	qsort_62_m_axi_gmem_ARBURST,
	qsort_62_m_axi_gmem_ARLOCK,
	qsort_62_m_axi_gmem_ARCACHE,
	qsort_62_m_axi_gmem_ARPROT,
	qsort_62_m_axi_gmem_ARQOS,
	qsort_62_m_axi_gmem_ARREGION,
	qsort_62_m_axi_gmem_ARUSER,
	qsort_62_m_axi_gmem_RREADY,
	qsort_62_m_axi_gmem_RVALID,
	qsort_62_m_axi_gmem_RID,
	qsort_62_m_axi_gmem_RDATA,
	qsort_62_m_axi_gmem_RRESP,
	qsort_62_m_axi_gmem_RLAST,
	qsort_62_m_axi_gmem_RUSER,
	qsort_62_m_axi_gmem_AWREADY,
	qsort_62_m_axi_gmem_AWVALID,
	qsort_62_m_axi_gmem_AWID,
	qsort_62_m_axi_gmem_AWADDR,
	qsort_62_m_axi_gmem_AWLEN,
	qsort_62_m_axi_gmem_AWSIZE,
	qsort_62_m_axi_gmem_AWBURST,
	qsort_62_m_axi_gmem_AWLOCK,
	qsort_62_m_axi_gmem_AWCACHE,
	qsort_62_m_axi_gmem_AWPROT,
	qsort_62_m_axi_gmem_AWQOS,
	qsort_62_m_axi_gmem_AWREGION,
	qsort_62_m_axi_gmem_AWUSER,
	qsort_62_m_axi_gmem_WREADY,
	qsort_62_m_axi_gmem_WVALID,
	qsort_62_m_axi_gmem_WDATA,
	qsort_62_m_axi_gmem_WSTRB,
	qsort_62_m_axi_gmem_WLAST,
	qsort_62_m_axi_gmem_WUSER,
	qsort_62_m_axi_gmem_BREADY,
	qsort_62_m_axi_gmem_BVALID,
	qsort_62_m_axi_gmem_BID,
	qsort_62_m_axi_gmem_BRESP,
	qsort_62_m_axi_gmem_BUSER,
	qsort_62_s_axi_control_ARREADY,
	qsort_62_s_axi_control_ARVALID,
	qsort_62_s_axi_control_ARADDR,
	qsort_62_s_axi_control_RREADY,
	qsort_62_s_axi_control_RVALID,
	qsort_62_s_axi_control_RDATA,
	qsort_62_s_axi_control_RRESP,
	qsort_62_s_axi_control_AWREADY,
	qsort_62_s_axi_control_AWVALID,
	qsort_62_s_axi_control_AWADDR,
	qsort_62_s_axi_control_WREADY,
	qsort_62_s_axi_control_WVALID,
	qsort_62_s_axi_control_WDATA,
	qsort_62_s_axi_control_WSTRB,
	qsort_62_s_axi_control_BREADY,
	qsort_62_s_axi_control_BVALID,
	qsort_62_s_axi_control_BRESP,
	qsort_63_m_axi_gmem_ARREADY,
	qsort_63_m_axi_gmem_ARVALID,
	qsort_63_m_axi_gmem_ARID,
	qsort_63_m_axi_gmem_ARADDR,
	qsort_63_m_axi_gmem_ARLEN,
	qsort_63_m_axi_gmem_ARSIZE,
	qsort_63_m_axi_gmem_ARBURST,
	qsort_63_m_axi_gmem_ARLOCK,
	qsort_63_m_axi_gmem_ARCACHE,
	qsort_63_m_axi_gmem_ARPROT,
	qsort_63_m_axi_gmem_ARQOS,
	qsort_63_m_axi_gmem_ARREGION,
	qsort_63_m_axi_gmem_ARUSER,
	qsort_63_m_axi_gmem_RREADY,
	qsort_63_m_axi_gmem_RVALID,
	qsort_63_m_axi_gmem_RID,
	qsort_63_m_axi_gmem_RDATA,
	qsort_63_m_axi_gmem_RRESP,
	qsort_63_m_axi_gmem_RLAST,
	qsort_63_m_axi_gmem_RUSER,
	qsort_63_m_axi_gmem_AWREADY,
	qsort_63_m_axi_gmem_AWVALID,
	qsort_63_m_axi_gmem_AWID,
	qsort_63_m_axi_gmem_AWADDR,
	qsort_63_m_axi_gmem_AWLEN,
	qsort_63_m_axi_gmem_AWSIZE,
	qsort_63_m_axi_gmem_AWBURST,
	qsort_63_m_axi_gmem_AWLOCK,
	qsort_63_m_axi_gmem_AWCACHE,
	qsort_63_m_axi_gmem_AWPROT,
	qsort_63_m_axi_gmem_AWQOS,
	qsort_63_m_axi_gmem_AWREGION,
	qsort_63_m_axi_gmem_AWUSER,
	qsort_63_m_axi_gmem_WREADY,
	qsort_63_m_axi_gmem_WVALID,
	qsort_63_m_axi_gmem_WDATA,
	qsort_63_m_axi_gmem_WSTRB,
	qsort_63_m_axi_gmem_WLAST,
	qsort_63_m_axi_gmem_WUSER,
	qsort_63_m_axi_gmem_BREADY,
	qsort_63_m_axi_gmem_BVALID,
	qsort_63_m_axi_gmem_BID,
	qsort_63_m_axi_gmem_BRESP,
	qsort_63_m_axi_gmem_BUSER,
	qsort_63_s_axi_control_ARREADY,
	qsort_63_s_axi_control_ARVALID,
	qsort_63_s_axi_control_ARADDR,
	qsort_63_s_axi_control_RREADY,
	qsort_63_s_axi_control_RVALID,
	qsort_63_s_axi_control_RDATA,
	qsort_63_s_axi_control_RRESP,
	qsort_63_s_axi_control_AWREADY,
	qsort_63_s_axi_control_AWVALID,
	qsort_63_s_axi_control_AWADDR,
	qsort_63_s_axi_control_WREADY,
	qsort_63_s_axi_control_WVALID,
	qsort_63_s_axi_control_WDATA,
	qsort_63_s_axi_control_WSTRB,
	qsort_63_s_axi_control_BREADY,
	qsort_63_s_axi_control_BVALID,
	qsort_63_s_axi_control_BRESP,
	qsort_schedulerAXI_0_ARREADY,
	qsort_schedulerAXI_0_ARVALID,
	qsort_schedulerAXI_0_ARID,
	qsort_schedulerAXI_0_ARADDR,
	qsort_schedulerAXI_0_ARLEN,
	qsort_schedulerAXI_0_ARSIZE,
	qsort_schedulerAXI_0_ARBURST,
	qsort_schedulerAXI_0_ARLOCK,
	qsort_schedulerAXI_0_ARCACHE,
	qsort_schedulerAXI_0_ARPROT,
	qsort_schedulerAXI_0_ARQOS,
	qsort_schedulerAXI_0_ARREGION,
	qsort_schedulerAXI_0_RREADY,
	qsort_schedulerAXI_0_RVALID,
	qsort_schedulerAXI_0_RID,
	qsort_schedulerAXI_0_RDATA,
	qsort_schedulerAXI_0_RRESP,
	qsort_schedulerAXI_0_RLAST,
	qsort_schedulerAXI_0_AWREADY,
	qsort_schedulerAXI_0_AWVALID,
	qsort_schedulerAXI_0_AWID,
	qsort_schedulerAXI_0_AWADDR,
	qsort_schedulerAXI_0_AWLEN,
	qsort_schedulerAXI_0_AWSIZE,
	qsort_schedulerAXI_0_AWBURST,
	qsort_schedulerAXI_0_AWLOCK,
	qsort_schedulerAXI_0_AWCACHE,
	qsort_schedulerAXI_0_AWPROT,
	qsort_schedulerAXI_0_AWQOS,
	qsort_schedulerAXI_0_AWREGION,
	qsort_schedulerAXI_0_WREADY,
	qsort_schedulerAXI_0_WVALID,
	qsort_schedulerAXI_0_WDATA,
	qsort_schedulerAXI_0_WSTRB,
	qsort_schedulerAXI_0_WLAST,
	qsort_schedulerAXI_0_BREADY,
	qsort_schedulerAXI_0_BVALID,
	qsort_schedulerAXI_0_BID,
	qsort_schedulerAXI_0_BRESP,
	sync_schedulerAXI_0_ARREADY,
	sync_schedulerAXI_0_ARVALID,
	sync_schedulerAXI_0_ARID,
	sync_schedulerAXI_0_ARADDR,
	sync_schedulerAXI_0_ARLEN,
	sync_schedulerAXI_0_ARSIZE,
	sync_schedulerAXI_0_ARBURST,
	sync_schedulerAXI_0_ARLOCK,
	sync_schedulerAXI_0_ARCACHE,
	sync_schedulerAXI_0_ARPROT,
	sync_schedulerAXI_0_ARQOS,
	sync_schedulerAXI_0_ARREGION,
	sync_schedulerAXI_0_RREADY,
	sync_schedulerAXI_0_RVALID,
	sync_schedulerAXI_0_RID,
	sync_schedulerAXI_0_RDATA,
	sync_schedulerAXI_0_RRESP,
	sync_schedulerAXI_0_RLAST,
	sync_schedulerAXI_0_AWREADY,
	sync_schedulerAXI_0_AWVALID,
	sync_schedulerAXI_0_AWID,
	sync_schedulerAXI_0_AWADDR,
	sync_schedulerAXI_0_AWLEN,
	sync_schedulerAXI_0_AWSIZE,
	sync_schedulerAXI_0_AWBURST,
	sync_schedulerAXI_0_AWLOCK,
	sync_schedulerAXI_0_AWCACHE,
	sync_schedulerAXI_0_AWPROT,
	sync_schedulerAXI_0_AWQOS,
	sync_schedulerAXI_0_AWREGION,
	sync_schedulerAXI_0_WREADY,
	sync_schedulerAXI_0_WVALID,
	sync_schedulerAXI_0_WDATA,
	sync_schedulerAXI_0_WSTRB,
	sync_schedulerAXI_0_WLAST,
	sync_schedulerAXI_0_BREADY,
	sync_schedulerAXI_0_BVALID,
	sync_schedulerAXI_0_BID,
	sync_schedulerAXI_0_BRESP,
	sync_closureAllocatorAXI_0_ARREADY,
	sync_closureAllocatorAXI_0_ARVALID,
	sync_closureAllocatorAXI_0_ARID,
	sync_closureAllocatorAXI_0_ARADDR,
	sync_closureAllocatorAXI_0_ARLEN,
	sync_closureAllocatorAXI_0_ARSIZE,
	sync_closureAllocatorAXI_0_ARBURST,
	sync_closureAllocatorAXI_0_ARLOCK,
	sync_closureAllocatorAXI_0_ARCACHE,
	sync_closureAllocatorAXI_0_ARPROT,
	sync_closureAllocatorAXI_0_ARQOS,
	sync_closureAllocatorAXI_0_ARREGION,
	sync_closureAllocatorAXI_0_RREADY,
	sync_closureAllocatorAXI_0_RVALID,
	sync_closureAllocatorAXI_0_RID,
	sync_closureAllocatorAXI_0_RDATA,
	sync_closureAllocatorAXI_0_RRESP,
	sync_closureAllocatorAXI_0_RLAST,
	sync_closureAllocatorAXI_0_AWREADY,
	sync_closureAllocatorAXI_0_AWVALID,
	sync_closureAllocatorAXI_0_AWID,
	sync_closureAllocatorAXI_0_AWADDR,
	sync_closureAllocatorAXI_0_AWLEN,
	sync_closureAllocatorAXI_0_AWSIZE,
	sync_closureAllocatorAXI_0_AWBURST,
	sync_closureAllocatorAXI_0_AWLOCK,
	sync_closureAllocatorAXI_0_AWCACHE,
	sync_closureAllocatorAXI_0_AWPROT,
	sync_closureAllocatorAXI_0_AWQOS,
	sync_closureAllocatorAXI_0_AWREGION,
	sync_closureAllocatorAXI_0_WREADY,
	sync_closureAllocatorAXI_0_WVALID,
	sync_closureAllocatorAXI_0_WDATA,
	sync_closureAllocatorAXI_0_WSTRB,
	sync_closureAllocatorAXI_0_WLAST,
	sync_closureAllocatorAXI_0_BREADY,
	sync_closureAllocatorAXI_0_BVALID,
	sync_closureAllocatorAXI_0_BID,
	sync_closureAllocatorAXI_0_BRESP,
	sync_closureAllocatorAXI_1_ARREADY,
	sync_closureAllocatorAXI_1_ARVALID,
	sync_closureAllocatorAXI_1_ARID,
	sync_closureAllocatorAXI_1_ARADDR,
	sync_closureAllocatorAXI_1_ARLEN,
	sync_closureAllocatorAXI_1_ARSIZE,
	sync_closureAllocatorAXI_1_ARBURST,
	sync_closureAllocatorAXI_1_ARLOCK,
	sync_closureAllocatorAXI_1_ARCACHE,
	sync_closureAllocatorAXI_1_ARPROT,
	sync_closureAllocatorAXI_1_ARQOS,
	sync_closureAllocatorAXI_1_ARREGION,
	sync_closureAllocatorAXI_1_RREADY,
	sync_closureAllocatorAXI_1_RVALID,
	sync_closureAllocatorAXI_1_RID,
	sync_closureAllocatorAXI_1_RDATA,
	sync_closureAllocatorAXI_1_RRESP,
	sync_closureAllocatorAXI_1_RLAST,
	sync_closureAllocatorAXI_1_AWREADY,
	sync_closureAllocatorAXI_1_AWVALID,
	sync_closureAllocatorAXI_1_AWID,
	sync_closureAllocatorAXI_1_AWADDR,
	sync_closureAllocatorAXI_1_AWLEN,
	sync_closureAllocatorAXI_1_AWSIZE,
	sync_closureAllocatorAXI_1_AWBURST,
	sync_closureAllocatorAXI_1_AWLOCK,
	sync_closureAllocatorAXI_1_AWCACHE,
	sync_closureAllocatorAXI_1_AWPROT,
	sync_closureAllocatorAXI_1_AWQOS,
	sync_closureAllocatorAXI_1_AWREGION,
	sync_closureAllocatorAXI_1_WREADY,
	sync_closureAllocatorAXI_1_WVALID,
	sync_closureAllocatorAXI_1_WDATA,
	sync_closureAllocatorAXI_1_WSTRB,
	sync_closureAllocatorAXI_1_WLAST,
	sync_closureAllocatorAXI_1_BREADY,
	sync_closureAllocatorAXI_1_BVALID,
	sync_closureAllocatorAXI_1_BID,
	sync_closureAllocatorAXI_1_BRESP,
	sync_closureAllocatorAXI_2_ARREADY,
	sync_closureAllocatorAXI_2_ARVALID,
	sync_closureAllocatorAXI_2_ARID,
	sync_closureAllocatorAXI_2_ARADDR,
	sync_closureAllocatorAXI_2_ARLEN,
	sync_closureAllocatorAXI_2_ARSIZE,
	sync_closureAllocatorAXI_2_ARBURST,
	sync_closureAllocatorAXI_2_ARLOCK,
	sync_closureAllocatorAXI_2_ARCACHE,
	sync_closureAllocatorAXI_2_ARPROT,
	sync_closureAllocatorAXI_2_ARQOS,
	sync_closureAllocatorAXI_2_ARREGION,
	sync_closureAllocatorAXI_2_RREADY,
	sync_closureAllocatorAXI_2_RVALID,
	sync_closureAllocatorAXI_2_RID,
	sync_closureAllocatorAXI_2_RDATA,
	sync_closureAllocatorAXI_2_RRESP,
	sync_closureAllocatorAXI_2_RLAST,
	sync_closureAllocatorAXI_2_AWREADY,
	sync_closureAllocatorAXI_2_AWVALID,
	sync_closureAllocatorAXI_2_AWID,
	sync_closureAllocatorAXI_2_AWADDR,
	sync_closureAllocatorAXI_2_AWLEN,
	sync_closureAllocatorAXI_2_AWSIZE,
	sync_closureAllocatorAXI_2_AWBURST,
	sync_closureAllocatorAXI_2_AWLOCK,
	sync_closureAllocatorAXI_2_AWCACHE,
	sync_closureAllocatorAXI_2_AWPROT,
	sync_closureAllocatorAXI_2_AWQOS,
	sync_closureAllocatorAXI_2_AWREGION,
	sync_closureAllocatorAXI_2_WREADY,
	sync_closureAllocatorAXI_2_WVALID,
	sync_closureAllocatorAXI_2_WDATA,
	sync_closureAllocatorAXI_2_WSTRB,
	sync_closureAllocatorAXI_2_WLAST,
	sync_closureAllocatorAXI_2_BREADY,
	sync_closureAllocatorAXI_2_BVALID,
	sync_closureAllocatorAXI_2_BID,
	sync_closureAllocatorAXI_2_BRESP,
	sync_closureAllocatorAXI_3_ARREADY,
	sync_closureAllocatorAXI_3_ARVALID,
	sync_closureAllocatorAXI_3_ARID,
	sync_closureAllocatorAXI_3_ARADDR,
	sync_closureAllocatorAXI_3_ARLEN,
	sync_closureAllocatorAXI_3_ARSIZE,
	sync_closureAllocatorAXI_3_ARBURST,
	sync_closureAllocatorAXI_3_ARLOCK,
	sync_closureAllocatorAXI_3_ARCACHE,
	sync_closureAllocatorAXI_3_ARPROT,
	sync_closureAllocatorAXI_3_ARQOS,
	sync_closureAllocatorAXI_3_ARREGION,
	sync_closureAllocatorAXI_3_RREADY,
	sync_closureAllocatorAXI_3_RVALID,
	sync_closureAllocatorAXI_3_RID,
	sync_closureAllocatorAXI_3_RDATA,
	sync_closureAllocatorAXI_3_RRESP,
	sync_closureAllocatorAXI_3_RLAST,
	sync_closureAllocatorAXI_3_AWREADY,
	sync_closureAllocatorAXI_3_AWVALID,
	sync_closureAllocatorAXI_3_AWID,
	sync_closureAllocatorAXI_3_AWADDR,
	sync_closureAllocatorAXI_3_AWLEN,
	sync_closureAllocatorAXI_3_AWSIZE,
	sync_closureAllocatorAXI_3_AWBURST,
	sync_closureAllocatorAXI_3_AWLOCK,
	sync_closureAllocatorAXI_3_AWCACHE,
	sync_closureAllocatorAXI_3_AWPROT,
	sync_closureAllocatorAXI_3_AWQOS,
	sync_closureAllocatorAXI_3_AWREGION,
	sync_closureAllocatorAXI_3_WREADY,
	sync_closureAllocatorAXI_3_WVALID,
	sync_closureAllocatorAXI_3_WDATA,
	sync_closureAllocatorAXI_3_WSTRB,
	sync_closureAllocatorAXI_3_WLAST,
	sync_closureAllocatorAXI_3_BREADY,
	sync_closureAllocatorAXI_3_BVALID,
	sync_closureAllocatorAXI_3_BID,
	sync_closureAllocatorAXI_3_BRESP,
	sync_argumentNotifierAXI_0_ARREADY,
	sync_argumentNotifierAXI_0_ARVALID,
	sync_argumentNotifierAXI_0_ARADDR,
	sync_argumentNotifierAXI_0_ARLEN,
	sync_argumentNotifierAXI_0_ARSIZE,
	sync_argumentNotifierAXI_0_ARBURST,
	sync_argumentNotifierAXI_0_ARLOCK,
	sync_argumentNotifierAXI_0_ARCACHE,
	sync_argumentNotifierAXI_0_ARPROT,
	sync_argumentNotifierAXI_0_ARQOS,
	sync_argumentNotifierAXI_0_ARREGION,
	sync_argumentNotifierAXI_0_RREADY,
	sync_argumentNotifierAXI_0_RVALID,
	sync_argumentNotifierAXI_0_RDATA,
	sync_argumentNotifierAXI_0_RRESP,
	sync_argumentNotifierAXI_0_RLAST,
	sync_argumentNotifierAXI_0_AWREADY,
	sync_argumentNotifierAXI_0_AWVALID,
	sync_argumentNotifierAXI_0_AWADDR,
	sync_argumentNotifierAXI_0_AWLEN,
	sync_argumentNotifierAXI_0_AWSIZE,
	sync_argumentNotifierAXI_0_AWBURST,
	sync_argumentNotifierAXI_0_AWLOCK,
	sync_argumentNotifierAXI_0_AWCACHE,
	sync_argumentNotifierAXI_0_AWPROT,
	sync_argumentNotifierAXI_0_AWQOS,
	sync_argumentNotifierAXI_0_AWREGION,
	sync_argumentNotifierAXI_0_WREADY,
	sync_argumentNotifierAXI_0_WVALID,
	sync_argumentNotifierAXI_0_WDATA,
	sync_argumentNotifierAXI_0_WSTRB,
	sync_argumentNotifierAXI_0_WLAST,
	sync_argumentNotifierAXI_0_BREADY,
	sync_argumentNotifierAXI_0_BVALID,
	sync_argumentNotifierAXI_0_BRESP,
	sync_argumentNotifierAXI_1_ARREADY,
	sync_argumentNotifierAXI_1_ARVALID,
	sync_argumentNotifierAXI_1_ARADDR,
	sync_argumentNotifierAXI_1_ARLEN,
	sync_argumentNotifierAXI_1_ARSIZE,
	sync_argumentNotifierAXI_1_ARBURST,
	sync_argumentNotifierAXI_1_ARLOCK,
	sync_argumentNotifierAXI_1_ARCACHE,
	sync_argumentNotifierAXI_1_ARPROT,
	sync_argumentNotifierAXI_1_ARQOS,
	sync_argumentNotifierAXI_1_ARREGION,
	sync_argumentNotifierAXI_1_RREADY,
	sync_argumentNotifierAXI_1_RVALID,
	sync_argumentNotifierAXI_1_RDATA,
	sync_argumentNotifierAXI_1_RRESP,
	sync_argumentNotifierAXI_1_RLAST,
	sync_argumentNotifierAXI_1_AWREADY,
	sync_argumentNotifierAXI_1_AWVALID,
	sync_argumentNotifierAXI_1_AWADDR,
	sync_argumentNotifierAXI_1_AWLEN,
	sync_argumentNotifierAXI_1_AWSIZE,
	sync_argumentNotifierAXI_1_AWBURST,
	sync_argumentNotifierAXI_1_AWLOCK,
	sync_argumentNotifierAXI_1_AWCACHE,
	sync_argumentNotifierAXI_1_AWPROT,
	sync_argumentNotifierAXI_1_AWQOS,
	sync_argumentNotifierAXI_1_AWREGION,
	sync_argumentNotifierAXI_1_WREADY,
	sync_argumentNotifierAXI_1_WVALID,
	sync_argumentNotifierAXI_1_WDATA,
	sync_argumentNotifierAXI_1_WSTRB,
	sync_argumentNotifierAXI_1_WLAST,
	sync_argumentNotifierAXI_1_BREADY,
	sync_argumentNotifierAXI_1_BVALID,
	sync_argumentNotifierAXI_1_BRESP,
	sync_argumentNotifierAXI_2_ARREADY,
	sync_argumentNotifierAXI_2_ARVALID,
	sync_argumentNotifierAXI_2_ARADDR,
	sync_argumentNotifierAXI_2_ARLEN,
	sync_argumentNotifierAXI_2_ARSIZE,
	sync_argumentNotifierAXI_2_ARBURST,
	sync_argumentNotifierAXI_2_ARLOCK,
	sync_argumentNotifierAXI_2_ARCACHE,
	sync_argumentNotifierAXI_2_ARPROT,
	sync_argumentNotifierAXI_2_ARQOS,
	sync_argumentNotifierAXI_2_ARREGION,
	sync_argumentNotifierAXI_2_RREADY,
	sync_argumentNotifierAXI_2_RVALID,
	sync_argumentNotifierAXI_2_RDATA,
	sync_argumentNotifierAXI_2_RRESP,
	sync_argumentNotifierAXI_2_RLAST,
	sync_argumentNotifierAXI_2_AWREADY,
	sync_argumentNotifierAXI_2_AWVALID,
	sync_argumentNotifierAXI_2_AWADDR,
	sync_argumentNotifierAXI_2_AWLEN,
	sync_argumentNotifierAXI_2_AWSIZE,
	sync_argumentNotifierAXI_2_AWBURST,
	sync_argumentNotifierAXI_2_AWLOCK,
	sync_argumentNotifierAXI_2_AWCACHE,
	sync_argumentNotifierAXI_2_AWPROT,
	sync_argumentNotifierAXI_2_AWQOS,
	sync_argumentNotifierAXI_2_AWREGION,
	sync_argumentNotifierAXI_2_WREADY,
	sync_argumentNotifierAXI_2_WVALID,
	sync_argumentNotifierAXI_2_WDATA,
	sync_argumentNotifierAXI_2_WSTRB,
	sync_argumentNotifierAXI_2_WLAST,
	sync_argumentNotifierAXI_2_BREADY,
	sync_argumentNotifierAXI_2_BVALID,
	sync_argumentNotifierAXI_2_BRESP,
	sync_argumentNotifierAXI_3_ARREADY,
	sync_argumentNotifierAXI_3_ARVALID,
	sync_argumentNotifierAXI_3_ARADDR,
	sync_argumentNotifierAXI_3_ARLEN,
	sync_argumentNotifierAXI_3_ARSIZE,
	sync_argumentNotifierAXI_3_ARBURST,
	sync_argumentNotifierAXI_3_ARLOCK,
	sync_argumentNotifierAXI_3_ARCACHE,
	sync_argumentNotifierAXI_3_ARPROT,
	sync_argumentNotifierAXI_3_ARQOS,
	sync_argumentNotifierAXI_3_ARREGION,
	sync_argumentNotifierAXI_3_RREADY,
	sync_argumentNotifierAXI_3_RVALID,
	sync_argumentNotifierAXI_3_RDATA,
	sync_argumentNotifierAXI_3_RRESP,
	sync_argumentNotifierAXI_3_RLAST,
	sync_argumentNotifierAXI_3_AWREADY,
	sync_argumentNotifierAXI_3_AWVALID,
	sync_argumentNotifierAXI_3_AWADDR,
	sync_argumentNotifierAXI_3_AWLEN,
	sync_argumentNotifierAXI_3_AWSIZE,
	sync_argumentNotifierAXI_3_AWBURST,
	sync_argumentNotifierAXI_3_AWLOCK,
	sync_argumentNotifierAXI_3_AWCACHE,
	sync_argumentNotifierAXI_3_AWPROT,
	sync_argumentNotifierAXI_3_AWQOS,
	sync_argumentNotifierAXI_3_AWREGION,
	sync_argumentNotifierAXI_3_WREADY,
	sync_argumentNotifierAXI_3_WVALID,
	sync_argumentNotifierAXI_3_WDATA,
	sync_argumentNotifierAXI_3_WSTRB,
	sync_argumentNotifierAXI_3_WLAST,
	sync_argumentNotifierAXI_3_BREADY,
	sync_argumentNotifierAXI_3_BVALID,
	sync_argumentNotifierAXI_3_BRESP,
	sync_argumentNotifierAXI_4_ARREADY,
	sync_argumentNotifierAXI_4_ARVALID,
	sync_argumentNotifierAXI_4_ARADDR,
	sync_argumentNotifierAXI_4_ARLEN,
	sync_argumentNotifierAXI_4_ARSIZE,
	sync_argumentNotifierAXI_4_ARBURST,
	sync_argumentNotifierAXI_4_ARLOCK,
	sync_argumentNotifierAXI_4_ARCACHE,
	sync_argumentNotifierAXI_4_ARPROT,
	sync_argumentNotifierAXI_4_ARQOS,
	sync_argumentNotifierAXI_4_ARREGION,
	sync_argumentNotifierAXI_4_RREADY,
	sync_argumentNotifierAXI_4_RVALID,
	sync_argumentNotifierAXI_4_RDATA,
	sync_argumentNotifierAXI_4_RRESP,
	sync_argumentNotifierAXI_4_RLAST,
	sync_argumentNotifierAXI_4_AWREADY,
	sync_argumentNotifierAXI_4_AWVALID,
	sync_argumentNotifierAXI_4_AWADDR,
	sync_argumentNotifierAXI_4_AWLEN,
	sync_argumentNotifierAXI_4_AWSIZE,
	sync_argumentNotifierAXI_4_AWBURST,
	sync_argumentNotifierAXI_4_AWLOCK,
	sync_argumentNotifierAXI_4_AWCACHE,
	sync_argumentNotifierAXI_4_AWPROT,
	sync_argumentNotifierAXI_4_AWQOS,
	sync_argumentNotifierAXI_4_AWREGION,
	sync_argumentNotifierAXI_4_WREADY,
	sync_argumentNotifierAXI_4_WVALID,
	sync_argumentNotifierAXI_4_WDATA,
	sync_argumentNotifierAXI_4_WSTRB,
	sync_argumentNotifierAXI_4_WLAST,
	sync_argumentNotifierAXI_4_BREADY,
	sync_argumentNotifierAXI_4_BVALID,
	sync_argumentNotifierAXI_4_BRESP,
	sync_argumentNotifierAXI_5_ARREADY,
	sync_argumentNotifierAXI_5_ARVALID,
	sync_argumentNotifierAXI_5_ARADDR,
	sync_argumentNotifierAXI_5_ARLEN,
	sync_argumentNotifierAXI_5_ARSIZE,
	sync_argumentNotifierAXI_5_ARBURST,
	sync_argumentNotifierAXI_5_ARLOCK,
	sync_argumentNotifierAXI_5_ARCACHE,
	sync_argumentNotifierAXI_5_ARPROT,
	sync_argumentNotifierAXI_5_ARQOS,
	sync_argumentNotifierAXI_5_ARREGION,
	sync_argumentNotifierAXI_5_RREADY,
	sync_argumentNotifierAXI_5_RVALID,
	sync_argumentNotifierAXI_5_RDATA,
	sync_argumentNotifierAXI_5_RRESP,
	sync_argumentNotifierAXI_5_RLAST,
	sync_argumentNotifierAXI_5_AWREADY,
	sync_argumentNotifierAXI_5_AWVALID,
	sync_argumentNotifierAXI_5_AWADDR,
	sync_argumentNotifierAXI_5_AWLEN,
	sync_argumentNotifierAXI_5_AWSIZE,
	sync_argumentNotifierAXI_5_AWBURST,
	sync_argumentNotifierAXI_5_AWLOCK,
	sync_argumentNotifierAXI_5_AWCACHE,
	sync_argumentNotifierAXI_5_AWPROT,
	sync_argumentNotifierAXI_5_AWQOS,
	sync_argumentNotifierAXI_5_AWREGION,
	sync_argumentNotifierAXI_5_WREADY,
	sync_argumentNotifierAXI_5_WVALID,
	sync_argumentNotifierAXI_5_WDATA,
	sync_argumentNotifierAXI_5_WSTRB,
	sync_argumentNotifierAXI_5_WLAST,
	sync_argumentNotifierAXI_5_BREADY,
	sync_argumentNotifierAXI_5_BVALID,
	sync_argumentNotifierAXI_5_BRESP,
	sync_argumentNotifierAXI_6_ARREADY,
	sync_argumentNotifierAXI_6_ARVALID,
	sync_argumentNotifierAXI_6_ARADDR,
	sync_argumentNotifierAXI_6_ARLEN,
	sync_argumentNotifierAXI_6_ARSIZE,
	sync_argumentNotifierAXI_6_ARBURST,
	sync_argumentNotifierAXI_6_ARLOCK,
	sync_argumentNotifierAXI_6_ARCACHE,
	sync_argumentNotifierAXI_6_ARPROT,
	sync_argumentNotifierAXI_6_ARQOS,
	sync_argumentNotifierAXI_6_ARREGION,
	sync_argumentNotifierAXI_6_RREADY,
	sync_argumentNotifierAXI_6_RVALID,
	sync_argumentNotifierAXI_6_RDATA,
	sync_argumentNotifierAXI_6_RRESP,
	sync_argumentNotifierAXI_6_RLAST,
	sync_argumentNotifierAXI_6_AWREADY,
	sync_argumentNotifierAXI_6_AWVALID,
	sync_argumentNotifierAXI_6_AWADDR,
	sync_argumentNotifierAXI_6_AWLEN,
	sync_argumentNotifierAXI_6_AWSIZE,
	sync_argumentNotifierAXI_6_AWBURST,
	sync_argumentNotifierAXI_6_AWLOCK,
	sync_argumentNotifierAXI_6_AWCACHE,
	sync_argumentNotifierAXI_6_AWPROT,
	sync_argumentNotifierAXI_6_AWQOS,
	sync_argumentNotifierAXI_6_AWREGION,
	sync_argumentNotifierAXI_6_WREADY,
	sync_argumentNotifierAXI_6_WVALID,
	sync_argumentNotifierAXI_6_WDATA,
	sync_argumentNotifierAXI_6_WSTRB,
	sync_argumentNotifierAXI_6_WLAST,
	sync_argumentNotifierAXI_6_BREADY,
	sync_argumentNotifierAXI_6_BVALID,
	sync_argumentNotifierAXI_6_BRESP,
	sync_argumentNotifierAXI_7_ARREADY,
	sync_argumentNotifierAXI_7_ARVALID,
	sync_argumentNotifierAXI_7_ARADDR,
	sync_argumentNotifierAXI_7_ARLEN,
	sync_argumentNotifierAXI_7_ARSIZE,
	sync_argumentNotifierAXI_7_ARBURST,
	sync_argumentNotifierAXI_7_ARLOCK,
	sync_argumentNotifierAXI_7_ARCACHE,
	sync_argumentNotifierAXI_7_ARPROT,
	sync_argumentNotifierAXI_7_ARQOS,
	sync_argumentNotifierAXI_7_ARREGION,
	sync_argumentNotifierAXI_7_RREADY,
	sync_argumentNotifierAXI_7_RVALID,
	sync_argumentNotifierAXI_7_RDATA,
	sync_argumentNotifierAXI_7_RRESP,
	sync_argumentNotifierAXI_7_RLAST,
	sync_argumentNotifierAXI_7_AWREADY,
	sync_argumentNotifierAXI_7_AWVALID,
	sync_argumentNotifierAXI_7_AWADDR,
	sync_argumentNotifierAXI_7_AWLEN,
	sync_argumentNotifierAXI_7_AWSIZE,
	sync_argumentNotifierAXI_7_AWBURST,
	sync_argumentNotifierAXI_7_AWLOCK,
	sync_argumentNotifierAXI_7_AWCACHE,
	sync_argumentNotifierAXI_7_AWPROT,
	sync_argumentNotifierAXI_7_AWQOS,
	sync_argumentNotifierAXI_7_AWREGION,
	sync_argumentNotifierAXI_7_WREADY,
	sync_argumentNotifierAXI_7_WVALID,
	sync_argumentNotifierAXI_7_WDATA,
	sync_argumentNotifierAXI_7_WSTRB,
	sync_argumentNotifierAXI_7_WLAST,
	sync_argumentNotifierAXI_7_BREADY,
	sync_argumentNotifierAXI_7_BVALID,
	sync_argumentNotifierAXI_7_BRESP,
	sync_argumentNotifierAXI_8_ARREADY,
	sync_argumentNotifierAXI_8_ARVALID,
	sync_argumentNotifierAXI_8_ARADDR,
	sync_argumentNotifierAXI_8_ARLEN,
	sync_argumentNotifierAXI_8_ARSIZE,
	sync_argumentNotifierAXI_8_ARBURST,
	sync_argumentNotifierAXI_8_ARLOCK,
	sync_argumentNotifierAXI_8_ARCACHE,
	sync_argumentNotifierAXI_8_ARPROT,
	sync_argumentNotifierAXI_8_ARQOS,
	sync_argumentNotifierAXI_8_ARREGION,
	sync_argumentNotifierAXI_8_RREADY,
	sync_argumentNotifierAXI_8_RVALID,
	sync_argumentNotifierAXI_8_RDATA,
	sync_argumentNotifierAXI_8_RRESP,
	sync_argumentNotifierAXI_8_RLAST,
	sync_argumentNotifierAXI_8_AWREADY,
	sync_argumentNotifierAXI_8_AWVALID,
	sync_argumentNotifierAXI_8_AWADDR,
	sync_argumentNotifierAXI_8_AWLEN,
	sync_argumentNotifierAXI_8_AWSIZE,
	sync_argumentNotifierAXI_8_AWBURST,
	sync_argumentNotifierAXI_8_AWLOCK,
	sync_argumentNotifierAXI_8_AWCACHE,
	sync_argumentNotifierAXI_8_AWPROT,
	sync_argumentNotifierAXI_8_AWQOS,
	sync_argumentNotifierAXI_8_AWREGION,
	sync_argumentNotifierAXI_8_WREADY,
	sync_argumentNotifierAXI_8_WVALID,
	sync_argumentNotifierAXI_8_WDATA,
	sync_argumentNotifierAXI_8_WSTRB,
	sync_argumentNotifierAXI_8_WLAST,
	sync_argumentNotifierAXI_8_BREADY,
	sync_argumentNotifierAXI_8_BVALID,
	sync_argumentNotifierAXI_8_BRESP,
	sync_argumentNotifierAXI_9_ARREADY,
	sync_argumentNotifierAXI_9_ARVALID,
	sync_argumentNotifierAXI_9_ARADDR,
	sync_argumentNotifierAXI_9_ARLEN,
	sync_argumentNotifierAXI_9_ARSIZE,
	sync_argumentNotifierAXI_9_ARBURST,
	sync_argumentNotifierAXI_9_ARLOCK,
	sync_argumentNotifierAXI_9_ARCACHE,
	sync_argumentNotifierAXI_9_ARPROT,
	sync_argumentNotifierAXI_9_ARQOS,
	sync_argumentNotifierAXI_9_ARREGION,
	sync_argumentNotifierAXI_9_RREADY,
	sync_argumentNotifierAXI_9_RVALID,
	sync_argumentNotifierAXI_9_RDATA,
	sync_argumentNotifierAXI_9_RRESP,
	sync_argumentNotifierAXI_9_RLAST,
	sync_argumentNotifierAXI_9_AWREADY,
	sync_argumentNotifierAXI_9_AWVALID,
	sync_argumentNotifierAXI_9_AWADDR,
	sync_argumentNotifierAXI_9_AWLEN,
	sync_argumentNotifierAXI_9_AWSIZE,
	sync_argumentNotifierAXI_9_AWBURST,
	sync_argumentNotifierAXI_9_AWLOCK,
	sync_argumentNotifierAXI_9_AWCACHE,
	sync_argumentNotifierAXI_9_AWPROT,
	sync_argumentNotifierAXI_9_AWQOS,
	sync_argumentNotifierAXI_9_AWREGION,
	sync_argumentNotifierAXI_9_WREADY,
	sync_argumentNotifierAXI_9_WVALID,
	sync_argumentNotifierAXI_9_WDATA,
	sync_argumentNotifierAXI_9_WSTRB,
	sync_argumentNotifierAXI_9_WLAST,
	sync_argumentNotifierAXI_9_BREADY,
	sync_argumentNotifierAXI_9_BVALID,
	sync_argumentNotifierAXI_9_BRESP,
	sync_argumentNotifierAXI_10_ARREADY,
	sync_argumentNotifierAXI_10_ARVALID,
	sync_argumentNotifierAXI_10_ARADDR,
	sync_argumentNotifierAXI_10_ARLEN,
	sync_argumentNotifierAXI_10_ARSIZE,
	sync_argumentNotifierAXI_10_ARBURST,
	sync_argumentNotifierAXI_10_ARLOCK,
	sync_argumentNotifierAXI_10_ARCACHE,
	sync_argumentNotifierAXI_10_ARPROT,
	sync_argumentNotifierAXI_10_ARQOS,
	sync_argumentNotifierAXI_10_ARREGION,
	sync_argumentNotifierAXI_10_RREADY,
	sync_argumentNotifierAXI_10_RVALID,
	sync_argumentNotifierAXI_10_RDATA,
	sync_argumentNotifierAXI_10_RRESP,
	sync_argumentNotifierAXI_10_RLAST,
	sync_argumentNotifierAXI_10_AWREADY,
	sync_argumentNotifierAXI_10_AWVALID,
	sync_argumentNotifierAXI_10_AWADDR,
	sync_argumentNotifierAXI_10_AWLEN,
	sync_argumentNotifierAXI_10_AWSIZE,
	sync_argumentNotifierAXI_10_AWBURST,
	sync_argumentNotifierAXI_10_AWLOCK,
	sync_argumentNotifierAXI_10_AWCACHE,
	sync_argumentNotifierAXI_10_AWPROT,
	sync_argumentNotifierAXI_10_AWQOS,
	sync_argumentNotifierAXI_10_AWREGION,
	sync_argumentNotifierAXI_10_WREADY,
	sync_argumentNotifierAXI_10_WVALID,
	sync_argumentNotifierAXI_10_WDATA,
	sync_argumentNotifierAXI_10_WSTRB,
	sync_argumentNotifierAXI_10_WLAST,
	sync_argumentNotifierAXI_10_BREADY,
	sync_argumentNotifierAXI_10_BVALID,
	sync_argumentNotifierAXI_10_BRESP,
	sync_argumentNotifierAXI_11_ARREADY,
	sync_argumentNotifierAXI_11_ARVALID,
	sync_argumentNotifierAXI_11_ARADDR,
	sync_argumentNotifierAXI_11_ARLEN,
	sync_argumentNotifierAXI_11_ARSIZE,
	sync_argumentNotifierAXI_11_ARBURST,
	sync_argumentNotifierAXI_11_ARLOCK,
	sync_argumentNotifierAXI_11_ARCACHE,
	sync_argumentNotifierAXI_11_ARPROT,
	sync_argumentNotifierAXI_11_ARQOS,
	sync_argumentNotifierAXI_11_ARREGION,
	sync_argumentNotifierAXI_11_RREADY,
	sync_argumentNotifierAXI_11_RVALID,
	sync_argumentNotifierAXI_11_RDATA,
	sync_argumentNotifierAXI_11_RRESP,
	sync_argumentNotifierAXI_11_RLAST,
	sync_argumentNotifierAXI_11_AWREADY,
	sync_argumentNotifierAXI_11_AWVALID,
	sync_argumentNotifierAXI_11_AWADDR,
	sync_argumentNotifierAXI_11_AWLEN,
	sync_argumentNotifierAXI_11_AWSIZE,
	sync_argumentNotifierAXI_11_AWBURST,
	sync_argumentNotifierAXI_11_AWLOCK,
	sync_argumentNotifierAXI_11_AWCACHE,
	sync_argumentNotifierAXI_11_AWPROT,
	sync_argumentNotifierAXI_11_AWQOS,
	sync_argumentNotifierAXI_11_AWREGION,
	sync_argumentNotifierAXI_11_WREADY,
	sync_argumentNotifierAXI_11_WVALID,
	sync_argumentNotifierAXI_11_WDATA,
	sync_argumentNotifierAXI_11_WSTRB,
	sync_argumentNotifierAXI_11_WLAST,
	sync_argumentNotifierAXI_11_BREADY,
	sync_argumentNotifierAXI_11_BVALID,
	sync_argumentNotifierAXI_11_BRESP,
	sync_argumentNotifierAXI_12_ARREADY,
	sync_argumentNotifierAXI_12_ARVALID,
	sync_argumentNotifierAXI_12_ARADDR,
	sync_argumentNotifierAXI_12_ARLEN,
	sync_argumentNotifierAXI_12_ARSIZE,
	sync_argumentNotifierAXI_12_ARBURST,
	sync_argumentNotifierAXI_12_ARLOCK,
	sync_argumentNotifierAXI_12_ARCACHE,
	sync_argumentNotifierAXI_12_ARPROT,
	sync_argumentNotifierAXI_12_ARQOS,
	sync_argumentNotifierAXI_12_ARREGION,
	sync_argumentNotifierAXI_12_RREADY,
	sync_argumentNotifierAXI_12_RVALID,
	sync_argumentNotifierAXI_12_RDATA,
	sync_argumentNotifierAXI_12_RRESP,
	sync_argumentNotifierAXI_12_RLAST,
	sync_argumentNotifierAXI_12_AWREADY,
	sync_argumentNotifierAXI_12_AWVALID,
	sync_argumentNotifierAXI_12_AWADDR,
	sync_argumentNotifierAXI_12_AWLEN,
	sync_argumentNotifierAXI_12_AWSIZE,
	sync_argumentNotifierAXI_12_AWBURST,
	sync_argumentNotifierAXI_12_AWLOCK,
	sync_argumentNotifierAXI_12_AWCACHE,
	sync_argumentNotifierAXI_12_AWPROT,
	sync_argumentNotifierAXI_12_AWQOS,
	sync_argumentNotifierAXI_12_AWREGION,
	sync_argumentNotifierAXI_12_WREADY,
	sync_argumentNotifierAXI_12_WVALID,
	sync_argumentNotifierAXI_12_WDATA,
	sync_argumentNotifierAXI_12_WSTRB,
	sync_argumentNotifierAXI_12_WLAST,
	sync_argumentNotifierAXI_12_BREADY,
	sync_argumentNotifierAXI_12_BVALID,
	sync_argumentNotifierAXI_12_BRESP,
	sync_argumentNotifierAXI_13_ARREADY,
	sync_argumentNotifierAXI_13_ARVALID,
	sync_argumentNotifierAXI_13_ARADDR,
	sync_argumentNotifierAXI_13_ARLEN,
	sync_argumentNotifierAXI_13_ARSIZE,
	sync_argumentNotifierAXI_13_ARBURST,
	sync_argumentNotifierAXI_13_ARLOCK,
	sync_argumentNotifierAXI_13_ARCACHE,
	sync_argumentNotifierAXI_13_ARPROT,
	sync_argumentNotifierAXI_13_ARQOS,
	sync_argumentNotifierAXI_13_ARREGION,
	sync_argumentNotifierAXI_13_RREADY,
	sync_argumentNotifierAXI_13_RVALID,
	sync_argumentNotifierAXI_13_RDATA,
	sync_argumentNotifierAXI_13_RRESP,
	sync_argumentNotifierAXI_13_RLAST,
	sync_argumentNotifierAXI_13_AWREADY,
	sync_argumentNotifierAXI_13_AWVALID,
	sync_argumentNotifierAXI_13_AWADDR,
	sync_argumentNotifierAXI_13_AWLEN,
	sync_argumentNotifierAXI_13_AWSIZE,
	sync_argumentNotifierAXI_13_AWBURST,
	sync_argumentNotifierAXI_13_AWLOCK,
	sync_argumentNotifierAXI_13_AWCACHE,
	sync_argumentNotifierAXI_13_AWPROT,
	sync_argumentNotifierAXI_13_AWQOS,
	sync_argumentNotifierAXI_13_AWREGION,
	sync_argumentNotifierAXI_13_WREADY,
	sync_argumentNotifierAXI_13_WVALID,
	sync_argumentNotifierAXI_13_WDATA,
	sync_argumentNotifierAXI_13_WSTRB,
	sync_argumentNotifierAXI_13_WLAST,
	sync_argumentNotifierAXI_13_BREADY,
	sync_argumentNotifierAXI_13_BVALID,
	sync_argumentNotifierAXI_13_BRESP,
	sync_argumentNotifierAXI_14_ARREADY,
	sync_argumentNotifierAXI_14_ARVALID,
	sync_argumentNotifierAXI_14_ARADDR,
	sync_argumentNotifierAXI_14_ARLEN,
	sync_argumentNotifierAXI_14_ARSIZE,
	sync_argumentNotifierAXI_14_ARBURST,
	sync_argumentNotifierAXI_14_ARLOCK,
	sync_argumentNotifierAXI_14_ARCACHE,
	sync_argumentNotifierAXI_14_ARPROT,
	sync_argumentNotifierAXI_14_ARQOS,
	sync_argumentNotifierAXI_14_ARREGION,
	sync_argumentNotifierAXI_14_RREADY,
	sync_argumentNotifierAXI_14_RVALID,
	sync_argumentNotifierAXI_14_RDATA,
	sync_argumentNotifierAXI_14_RRESP,
	sync_argumentNotifierAXI_14_RLAST,
	sync_argumentNotifierAXI_14_AWREADY,
	sync_argumentNotifierAXI_14_AWVALID,
	sync_argumentNotifierAXI_14_AWADDR,
	sync_argumentNotifierAXI_14_AWLEN,
	sync_argumentNotifierAXI_14_AWSIZE,
	sync_argumentNotifierAXI_14_AWBURST,
	sync_argumentNotifierAXI_14_AWLOCK,
	sync_argumentNotifierAXI_14_AWCACHE,
	sync_argumentNotifierAXI_14_AWPROT,
	sync_argumentNotifierAXI_14_AWQOS,
	sync_argumentNotifierAXI_14_AWREGION,
	sync_argumentNotifierAXI_14_WREADY,
	sync_argumentNotifierAXI_14_WVALID,
	sync_argumentNotifierAXI_14_WDATA,
	sync_argumentNotifierAXI_14_WSTRB,
	sync_argumentNotifierAXI_14_WLAST,
	sync_argumentNotifierAXI_14_BREADY,
	sync_argumentNotifierAXI_14_BVALID,
	sync_argumentNotifierAXI_14_BRESP,
	sync_argumentNotifierAXI_15_ARREADY,
	sync_argumentNotifierAXI_15_ARVALID,
	sync_argumentNotifierAXI_15_ARADDR,
	sync_argumentNotifierAXI_15_ARLEN,
	sync_argumentNotifierAXI_15_ARSIZE,
	sync_argumentNotifierAXI_15_ARBURST,
	sync_argumentNotifierAXI_15_ARLOCK,
	sync_argumentNotifierAXI_15_ARCACHE,
	sync_argumentNotifierAXI_15_ARPROT,
	sync_argumentNotifierAXI_15_ARQOS,
	sync_argumentNotifierAXI_15_ARREGION,
	sync_argumentNotifierAXI_15_RREADY,
	sync_argumentNotifierAXI_15_RVALID,
	sync_argumentNotifierAXI_15_RDATA,
	sync_argumentNotifierAXI_15_RRESP,
	sync_argumentNotifierAXI_15_RLAST,
	sync_argumentNotifierAXI_15_AWREADY,
	sync_argumentNotifierAXI_15_AWVALID,
	sync_argumentNotifierAXI_15_AWADDR,
	sync_argumentNotifierAXI_15_AWLEN,
	sync_argumentNotifierAXI_15_AWSIZE,
	sync_argumentNotifierAXI_15_AWBURST,
	sync_argumentNotifierAXI_15_AWLOCK,
	sync_argumentNotifierAXI_15_AWCACHE,
	sync_argumentNotifierAXI_15_AWPROT,
	sync_argumentNotifierAXI_15_AWQOS,
	sync_argumentNotifierAXI_15_AWREGION,
	sync_argumentNotifierAXI_15_WREADY,
	sync_argumentNotifierAXI_15_WVALID,
	sync_argumentNotifierAXI_15_WDATA,
	sync_argumentNotifierAXI_15_WSTRB,
	sync_argumentNotifierAXI_15_WLAST,
	sync_argumentNotifierAXI_15_BREADY,
	sync_argumentNotifierAXI_15_BVALID,
	sync_argumentNotifierAXI_15_BRESP,
	sync_argumentNotifierAXI_16_ARREADY,
	sync_argumentNotifierAXI_16_ARVALID,
	sync_argumentNotifierAXI_16_ARADDR,
	sync_argumentNotifierAXI_16_ARLEN,
	sync_argumentNotifierAXI_16_ARSIZE,
	sync_argumentNotifierAXI_16_ARBURST,
	sync_argumentNotifierAXI_16_ARLOCK,
	sync_argumentNotifierAXI_16_ARCACHE,
	sync_argumentNotifierAXI_16_ARPROT,
	sync_argumentNotifierAXI_16_ARQOS,
	sync_argumentNotifierAXI_16_ARREGION,
	sync_argumentNotifierAXI_16_RREADY,
	sync_argumentNotifierAXI_16_RVALID,
	sync_argumentNotifierAXI_16_RDATA,
	sync_argumentNotifierAXI_16_RRESP,
	sync_argumentNotifierAXI_16_RLAST,
	sync_argumentNotifierAXI_16_AWREADY,
	sync_argumentNotifierAXI_16_AWVALID,
	sync_argumentNotifierAXI_16_AWADDR,
	sync_argumentNotifierAXI_16_AWLEN,
	sync_argumentNotifierAXI_16_AWSIZE,
	sync_argumentNotifierAXI_16_AWBURST,
	sync_argumentNotifierAXI_16_AWLOCK,
	sync_argumentNotifierAXI_16_AWCACHE,
	sync_argumentNotifierAXI_16_AWPROT,
	sync_argumentNotifierAXI_16_AWQOS,
	sync_argumentNotifierAXI_16_AWREGION,
	sync_argumentNotifierAXI_16_WREADY,
	sync_argumentNotifierAXI_16_WVALID,
	sync_argumentNotifierAXI_16_WDATA,
	sync_argumentNotifierAXI_16_WSTRB,
	sync_argumentNotifierAXI_16_WLAST,
	sync_argumentNotifierAXI_16_BREADY,
	sync_argumentNotifierAXI_16_BVALID,
	sync_argumentNotifierAXI_16_BRESP,
	sync_argumentNotifierAXI_17_ARREADY,
	sync_argumentNotifierAXI_17_ARVALID,
	sync_argumentNotifierAXI_17_ARADDR,
	sync_argumentNotifierAXI_17_ARLEN,
	sync_argumentNotifierAXI_17_ARSIZE,
	sync_argumentNotifierAXI_17_ARBURST,
	sync_argumentNotifierAXI_17_ARLOCK,
	sync_argumentNotifierAXI_17_ARCACHE,
	sync_argumentNotifierAXI_17_ARPROT,
	sync_argumentNotifierAXI_17_ARQOS,
	sync_argumentNotifierAXI_17_ARREGION,
	sync_argumentNotifierAXI_17_RREADY,
	sync_argumentNotifierAXI_17_RVALID,
	sync_argumentNotifierAXI_17_RDATA,
	sync_argumentNotifierAXI_17_RRESP,
	sync_argumentNotifierAXI_17_RLAST,
	sync_argumentNotifierAXI_17_AWREADY,
	sync_argumentNotifierAXI_17_AWVALID,
	sync_argumentNotifierAXI_17_AWADDR,
	sync_argumentNotifierAXI_17_AWLEN,
	sync_argumentNotifierAXI_17_AWSIZE,
	sync_argumentNotifierAXI_17_AWBURST,
	sync_argumentNotifierAXI_17_AWLOCK,
	sync_argumentNotifierAXI_17_AWCACHE,
	sync_argumentNotifierAXI_17_AWPROT,
	sync_argumentNotifierAXI_17_AWQOS,
	sync_argumentNotifierAXI_17_AWREGION,
	sync_argumentNotifierAXI_17_WREADY,
	sync_argumentNotifierAXI_17_WVALID,
	sync_argumentNotifierAXI_17_WDATA,
	sync_argumentNotifierAXI_17_WSTRB,
	sync_argumentNotifierAXI_17_WLAST,
	sync_argumentNotifierAXI_17_BREADY,
	sync_argumentNotifierAXI_17_BVALID,
	sync_argumentNotifierAXI_17_BRESP,
	sync_argumentNotifierAXI_18_ARREADY,
	sync_argumentNotifierAXI_18_ARVALID,
	sync_argumentNotifierAXI_18_ARADDR,
	sync_argumentNotifierAXI_18_ARLEN,
	sync_argumentNotifierAXI_18_ARSIZE,
	sync_argumentNotifierAXI_18_ARBURST,
	sync_argumentNotifierAXI_18_ARLOCK,
	sync_argumentNotifierAXI_18_ARCACHE,
	sync_argumentNotifierAXI_18_ARPROT,
	sync_argumentNotifierAXI_18_ARQOS,
	sync_argumentNotifierAXI_18_ARREGION,
	sync_argumentNotifierAXI_18_RREADY,
	sync_argumentNotifierAXI_18_RVALID,
	sync_argumentNotifierAXI_18_RDATA,
	sync_argumentNotifierAXI_18_RRESP,
	sync_argumentNotifierAXI_18_RLAST,
	sync_argumentNotifierAXI_18_AWREADY,
	sync_argumentNotifierAXI_18_AWVALID,
	sync_argumentNotifierAXI_18_AWADDR,
	sync_argumentNotifierAXI_18_AWLEN,
	sync_argumentNotifierAXI_18_AWSIZE,
	sync_argumentNotifierAXI_18_AWBURST,
	sync_argumentNotifierAXI_18_AWLOCK,
	sync_argumentNotifierAXI_18_AWCACHE,
	sync_argumentNotifierAXI_18_AWPROT,
	sync_argumentNotifierAXI_18_AWQOS,
	sync_argumentNotifierAXI_18_AWREGION,
	sync_argumentNotifierAXI_18_WREADY,
	sync_argumentNotifierAXI_18_WVALID,
	sync_argumentNotifierAXI_18_WDATA,
	sync_argumentNotifierAXI_18_WSTRB,
	sync_argumentNotifierAXI_18_WLAST,
	sync_argumentNotifierAXI_18_BREADY,
	sync_argumentNotifierAXI_18_BVALID,
	sync_argumentNotifierAXI_18_BRESP,
	sync_argumentNotifierAXI_19_ARREADY,
	sync_argumentNotifierAXI_19_ARVALID,
	sync_argumentNotifierAXI_19_ARADDR,
	sync_argumentNotifierAXI_19_ARLEN,
	sync_argumentNotifierAXI_19_ARSIZE,
	sync_argumentNotifierAXI_19_ARBURST,
	sync_argumentNotifierAXI_19_ARLOCK,
	sync_argumentNotifierAXI_19_ARCACHE,
	sync_argumentNotifierAXI_19_ARPROT,
	sync_argumentNotifierAXI_19_ARQOS,
	sync_argumentNotifierAXI_19_ARREGION,
	sync_argumentNotifierAXI_19_RREADY,
	sync_argumentNotifierAXI_19_RVALID,
	sync_argumentNotifierAXI_19_RDATA,
	sync_argumentNotifierAXI_19_RRESP,
	sync_argumentNotifierAXI_19_RLAST,
	sync_argumentNotifierAXI_19_AWREADY,
	sync_argumentNotifierAXI_19_AWVALID,
	sync_argumentNotifierAXI_19_AWADDR,
	sync_argumentNotifierAXI_19_AWLEN,
	sync_argumentNotifierAXI_19_AWSIZE,
	sync_argumentNotifierAXI_19_AWBURST,
	sync_argumentNotifierAXI_19_AWLOCK,
	sync_argumentNotifierAXI_19_AWCACHE,
	sync_argumentNotifierAXI_19_AWPROT,
	sync_argumentNotifierAXI_19_AWQOS,
	sync_argumentNotifierAXI_19_AWREGION,
	sync_argumentNotifierAXI_19_WREADY,
	sync_argumentNotifierAXI_19_WVALID,
	sync_argumentNotifierAXI_19_WDATA,
	sync_argumentNotifierAXI_19_WSTRB,
	sync_argumentNotifierAXI_19_WLAST,
	sync_argumentNotifierAXI_19_BREADY,
	sync_argumentNotifierAXI_19_BVALID,
	sync_argumentNotifierAXI_19_BRESP,
	sync_argumentNotifierAXI_20_ARREADY,
	sync_argumentNotifierAXI_20_ARVALID,
	sync_argumentNotifierAXI_20_ARADDR,
	sync_argumentNotifierAXI_20_ARLEN,
	sync_argumentNotifierAXI_20_ARSIZE,
	sync_argumentNotifierAXI_20_ARBURST,
	sync_argumentNotifierAXI_20_ARLOCK,
	sync_argumentNotifierAXI_20_ARCACHE,
	sync_argumentNotifierAXI_20_ARPROT,
	sync_argumentNotifierAXI_20_ARQOS,
	sync_argumentNotifierAXI_20_ARREGION,
	sync_argumentNotifierAXI_20_RREADY,
	sync_argumentNotifierAXI_20_RVALID,
	sync_argumentNotifierAXI_20_RDATA,
	sync_argumentNotifierAXI_20_RRESP,
	sync_argumentNotifierAXI_20_RLAST,
	sync_argumentNotifierAXI_20_AWREADY,
	sync_argumentNotifierAXI_20_AWVALID,
	sync_argumentNotifierAXI_20_AWADDR,
	sync_argumentNotifierAXI_20_AWLEN,
	sync_argumentNotifierAXI_20_AWSIZE,
	sync_argumentNotifierAXI_20_AWBURST,
	sync_argumentNotifierAXI_20_AWLOCK,
	sync_argumentNotifierAXI_20_AWCACHE,
	sync_argumentNotifierAXI_20_AWPROT,
	sync_argumentNotifierAXI_20_AWQOS,
	sync_argumentNotifierAXI_20_AWREGION,
	sync_argumentNotifierAXI_20_WREADY,
	sync_argumentNotifierAXI_20_WVALID,
	sync_argumentNotifierAXI_20_WDATA,
	sync_argumentNotifierAXI_20_WSTRB,
	sync_argumentNotifierAXI_20_WLAST,
	sync_argumentNotifierAXI_20_BREADY,
	sync_argumentNotifierAXI_20_BVALID,
	sync_argumentNotifierAXI_20_BRESP,
	sync_argumentNotifierAXI_21_ARREADY,
	sync_argumentNotifierAXI_21_ARVALID,
	sync_argumentNotifierAXI_21_ARADDR,
	sync_argumentNotifierAXI_21_ARLEN,
	sync_argumentNotifierAXI_21_ARSIZE,
	sync_argumentNotifierAXI_21_ARBURST,
	sync_argumentNotifierAXI_21_ARLOCK,
	sync_argumentNotifierAXI_21_ARCACHE,
	sync_argumentNotifierAXI_21_ARPROT,
	sync_argumentNotifierAXI_21_ARQOS,
	sync_argumentNotifierAXI_21_ARREGION,
	sync_argumentNotifierAXI_21_RREADY,
	sync_argumentNotifierAXI_21_RVALID,
	sync_argumentNotifierAXI_21_RDATA,
	sync_argumentNotifierAXI_21_RRESP,
	sync_argumentNotifierAXI_21_RLAST,
	sync_argumentNotifierAXI_21_AWREADY,
	sync_argumentNotifierAXI_21_AWVALID,
	sync_argumentNotifierAXI_21_AWADDR,
	sync_argumentNotifierAXI_21_AWLEN,
	sync_argumentNotifierAXI_21_AWSIZE,
	sync_argumentNotifierAXI_21_AWBURST,
	sync_argumentNotifierAXI_21_AWLOCK,
	sync_argumentNotifierAXI_21_AWCACHE,
	sync_argumentNotifierAXI_21_AWPROT,
	sync_argumentNotifierAXI_21_AWQOS,
	sync_argumentNotifierAXI_21_AWREGION,
	sync_argumentNotifierAXI_21_WREADY,
	sync_argumentNotifierAXI_21_WVALID,
	sync_argumentNotifierAXI_21_WDATA,
	sync_argumentNotifierAXI_21_WSTRB,
	sync_argumentNotifierAXI_21_WLAST,
	sync_argumentNotifierAXI_21_BREADY,
	sync_argumentNotifierAXI_21_BVALID,
	sync_argumentNotifierAXI_21_BRESP,
	sync_argumentNotifierAXI_22_ARREADY,
	sync_argumentNotifierAXI_22_ARVALID,
	sync_argumentNotifierAXI_22_ARADDR,
	sync_argumentNotifierAXI_22_ARLEN,
	sync_argumentNotifierAXI_22_ARSIZE,
	sync_argumentNotifierAXI_22_ARBURST,
	sync_argumentNotifierAXI_22_ARLOCK,
	sync_argumentNotifierAXI_22_ARCACHE,
	sync_argumentNotifierAXI_22_ARPROT,
	sync_argumentNotifierAXI_22_ARQOS,
	sync_argumentNotifierAXI_22_ARREGION,
	sync_argumentNotifierAXI_22_RREADY,
	sync_argumentNotifierAXI_22_RVALID,
	sync_argumentNotifierAXI_22_RDATA,
	sync_argumentNotifierAXI_22_RRESP,
	sync_argumentNotifierAXI_22_RLAST,
	sync_argumentNotifierAXI_22_AWREADY,
	sync_argumentNotifierAXI_22_AWVALID,
	sync_argumentNotifierAXI_22_AWADDR,
	sync_argumentNotifierAXI_22_AWLEN,
	sync_argumentNotifierAXI_22_AWSIZE,
	sync_argumentNotifierAXI_22_AWBURST,
	sync_argumentNotifierAXI_22_AWLOCK,
	sync_argumentNotifierAXI_22_AWCACHE,
	sync_argumentNotifierAXI_22_AWPROT,
	sync_argumentNotifierAXI_22_AWQOS,
	sync_argumentNotifierAXI_22_AWREGION,
	sync_argumentNotifierAXI_22_WREADY,
	sync_argumentNotifierAXI_22_WVALID,
	sync_argumentNotifierAXI_22_WDATA,
	sync_argumentNotifierAXI_22_WSTRB,
	sync_argumentNotifierAXI_22_WLAST,
	sync_argumentNotifierAXI_22_BREADY,
	sync_argumentNotifierAXI_22_BVALID,
	sync_argumentNotifierAXI_22_BRESP,
	sync_argumentNotifierAXI_23_ARREADY,
	sync_argumentNotifierAXI_23_ARVALID,
	sync_argumentNotifierAXI_23_ARADDR,
	sync_argumentNotifierAXI_23_ARLEN,
	sync_argumentNotifierAXI_23_ARSIZE,
	sync_argumentNotifierAXI_23_ARBURST,
	sync_argumentNotifierAXI_23_ARLOCK,
	sync_argumentNotifierAXI_23_ARCACHE,
	sync_argumentNotifierAXI_23_ARPROT,
	sync_argumentNotifierAXI_23_ARQOS,
	sync_argumentNotifierAXI_23_ARREGION,
	sync_argumentNotifierAXI_23_RREADY,
	sync_argumentNotifierAXI_23_RVALID,
	sync_argumentNotifierAXI_23_RDATA,
	sync_argumentNotifierAXI_23_RRESP,
	sync_argumentNotifierAXI_23_RLAST,
	sync_argumentNotifierAXI_23_AWREADY,
	sync_argumentNotifierAXI_23_AWVALID,
	sync_argumentNotifierAXI_23_AWADDR,
	sync_argumentNotifierAXI_23_AWLEN,
	sync_argumentNotifierAXI_23_AWSIZE,
	sync_argumentNotifierAXI_23_AWBURST,
	sync_argumentNotifierAXI_23_AWLOCK,
	sync_argumentNotifierAXI_23_AWCACHE,
	sync_argumentNotifierAXI_23_AWPROT,
	sync_argumentNotifierAXI_23_AWQOS,
	sync_argumentNotifierAXI_23_AWREGION,
	sync_argumentNotifierAXI_23_WREADY,
	sync_argumentNotifierAXI_23_WVALID,
	sync_argumentNotifierAXI_23_WDATA,
	sync_argumentNotifierAXI_23_WSTRB,
	sync_argumentNotifierAXI_23_WLAST,
	sync_argumentNotifierAXI_23_BREADY,
	sync_argumentNotifierAXI_23_BVALID,
	sync_argumentNotifierAXI_23_BRESP,
	sync_argumentNotifierAXI_24_ARREADY,
	sync_argumentNotifierAXI_24_ARVALID,
	sync_argumentNotifierAXI_24_ARADDR,
	sync_argumentNotifierAXI_24_ARLEN,
	sync_argumentNotifierAXI_24_ARSIZE,
	sync_argumentNotifierAXI_24_ARBURST,
	sync_argumentNotifierAXI_24_ARLOCK,
	sync_argumentNotifierAXI_24_ARCACHE,
	sync_argumentNotifierAXI_24_ARPROT,
	sync_argumentNotifierAXI_24_ARQOS,
	sync_argumentNotifierAXI_24_ARREGION,
	sync_argumentNotifierAXI_24_RREADY,
	sync_argumentNotifierAXI_24_RVALID,
	sync_argumentNotifierAXI_24_RDATA,
	sync_argumentNotifierAXI_24_RRESP,
	sync_argumentNotifierAXI_24_RLAST,
	sync_argumentNotifierAXI_24_AWREADY,
	sync_argumentNotifierAXI_24_AWVALID,
	sync_argumentNotifierAXI_24_AWADDR,
	sync_argumentNotifierAXI_24_AWLEN,
	sync_argumentNotifierAXI_24_AWSIZE,
	sync_argumentNotifierAXI_24_AWBURST,
	sync_argumentNotifierAXI_24_AWLOCK,
	sync_argumentNotifierAXI_24_AWCACHE,
	sync_argumentNotifierAXI_24_AWPROT,
	sync_argumentNotifierAXI_24_AWQOS,
	sync_argumentNotifierAXI_24_AWREGION,
	sync_argumentNotifierAXI_24_WREADY,
	sync_argumentNotifierAXI_24_WVALID,
	sync_argumentNotifierAXI_24_WDATA,
	sync_argumentNotifierAXI_24_WSTRB,
	sync_argumentNotifierAXI_24_WLAST,
	sync_argumentNotifierAXI_24_BREADY,
	sync_argumentNotifierAXI_24_BVALID,
	sync_argumentNotifierAXI_24_BRESP,
	sync_argumentNotifierAXI_25_ARREADY,
	sync_argumentNotifierAXI_25_ARVALID,
	sync_argumentNotifierAXI_25_ARADDR,
	sync_argumentNotifierAXI_25_ARLEN,
	sync_argumentNotifierAXI_25_ARSIZE,
	sync_argumentNotifierAXI_25_ARBURST,
	sync_argumentNotifierAXI_25_ARLOCK,
	sync_argumentNotifierAXI_25_ARCACHE,
	sync_argumentNotifierAXI_25_ARPROT,
	sync_argumentNotifierAXI_25_ARQOS,
	sync_argumentNotifierAXI_25_ARREGION,
	sync_argumentNotifierAXI_25_RREADY,
	sync_argumentNotifierAXI_25_RVALID,
	sync_argumentNotifierAXI_25_RDATA,
	sync_argumentNotifierAXI_25_RRESP,
	sync_argumentNotifierAXI_25_RLAST,
	sync_argumentNotifierAXI_25_AWREADY,
	sync_argumentNotifierAXI_25_AWVALID,
	sync_argumentNotifierAXI_25_AWADDR,
	sync_argumentNotifierAXI_25_AWLEN,
	sync_argumentNotifierAXI_25_AWSIZE,
	sync_argumentNotifierAXI_25_AWBURST,
	sync_argumentNotifierAXI_25_AWLOCK,
	sync_argumentNotifierAXI_25_AWCACHE,
	sync_argumentNotifierAXI_25_AWPROT,
	sync_argumentNotifierAXI_25_AWQOS,
	sync_argumentNotifierAXI_25_AWREGION,
	sync_argumentNotifierAXI_25_WREADY,
	sync_argumentNotifierAXI_25_WVALID,
	sync_argumentNotifierAXI_25_WDATA,
	sync_argumentNotifierAXI_25_WSTRB,
	sync_argumentNotifierAXI_25_WLAST,
	sync_argumentNotifierAXI_25_BREADY,
	sync_argumentNotifierAXI_25_BVALID,
	sync_argumentNotifierAXI_25_BRESP,
	sync_argumentNotifierAXI_26_ARREADY,
	sync_argumentNotifierAXI_26_ARVALID,
	sync_argumentNotifierAXI_26_ARADDR,
	sync_argumentNotifierAXI_26_ARLEN,
	sync_argumentNotifierAXI_26_ARSIZE,
	sync_argumentNotifierAXI_26_ARBURST,
	sync_argumentNotifierAXI_26_ARLOCK,
	sync_argumentNotifierAXI_26_ARCACHE,
	sync_argumentNotifierAXI_26_ARPROT,
	sync_argumentNotifierAXI_26_ARQOS,
	sync_argumentNotifierAXI_26_ARREGION,
	sync_argumentNotifierAXI_26_RREADY,
	sync_argumentNotifierAXI_26_RVALID,
	sync_argumentNotifierAXI_26_RDATA,
	sync_argumentNotifierAXI_26_RRESP,
	sync_argumentNotifierAXI_26_RLAST,
	sync_argumentNotifierAXI_26_AWREADY,
	sync_argumentNotifierAXI_26_AWVALID,
	sync_argumentNotifierAXI_26_AWADDR,
	sync_argumentNotifierAXI_26_AWLEN,
	sync_argumentNotifierAXI_26_AWSIZE,
	sync_argumentNotifierAXI_26_AWBURST,
	sync_argumentNotifierAXI_26_AWLOCK,
	sync_argumentNotifierAXI_26_AWCACHE,
	sync_argumentNotifierAXI_26_AWPROT,
	sync_argumentNotifierAXI_26_AWQOS,
	sync_argumentNotifierAXI_26_AWREGION,
	sync_argumentNotifierAXI_26_WREADY,
	sync_argumentNotifierAXI_26_WVALID,
	sync_argumentNotifierAXI_26_WDATA,
	sync_argumentNotifierAXI_26_WSTRB,
	sync_argumentNotifierAXI_26_WLAST,
	sync_argumentNotifierAXI_26_BREADY,
	sync_argumentNotifierAXI_26_BVALID,
	sync_argumentNotifierAXI_26_BRESP,
	sync_argumentNotifierAXI_27_ARREADY,
	sync_argumentNotifierAXI_27_ARVALID,
	sync_argumentNotifierAXI_27_ARADDR,
	sync_argumentNotifierAXI_27_ARLEN,
	sync_argumentNotifierAXI_27_ARSIZE,
	sync_argumentNotifierAXI_27_ARBURST,
	sync_argumentNotifierAXI_27_ARLOCK,
	sync_argumentNotifierAXI_27_ARCACHE,
	sync_argumentNotifierAXI_27_ARPROT,
	sync_argumentNotifierAXI_27_ARQOS,
	sync_argumentNotifierAXI_27_ARREGION,
	sync_argumentNotifierAXI_27_RREADY,
	sync_argumentNotifierAXI_27_RVALID,
	sync_argumentNotifierAXI_27_RDATA,
	sync_argumentNotifierAXI_27_RRESP,
	sync_argumentNotifierAXI_27_RLAST,
	sync_argumentNotifierAXI_27_AWREADY,
	sync_argumentNotifierAXI_27_AWVALID,
	sync_argumentNotifierAXI_27_AWADDR,
	sync_argumentNotifierAXI_27_AWLEN,
	sync_argumentNotifierAXI_27_AWSIZE,
	sync_argumentNotifierAXI_27_AWBURST,
	sync_argumentNotifierAXI_27_AWLOCK,
	sync_argumentNotifierAXI_27_AWCACHE,
	sync_argumentNotifierAXI_27_AWPROT,
	sync_argumentNotifierAXI_27_AWQOS,
	sync_argumentNotifierAXI_27_AWREGION,
	sync_argumentNotifierAXI_27_WREADY,
	sync_argumentNotifierAXI_27_WVALID,
	sync_argumentNotifierAXI_27_WDATA,
	sync_argumentNotifierAXI_27_WSTRB,
	sync_argumentNotifierAXI_27_WLAST,
	sync_argumentNotifierAXI_27_BREADY,
	sync_argumentNotifierAXI_27_BVALID,
	sync_argumentNotifierAXI_27_BRESP,
	sync_argumentNotifierAXI_28_ARREADY,
	sync_argumentNotifierAXI_28_ARVALID,
	sync_argumentNotifierAXI_28_ARADDR,
	sync_argumentNotifierAXI_28_ARLEN,
	sync_argumentNotifierAXI_28_ARSIZE,
	sync_argumentNotifierAXI_28_ARBURST,
	sync_argumentNotifierAXI_28_ARLOCK,
	sync_argumentNotifierAXI_28_ARCACHE,
	sync_argumentNotifierAXI_28_ARPROT,
	sync_argumentNotifierAXI_28_ARQOS,
	sync_argumentNotifierAXI_28_ARREGION,
	sync_argumentNotifierAXI_28_RREADY,
	sync_argumentNotifierAXI_28_RVALID,
	sync_argumentNotifierAXI_28_RDATA,
	sync_argumentNotifierAXI_28_RRESP,
	sync_argumentNotifierAXI_28_RLAST,
	sync_argumentNotifierAXI_28_AWREADY,
	sync_argumentNotifierAXI_28_AWVALID,
	sync_argumentNotifierAXI_28_AWADDR,
	sync_argumentNotifierAXI_28_AWLEN,
	sync_argumentNotifierAXI_28_AWSIZE,
	sync_argumentNotifierAXI_28_AWBURST,
	sync_argumentNotifierAXI_28_AWLOCK,
	sync_argumentNotifierAXI_28_AWCACHE,
	sync_argumentNotifierAXI_28_AWPROT,
	sync_argumentNotifierAXI_28_AWQOS,
	sync_argumentNotifierAXI_28_AWREGION,
	sync_argumentNotifierAXI_28_WREADY,
	sync_argumentNotifierAXI_28_WVALID,
	sync_argumentNotifierAXI_28_WDATA,
	sync_argumentNotifierAXI_28_WSTRB,
	sync_argumentNotifierAXI_28_WLAST,
	sync_argumentNotifierAXI_28_BREADY,
	sync_argumentNotifierAXI_28_BVALID,
	sync_argumentNotifierAXI_28_BRESP,
	sync_argumentNotifierAXI_29_ARREADY,
	sync_argumentNotifierAXI_29_ARVALID,
	sync_argumentNotifierAXI_29_ARADDR,
	sync_argumentNotifierAXI_29_ARLEN,
	sync_argumentNotifierAXI_29_ARSIZE,
	sync_argumentNotifierAXI_29_ARBURST,
	sync_argumentNotifierAXI_29_ARLOCK,
	sync_argumentNotifierAXI_29_ARCACHE,
	sync_argumentNotifierAXI_29_ARPROT,
	sync_argumentNotifierAXI_29_ARQOS,
	sync_argumentNotifierAXI_29_ARREGION,
	sync_argumentNotifierAXI_29_RREADY,
	sync_argumentNotifierAXI_29_RVALID,
	sync_argumentNotifierAXI_29_RDATA,
	sync_argumentNotifierAXI_29_RRESP,
	sync_argumentNotifierAXI_29_RLAST,
	sync_argumentNotifierAXI_29_AWREADY,
	sync_argumentNotifierAXI_29_AWVALID,
	sync_argumentNotifierAXI_29_AWADDR,
	sync_argumentNotifierAXI_29_AWLEN,
	sync_argumentNotifierAXI_29_AWSIZE,
	sync_argumentNotifierAXI_29_AWBURST,
	sync_argumentNotifierAXI_29_AWLOCK,
	sync_argumentNotifierAXI_29_AWCACHE,
	sync_argumentNotifierAXI_29_AWPROT,
	sync_argumentNotifierAXI_29_AWQOS,
	sync_argumentNotifierAXI_29_AWREGION,
	sync_argumentNotifierAXI_29_WREADY,
	sync_argumentNotifierAXI_29_WVALID,
	sync_argumentNotifierAXI_29_WDATA,
	sync_argumentNotifierAXI_29_WSTRB,
	sync_argumentNotifierAXI_29_WLAST,
	sync_argumentNotifierAXI_29_BREADY,
	sync_argumentNotifierAXI_29_BVALID,
	sync_argumentNotifierAXI_29_BRESP,
	sync_argumentNotifierAXI_30_ARREADY,
	sync_argumentNotifierAXI_30_ARVALID,
	sync_argumentNotifierAXI_30_ARADDR,
	sync_argumentNotifierAXI_30_ARLEN,
	sync_argumentNotifierAXI_30_ARSIZE,
	sync_argumentNotifierAXI_30_ARBURST,
	sync_argumentNotifierAXI_30_ARLOCK,
	sync_argumentNotifierAXI_30_ARCACHE,
	sync_argumentNotifierAXI_30_ARPROT,
	sync_argumentNotifierAXI_30_ARQOS,
	sync_argumentNotifierAXI_30_ARREGION,
	sync_argumentNotifierAXI_30_RREADY,
	sync_argumentNotifierAXI_30_RVALID,
	sync_argumentNotifierAXI_30_RDATA,
	sync_argumentNotifierAXI_30_RRESP,
	sync_argumentNotifierAXI_30_RLAST,
	sync_argumentNotifierAXI_30_AWREADY,
	sync_argumentNotifierAXI_30_AWVALID,
	sync_argumentNotifierAXI_30_AWADDR,
	sync_argumentNotifierAXI_30_AWLEN,
	sync_argumentNotifierAXI_30_AWSIZE,
	sync_argumentNotifierAXI_30_AWBURST,
	sync_argumentNotifierAXI_30_AWLOCK,
	sync_argumentNotifierAXI_30_AWCACHE,
	sync_argumentNotifierAXI_30_AWPROT,
	sync_argumentNotifierAXI_30_AWQOS,
	sync_argumentNotifierAXI_30_AWREGION,
	sync_argumentNotifierAXI_30_WREADY,
	sync_argumentNotifierAXI_30_WVALID,
	sync_argumentNotifierAXI_30_WDATA,
	sync_argumentNotifierAXI_30_WSTRB,
	sync_argumentNotifierAXI_30_WLAST,
	sync_argumentNotifierAXI_30_BREADY,
	sync_argumentNotifierAXI_30_BVALID,
	sync_argumentNotifierAXI_30_BRESP,
	sync_argumentNotifierAXI_31_ARREADY,
	sync_argumentNotifierAXI_31_ARVALID,
	sync_argumentNotifierAXI_31_ARADDR,
	sync_argumentNotifierAXI_31_ARLEN,
	sync_argumentNotifierAXI_31_ARSIZE,
	sync_argumentNotifierAXI_31_ARBURST,
	sync_argumentNotifierAXI_31_ARLOCK,
	sync_argumentNotifierAXI_31_ARCACHE,
	sync_argumentNotifierAXI_31_ARPROT,
	sync_argumentNotifierAXI_31_ARQOS,
	sync_argumentNotifierAXI_31_ARREGION,
	sync_argumentNotifierAXI_31_RREADY,
	sync_argumentNotifierAXI_31_RVALID,
	sync_argumentNotifierAXI_31_RDATA,
	sync_argumentNotifierAXI_31_RRESP,
	sync_argumentNotifierAXI_31_RLAST,
	sync_argumentNotifierAXI_31_AWREADY,
	sync_argumentNotifierAXI_31_AWVALID,
	sync_argumentNotifierAXI_31_AWADDR,
	sync_argumentNotifierAXI_31_AWLEN,
	sync_argumentNotifierAXI_31_AWSIZE,
	sync_argumentNotifierAXI_31_AWBURST,
	sync_argumentNotifierAXI_31_AWLOCK,
	sync_argumentNotifierAXI_31_AWCACHE,
	sync_argumentNotifierAXI_31_AWPROT,
	sync_argumentNotifierAXI_31_AWQOS,
	sync_argumentNotifierAXI_31_AWREGION,
	sync_argumentNotifierAXI_31_WREADY,
	sync_argumentNotifierAXI_31_WVALID,
	sync_argumentNotifierAXI_31_WDATA,
	sync_argumentNotifierAXI_31_WSTRB,
	sync_argumentNotifierAXI_31_WLAST,
	sync_argumentNotifierAXI_31_BREADY,
	sync_argumentNotifierAXI_31_BVALID,
	sync_argumentNotifierAXI_31_BRESP
);
	input clock;
	input reset;
	output wire s_axil_mgmt_hardcilk_ARREADY;
	input s_axil_mgmt_hardcilk_ARVALID;
	input [11:0] s_axil_mgmt_hardcilk_ARADDR;
	input [2:0] s_axil_mgmt_hardcilk_ARPROT;
	input s_axil_mgmt_hardcilk_RREADY;
	output wire s_axil_mgmt_hardcilk_RVALID;
	output wire [63:0] s_axil_mgmt_hardcilk_RDATA;
	output wire [1:0] s_axil_mgmt_hardcilk_RRESP;
	output wire s_axil_mgmt_hardcilk_AWREADY;
	input s_axil_mgmt_hardcilk_AWVALID;
	input [11:0] s_axil_mgmt_hardcilk_AWADDR;
	input [2:0] s_axil_mgmt_hardcilk_AWPROT;
	output wire s_axil_mgmt_hardcilk_WREADY;
	input s_axil_mgmt_hardcilk_WVALID;
	input [63:0] s_axil_mgmt_hardcilk_WDATA;
	input [7:0] s_axil_mgmt_hardcilk_WSTRB;
	input s_axil_mgmt_hardcilk_BREADY;
	output wire s_axil_mgmt_hardcilk_BVALID;
	output wire [1:0] s_axil_mgmt_hardcilk_BRESP;
	input qsort_0_m_axi_gmem_ARREADY;
	output wire qsort_0_m_axi_gmem_ARVALID;
	output wire qsort_0_m_axi_gmem_ARID;
	output wire [63:0] qsort_0_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_0_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_0_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_0_m_axi_gmem_ARBURST;
	output wire qsort_0_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_0_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_0_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_0_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_0_m_axi_gmem_ARREGION;
	output wire qsort_0_m_axi_gmem_ARUSER;
	output wire qsort_0_m_axi_gmem_RREADY;
	input qsort_0_m_axi_gmem_RVALID;
	input qsort_0_m_axi_gmem_RID;
	input [63:0] qsort_0_m_axi_gmem_RDATA;
	input [1:0] qsort_0_m_axi_gmem_RRESP;
	input qsort_0_m_axi_gmem_RLAST;
	input qsort_0_m_axi_gmem_RUSER;
	input qsort_0_m_axi_gmem_AWREADY;
	output wire qsort_0_m_axi_gmem_AWVALID;
	output wire qsort_0_m_axi_gmem_AWID;
	output wire [63:0] qsort_0_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_0_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_0_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_0_m_axi_gmem_AWBURST;
	output wire qsort_0_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_0_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_0_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_0_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_0_m_axi_gmem_AWREGION;
	output wire qsort_0_m_axi_gmem_AWUSER;
	input qsort_0_m_axi_gmem_WREADY;
	output wire qsort_0_m_axi_gmem_WVALID;
	output wire [63:0] qsort_0_m_axi_gmem_WDATA;
	output wire [7:0] qsort_0_m_axi_gmem_WSTRB;
	output wire qsort_0_m_axi_gmem_WLAST;
	output wire qsort_0_m_axi_gmem_WUSER;
	output wire qsort_0_m_axi_gmem_BREADY;
	input qsort_0_m_axi_gmem_BVALID;
	input qsort_0_m_axi_gmem_BID;
	input [1:0] qsort_0_m_axi_gmem_BRESP;
	input qsort_0_m_axi_gmem_BUSER;
	output wire qsort_0_s_axi_control_ARREADY;
	input qsort_0_s_axi_control_ARVALID;
	input [5:0] qsort_0_s_axi_control_ARADDR;
	input qsort_0_s_axi_control_RREADY;
	output wire qsort_0_s_axi_control_RVALID;
	output wire [31:0] qsort_0_s_axi_control_RDATA;
	output wire [1:0] qsort_0_s_axi_control_RRESP;
	output wire qsort_0_s_axi_control_AWREADY;
	input qsort_0_s_axi_control_AWVALID;
	input [5:0] qsort_0_s_axi_control_AWADDR;
	output wire qsort_0_s_axi_control_WREADY;
	input qsort_0_s_axi_control_WVALID;
	input [31:0] qsort_0_s_axi_control_WDATA;
	input [3:0] qsort_0_s_axi_control_WSTRB;
	input qsort_0_s_axi_control_BREADY;
	output wire qsort_0_s_axi_control_BVALID;
	output wire [1:0] qsort_0_s_axi_control_BRESP;
	input qsort_1_m_axi_gmem_ARREADY;
	output wire qsort_1_m_axi_gmem_ARVALID;
	output wire qsort_1_m_axi_gmem_ARID;
	output wire [63:0] qsort_1_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_1_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_1_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_1_m_axi_gmem_ARBURST;
	output wire qsort_1_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_1_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_1_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_1_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_1_m_axi_gmem_ARREGION;
	output wire qsort_1_m_axi_gmem_ARUSER;
	output wire qsort_1_m_axi_gmem_RREADY;
	input qsort_1_m_axi_gmem_RVALID;
	input qsort_1_m_axi_gmem_RID;
	input [63:0] qsort_1_m_axi_gmem_RDATA;
	input [1:0] qsort_1_m_axi_gmem_RRESP;
	input qsort_1_m_axi_gmem_RLAST;
	input qsort_1_m_axi_gmem_RUSER;
	input qsort_1_m_axi_gmem_AWREADY;
	output wire qsort_1_m_axi_gmem_AWVALID;
	output wire qsort_1_m_axi_gmem_AWID;
	output wire [63:0] qsort_1_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_1_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_1_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_1_m_axi_gmem_AWBURST;
	output wire qsort_1_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_1_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_1_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_1_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_1_m_axi_gmem_AWREGION;
	output wire qsort_1_m_axi_gmem_AWUSER;
	input qsort_1_m_axi_gmem_WREADY;
	output wire qsort_1_m_axi_gmem_WVALID;
	output wire [63:0] qsort_1_m_axi_gmem_WDATA;
	output wire [7:0] qsort_1_m_axi_gmem_WSTRB;
	output wire qsort_1_m_axi_gmem_WLAST;
	output wire qsort_1_m_axi_gmem_WUSER;
	output wire qsort_1_m_axi_gmem_BREADY;
	input qsort_1_m_axi_gmem_BVALID;
	input qsort_1_m_axi_gmem_BID;
	input [1:0] qsort_1_m_axi_gmem_BRESP;
	input qsort_1_m_axi_gmem_BUSER;
	output wire qsort_1_s_axi_control_ARREADY;
	input qsort_1_s_axi_control_ARVALID;
	input [5:0] qsort_1_s_axi_control_ARADDR;
	input qsort_1_s_axi_control_RREADY;
	output wire qsort_1_s_axi_control_RVALID;
	output wire [31:0] qsort_1_s_axi_control_RDATA;
	output wire [1:0] qsort_1_s_axi_control_RRESP;
	output wire qsort_1_s_axi_control_AWREADY;
	input qsort_1_s_axi_control_AWVALID;
	input [5:0] qsort_1_s_axi_control_AWADDR;
	output wire qsort_1_s_axi_control_WREADY;
	input qsort_1_s_axi_control_WVALID;
	input [31:0] qsort_1_s_axi_control_WDATA;
	input [3:0] qsort_1_s_axi_control_WSTRB;
	input qsort_1_s_axi_control_BREADY;
	output wire qsort_1_s_axi_control_BVALID;
	output wire [1:0] qsort_1_s_axi_control_BRESP;
	input qsort_2_m_axi_gmem_ARREADY;
	output wire qsort_2_m_axi_gmem_ARVALID;
	output wire qsort_2_m_axi_gmem_ARID;
	output wire [63:0] qsort_2_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_2_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_2_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_2_m_axi_gmem_ARBURST;
	output wire qsort_2_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_2_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_2_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_2_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_2_m_axi_gmem_ARREGION;
	output wire qsort_2_m_axi_gmem_ARUSER;
	output wire qsort_2_m_axi_gmem_RREADY;
	input qsort_2_m_axi_gmem_RVALID;
	input qsort_2_m_axi_gmem_RID;
	input [63:0] qsort_2_m_axi_gmem_RDATA;
	input [1:0] qsort_2_m_axi_gmem_RRESP;
	input qsort_2_m_axi_gmem_RLAST;
	input qsort_2_m_axi_gmem_RUSER;
	input qsort_2_m_axi_gmem_AWREADY;
	output wire qsort_2_m_axi_gmem_AWVALID;
	output wire qsort_2_m_axi_gmem_AWID;
	output wire [63:0] qsort_2_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_2_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_2_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_2_m_axi_gmem_AWBURST;
	output wire qsort_2_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_2_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_2_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_2_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_2_m_axi_gmem_AWREGION;
	output wire qsort_2_m_axi_gmem_AWUSER;
	input qsort_2_m_axi_gmem_WREADY;
	output wire qsort_2_m_axi_gmem_WVALID;
	output wire [63:0] qsort_2_m_axi_gmem_WDATA;
	output wire [7:0] qsort_2_m_axi_gmem_WSTRB;
	output wire qsort_2_m_axi_gmem_WLAST;
	output wire qsort_2_m_axi_gmem_WUSER;
	output wire qsort_2_m_axi_gmem_BREADY;
	input qsort_2_m_axi_gmem_BVALID;
	input qsort_2_m_axi_gmem_BID;
	input [1:0] qsort_2_m_axi_gmem_BRESP;
	input qsort_2_m_axi_gmem_BUSER;
	output wire qsort_2_s_axi_control_ARREADY;
	input qsort_2_s_axi_control_ARVALID;
	input [5:0] qsort_2_s_axi_control_ARADDR;
	input qsort_2_s_axi_control_RREADY;
	output wire qsort_2_s_axi_control_RVALID;
	output wire [31:0] qsort_2_s_axi_control_RDATA;
	output wire [1:0] qsort_2_s_axi_control_RRESP;
	output wire qsort_2_s_axi_control_AWREADY;
	input qsort_2_s_axi_control_AWVALID;
	input [5:0] qsort_2_s_axi_control_AWADDR;
	output wire qsort_2_s_axi_control_WREADY;
	input qsort_2_s_axi_control_WVALID;
	input [31:0] qsort_2_s_axi_control_WDATA;
	input [3:0] qsort_2_s_axi_control_WSTRB;
	input qsort_2_s_axi_control_BREADY;
	output wire qsort_2_s_axi_control_BVALID;
	output wire [1:0] qsort_2_s_axi_control_BRESP;
	input qsort_3_m_axi_gmem_ARREADY;
	output wire qsort_3_m_axi_gmem_ARVALID;
	output wire qsort_3_m_axi_gmem_ARID;
	output wire [63:0] qsort_3_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_3_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_3_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_3_m_axi_gmem_ARBURST;
	output wire qsort_3_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_3_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_3_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_3_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_3_m_axi_gmem_ARREGION;
	output wire qsort_3_m_axi_gmem_ARUSER;
	output wire qsort_3_m_axi_gmem_RREADY;
	input qsort_3_m_axi_gmem_RVALID;
	input qsort_3_m_axi_gmem_RID;
	input [63:0] qsort_3_m_axi_gmem_RDATA;
	input [1:0] qsort_3_m_axi_gmem_RRESP;
	input qsort_3_m_axi_gmem_RLAST;
	input qsort_3_m_axi_gmem_RUSER;
	input qsort_3_m_axi_gmem_AWREADY;
	output wire qsort_3_m_axi_gmem_AWVALID;
	output wire qsort_3_m_axi_gmem_AWID;
	output wire [63:0] qsort_3_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_3_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_3_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_3_m_axi_gmem_AWBURST;
	output wire qsort_3_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_3_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_3_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_3_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_3_m_axi_gmem_AWREGION;
	output wire qsort_3_m_axi_gmem_AWUSER;
	input qsort_3_m_axi_gmem_WREADY;
	output wire qsort_3_m_axi_gmem_WVALID;
	output wire [63:0] qsort_3_m_axi_gmem_WDATA;
	output wire [7:0] qsort_3_m_axi_gmem_WSTRB;
	output wire qsort_3_m_axi_gmem_WLAST;
	output wire qsort_3_m_axi_gmem_WUSER;
	output wire qsort_3_m_axi_gmem_BREADY;
	input qsort_3_m_axi_gmem_BVALID;
	input qsort_3_m_axi_gmem_BID;
	input [1:0] qsort_3_m_axi_gmem_BRESP;
	input qsort_3_m_axi_gmem_BUSER;
	output wire qsort_3_s_axi_control_ARREADY;
	input qsort_3_s_axi_control_ARVALID;
	input [5:0] qsort_3_s_axi_control_ARADDR;
	input qsort_3_s_axi_control_RREADY;
	output wire qsort_3_s_axi_control_RVALID;
	output wire [31:0] qsort_3_s_axi_control_RDATA;
	output wire [1:0] qsort_3_s_axi_control_RRESP;
	output wire qsort_3_s_axi_control_AWREADY;
	input qsort_3_s_axi_control_AWVALID;
	input [5:0] qsort_3_s_axi_control_AWADDR;
	output wire qsort_3_s_axi_control_WREADY;
	input qsort_3_s_axi_control_WVALID;
	input [31:0] qsort_3_s_axi_control_WDATA;
	input [3:0] qsort_3_s_axi_control_WSTRB;
	input qsort_3_s_axi_control_BREADY;
	output wire qsort_3_s_axi_control_BVALID;
	output wire [1:0] qsort_3_s_axi_control_BRESP;
	input qsort_4_m_axi_gmem_ARREADY;
	output wire qsort_4_m_axi_gmem_ARVALID;
	output wire qsort_4_m_axi_gmem_ARID;
	output wire [63:0] qsort_4_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_4_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_4_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_4_m_axi_gmem_ARBURST;
	output wire qsort_4_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_4_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_4_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_4_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_4_m_axi_gmem_ARREGION;
	output wire qsort_4_m_axi_gmem_ARUSER;
	output wire qsort_4_m_axi_gmem_RREADY;
	input qsort_4_m_axi_gmem_RVALID;
	input qsort_4_m_axi_gmem_RID;
	input [63:0] qsort_4_m_axi_gmem_RDATA;
	input [1:0] qsort_4_m_axi_gmem_RRESP;
	input qsort_4_m_axi_gmem_RLAST;
	input qsort_4_m_axi_gmem_RUSER;
	input qsort_4_m_axi_gmem_AWREADY;
	output wire qsort_4_m_axi_gmem_AWVALID;
	output wire qsort_4_m_axi_gmem_AWID;
	output wire [63:0] qsort_4_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_4_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_4_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_4_m_axi_gmem_AWBURST;
	output wire qsort_4_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_4_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_4_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_4_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_4_m_axi_gmem_AWREGION;
	output wire qsort_4_m_axi_gmem_AWUSER;
	input qsort_4_m_axi_gmem_WREADY;
	output wire qsort_4_m_axi_gmem_WVALID;
	output wire [63:0] qsort_4_m_axi_gmem_WDATA;
	output wire [7:0] qsort_4_m_axi_gmem_WSTRB;
	output wire qsort_4_m_axi_gmem_WLAST;
	output wire qsort_4_m_axi_gmem_WUSER;
	output wire qsort_4_m_axi_gmem_BREADY;
	input qsort_4_m_axi_gmem_BVALID;
	input qsort_4_m_axi_gmem_BID;
	input [1:0] qsort_4_m_axi_gmem_BRESP;
	input qsort_4_m_axi_gmem_BUSER;
	output wire qsort_4_s_axi_control_ARREADY;
	input qsort_4_s_axi_control_ARVALID;
	input [5:0] qsort_4_s_axi_control_ARADDR;
	input qsort_4_s_axi_control_RREADY;
	output wire qsort_4_s_axi_control_RVALID;
	output wire [31:0] qsort_4_s_axi_control_RDATA;
	output wire [1:0] qsort_4_s_axi_control_RRESP;
	output wire qsort_4_s_axi_control_AWREADY;
	input qsort_4_s_axi_control_AWVALID;
	input [5:0] qsort_4_s_axi_control_AWADDR;
	output wire qsort_4_s_axi_control_WREADY;
	input qsort_4_s_axi_control_WVALID;
	input [31:0] qsort_4_s_axi_control_WDATA;
	input [3:0] qsort_4_s_axi_control_WSTRB;
	input qsort_4_s_axi_control_BREADY;
	output wire qsort_4_s_axi_control_BVALID;
	output wire [1:0] qsort_4_s_axi_control_BRESP;
	input qsort_5_m_axi_gmem_ARREADY;
	output wire qsort_5_m_axi_gmem_ARVALID;
	output wire qsort_5_m_axi_gmem_ARID;
	output wire [63:0] qsort_5_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_5_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_5_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_5_m_axi_gmem_ARBURST;
	output wire qsort_5_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_5_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_5_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_5_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_5_m_axi_gmem_ARREGION;
	output wire qsort_5_m_axi_gmem_ARUSER;
	output wire qsort_5_m_axi_gmem_RREADY;
	input qsort_5_m_axi_gmem_RVALID;
	input qsort_5_m_axi_gmem_RID;
	input [63:0] qsort_5_m_axi_gmem_RDATA;
	input [1:0] qsort_5_m_axi_gmem_RRESP;
	input qsort_5_m_axi_gmem_RLAST;
	input qsort_5_m_axi_gmem_RUSER;
	input qsort_5_m_axi_gmem_AWREADY;
	output wire qsort_5_m_axi_gmem_AWVALID;
	output wire qsort_5_m_axi_gmem_AWID;
	output wire [63:0] qsort_5_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_5_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_5_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_5_m_axi_gmem_AWBURST;
	output wire qsort_5_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_5_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_5_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_5_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_5_m_axi_gmem_AWREGION;
	output wire qsort_5_m_axi_gmem_AWUSER;
	input qsort_5_m_axi_gmem_WREADY;
	output wire qsort_5_m_axi_gmem_WVALID;
	output wire [63:0] qsort_5_m_axi_gmem_WDATA;
	output wire [7:0] qsort_5_m_axi_gmem_WSTRB;
	output wire qsort_5_m_axi_gmem_WLAST;
	output wire qsort_5_m_axi_gmem_WUSER;
	output wire qsort_5_m_axi_gmem_BREADY;
	input qsort_5_m_axi_gmem_BVALID;
	input qsort_5_m_axi_gmem_BID;
	input [1:0] qsort_5_m_axi_gmem_BRESP;
	input qsort_5_m_axi_gmem_BUSER;
	output wire qsort_5_s_axi_control_ARREADY;
	input qsort_5_s_axi_control_ARVALID;
	input [5:0] qsort_5_s_axi_control_ARADDR;
	input qsort_5_s_axi_control_RREADY;
	output wire qsort_5_s_axi_control_RVALID;
	output wire [31:0] qsort_5_s_axi_control_RDATA;
	output wire [1:0] qsort_5_s_axi_control_RRESP;
	output wire qsort_5_s_axi_control_AWREADY;
	input qsort_5_s_axi_control_AWVALID;
	input [5:0] qsort_5_s_axi_control_AWADDR;
	output wire qsort_5_s_axi_control_WREADY;
	input qsort_5_s_axi_control_WVALID;
	input [31:0] qsort_5_s_axi_control_WDATA;
	input [3:0] qsort_5_s_axi_control_WSTRB;
	input qsort_5_s_axi_control_BREADY;
	output wire qsort_5_s_axi_control_BVALID;
	output wire [1:0] qsort_5_s_axi_control_BRESP;
	input qsort_6_m_axi_gmem_ARREADY;
	output wire qsort_6_m_axi_gmem_ARVALID;
	output wire qsort_6_m_axi_gmem_ARID;
	output wire [63:0] qsort_6_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_6_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_6_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_6_m_axi_gmem_ARBURST;
	output wire qsort_6_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_6_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_6_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_6_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_6_m_axi_gmem_ARREGION;
	output wire qsort_6_m_axi_gmem_ARUSER;
	output wire qsort_6_m_axi_gmem_RREADY;
	input qsort_6_m_axi_gmem_RVALID;
	input qsort_6_m_axi_gmem_RID;
	input [63:0] qsort_6_m_axi_gmem_RDATA;
	input [1:0] qsort_6_m_axi_gmem_RRESP;
	input qsort_6_m_axi_gmem_RLAST;
	input qsort_6_m_axi_gmem_RUSER;
	input qsort_6_m_axi_gmem_AWREADY;
	output wire qsort_6_m_axi_gmem_AWVALID;
	output wire qsort_6_m_axi_gmem_AWID;
	output wire [63:0] qsort_6_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_6_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_6_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_6_m_axi_gmem_AWBURST;
	output wire qsort_6_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_6_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_6_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_6_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_6_m_axi_gmem_AWREGION;
	output wire qsort_6_m_axi_gmem_AWUSER;
	input qsort_6_m_axi_gmem_WREADY;
	output wire qsort_6_m_axi_gmem_WVALID;
	output wire [63:0] qsort_6_m_axi_gmem_WDATA;
	output wire [7:0] qsort_6_m_axi_gmem_WSTRB;
	output wire qsort_6_m_axi_gmem_WLAST;
	output wire qsort_6_m_axi_gmem_WUSER;
	output wire qsort_6_m_axi_gmem_BREADY;
	input qsort_6_m_axi_gmem_BVALID;
	input qsort_6_m_axi_gmem_BID;
	input [1:0] qsort_6_m_axi_gmem_BRESP;
	input qsort_6_m_axi_gmem_BUSER;
	output wire qsort_6_s_axi_control_ARREADY;
	input qsort_6_s_axi_control_ARVALID;
	input [5:0] qsort_6_s_axi_control_ARADDR;
	input qsort_6_s_axi_control_RREADY;
	output wire qsort_6_s_axi_control_RVALID;
	output wire [31:0] qsort_6_s_axi_control_RDATA;
	output wire [1:0] qsort_6_s_axi_control_RRESP;
	output wire qsort_6_s_axi_control_AWREADY;
	input qsort_6_s_axi_control_AWVALID;
	input [5:0] qsort_6_s_axi_control_AWADDR;
	output wire qsort_6_s_axi_control_WREADY;
	input qsort_6_s_axi_control_WVALID;
	input [31:0] qsort_6_s_axi_control_WDATA;
	input [3:0] qsort_6_s_axi_control_WSTRB;
	input qsort_6_s_axi_control_BREADY;
	output wire qsort_6_s_axi_control_BVALID;
	output wire [1:0] qsort_6_s_axi_control_BRESP;
	input qsort_7_m_axi_gmem_ARREADY;
	output wire qsort_7_m_axi_gmem_ARVALID;
	output wire qsort_7_m_axi_gmem_ARID;
	output wire [63:0] qsort_7_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_7_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_7_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_7_m_axi_gmem_ARBURST;
	output wire qsort_7_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_7_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_7_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_7_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_7_m_axi_gmem_ARREGION;
	output wire qsort_7_m_axi_gmem_ARUSER;
	output wire qsort_7_m_axi_gmem_RREADY;
	input qsort_7_m_axi_gmem_RVALID;
	input qsort_7_m_axi_gmem_RID;
	input [63:0] qsort_7_m_axi_gmem_RDATA;
	input [1:0] qsort_7_m_axi_gmem_RRESP;
	input qsort_7_m_axi_gmem_RLAST;
	input qsort_7_m_axi_gmem_RUSER;
	input qsort_7_m_axi_gmem_AWREADY;
	output wire qsort_7_m_axi_gmem_AWVALID;
	output wire qsort_7_m_axi_gmem_AWID;
	output wire [63:0] qsort_7_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_7_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_7_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_7_m_axi_gmem_AWBURST;
	output wire qsort_7_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_7_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_7_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_7_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_7_m_axi_gmem_AWREGION;
	output wire qsort_7_m_axi_gmem_AWUSER;
	input qsort_7_m_axi_gmem_WREADY;
	output wire qsort_7_m_axi_gmem_WVALID;
	output wire [63:0] qsort_7_m_axi_gmem_WDATA;
	output wire [7:0] qsort_7_m_axi_gmem_WSTRB;
	output wire qsort_7_m_axi_gmem_WLAST;
	output wire qsort_7_m_axi_gmem_WUSER;
	output wire qsort_7_m_axi_gmem_BREADY;
	input qsort_7_m_axi_gmem_BVALID;
	input qsort_7_m_axi_gmem_BID;
	input [1:0] qsort_7_m_axi_gmem_BRESP;
	input qsort_7_m_axi_gmem_BUSER;
	output wire qsort_7_s_axi_control_ARREADY;
	input qsort_7_s_axi_control_ARVALID;
	input [5:0] qsort_7_s_axi_control_ARADDR;
	input qsort_7_s_axi_control_RREADY;
	output wire qsort_7_s_axi_control_RVALID;
	output wire [31:0] qsort_7_s_axi_control_RDATA;
	output wire [1:0] qsort_7_s_axi_control_RRESP;
	output wire qsort_7_s_axi_control_AWREADY;
	input qsort_7_s_axi_control_AWVALID;
	input [5:0] qsort_7_s_axi_control_AWADDR;
	output wire qsort_7_s_axi_control_WREADY;
	input qsort_7_s_axi_control_WVALID;
	input [31:0] qsort_7_s_axi_control_WDATA;
	input [3:0] qsort_7_s_axi_control_WSTRB;
	input qsort_7_s_axi_control_BREADY;
	output wire qsort_7_s_axi_control_BVALID;
	output wire [1:0] qsort_7_s_axi_control_BRESP;
	input qsort_8_m_axi_gmem_ARREADY;
	output wire qsort_8_m_axi_gmem_ARVALID;
	output wire qsort_8_m_axi_gmem_ARID;
	output wire [63:0] qsort_8_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_8_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_8_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_8_m_axi_gmem_ARBURST;
	output wire qsort_8_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_8_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_8_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_8_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_8_m_axi_gmem_ARREGION;
	output wire qsort_8_m_axi_gmem_ARUSER;
	output wire qsort_8_m_axi_gmem_RREADY;
	input qsort_8_m_axi_gmem_RVALID;
	input qsort_8_m_axi_gmem_RID;
	input [63:0] qsort_8_m_axi_gmem_RDATA;
	input [1:0] qsort_8_m_axi_gmem_RRESP;
	input qsort_8_m_axi_gmem_RLAST;
	input qsort_8_m_axi_gmem_RUSER;
	input qsort_8_m_axi_gmem_AWREADY;
	output wire qsort_8_m_axi_gmem_AWVALID;
	output wire qsort_8_m_axi_gmem_AWID;
	output wire [63:0] qsort_8_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_8_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_8_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_8_m_axi_gmem_AWBURST;
	output wire qsort_8_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_8_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_8_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_8_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_8_m_axi_gmem_AWREGION;
	output wire qsort_8_m_axi_gmem_AWUSER;
	input qsort_8_m_axi_gmem_WREADY;
	output wire qsort_8_m_axi_gmem_WVALID;
	output wire [63:0] qsort_8_m_axi_gmem_WDATA;
	output wire [7:0] qsort_8_m_axi_gmem_WSTRB;
	output wire qsort_8_m_axi_gmem_WLAST;
	output wire qsort_8_m_axi_gmem_WUSER;
	output wire qsort_8_m_axi_gmem_BREADY;
	input qsort_8_m_axi_gmem_BVALID;
	input qsort_8_m_axi_gmem_BID;
	input [1:0] qsort_8_m_axi_gmem_BRESP;
	input qsort_8_m_axi_gmem_BUSER;
	output wire qsort_8_s_axi_control_ARREADY;
	input qsort_8_s_axi_control_ARVALID;
	input [5:0] qsort_8_s_axi_control_ARADDR;
	input qsort_8_s_axi_control_RREADY;
	output wire qsort_8_s_axi_control_RVALID;
	output wire [31:0] qsort_8_s_axi_control_RDATA;
	output wire [1:0] qsort_8_s_axi_control_RRESP;
	output wire qsort_8_s_axi_control_AWREADY;
	input qsort_8_s_axi_control_AWVALID;
	input [5:0] qsort_8_s_axi_control_AWADDR;
	output wire qsort_8_s_axi_control_WREADY;
	input qsort_8_s_axi_control_WVALID;
	input [31:0] qsort_8_s_axi_control_WDATA;
	input [3:0] qsort_8_s_axi_control_WSTRB;
	input qsort_8_s_axi_control_BREADY;
	output wire qsort_8_s_axi_control_BVALID;
	output wire [1:0] qsort_8_s_axi_control_BRESP;
	input qsort_9_m_axi_gmem_ARREADY;
	output wire qsort_9_m_axi_gmem_ARVALID;
	output wire qsort_9_m_axi_gmem_ARID;
	output wire [63:0] qsort_9_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_9_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_9_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_9_m_axi_gmem_ARBURST;
	output wire qsort_9_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_9_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_9_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_9_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_9_m_axi_gmem_ARREGION;
	output wire qsort_9_m_axi_gmem_ARUSER;
	output wire qsort_9_m_axi_gmem_RREADY;
	input qsort_9_m_axi_gmem_RVALID;
	input qsort_9_m_axi_gmem_RID;
	input [63:0] qsort_9_m_axi_gmem_RDATA;
	input [1:0] qsort_9_m_axi_gmem_RRESP;
	input qsort_9_m_axi_gmem_RLAST;
	input qsort_9_m_axi_gmem_RUSER;
	input qsort_9_m_axi_gmem_AWREADY;
	output wire qsort_9_m_axi_gmem_AWVALID;
	output wire qsort_9_m_axi_gmem_AWID;
	output wire [63:0] qsort_9_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_9_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_9_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_9_m_axi_gmem_AWBURST;
	output wire qsort_9_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_9_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_9_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_9_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_9_m_axi_gmem_AWREGION;
	output wire qsort_9_m_axi_gmem_AWUSER;
	input qsort_9_m_axi_gmem_WREADY;
	output wire qsort_9_m_axi_gmem_WVALID;
	output wire [63:0] qsort_9_m_axi_gmem_WDATA;
	output wire [7:0] qsort_9_m_axi_gmem_WSTRB;
	output wire qsort_9_m_axi_gmem_WLAST;
	output wire qsort_9_m_axi_gmem_WUSER;
	output wire qsort_9_m_axi_gmem_BREADY;
	input qsort_9_m_axi_gmem_BVALID;
	input qsort_9_m_axi_gmem_BID;
	input [1:0] qsort_9_m_axi_gmem_BRESP;
	input qsort_9_m_axi_gmem_BUSER;
	output wire qsort_9_s_axi_control_ARREADY;
	input qsort_9_s_axi_control_ARVALID;
	input [5:0] qsort_9_s_axi_control_ARADDR;
	input qsort_9_s_axi_control_RREADY;
	output wire qsort_9_s_axi_control_RVALID;
	output wire [31:0] qsort_9_s_axi_control_RDATA;
	output wire [1:0] qsort_9_s_axi_control_RRESP;
	output wire qsort_9_s_axi_control_AWREADY;
	input qsort_9_s_axi_control_AWVALID;
	input [5:0] qsort_9_s_axi_control_AWADDR;
	output wire qsort_9_s_axi_control_WREADY;
	input qsort_9_s_axi_control_WVALID;
	input [31:0] qsort_9_s_axi_control_WDATA;
	input [3:0] qsort_9_s_axi_control_WSTRB;
	input qsort_9_s_axi_control_BREADY;
	output wire qsort_9_s_axi_control_BVALID;
	output wire [1:0] qsort_9_s_axi_control_BRESP;
	input qsort_10_m_axi_gmem_ARREADY;
	output wire qsort_10_m_axi_gmem_ARVALID;
	output wire qsort_10_m_axi_gmem_ARID;
	output wire [63:0] qsort_10_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_10_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_10_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_10_m_axi_gmem_ARBURST;
	output wire qsort_10_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_10_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_10_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_10_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_10_m_axi_gmem_ARREGION;
	output wire qsort_10_m_axi_gmem_ARUSER;
	output wire qsort_10_m_axi_gmem_RREADY;
	input qsort_10_m_axi_gmem_RVALID;
	input qsort_10_m_axi_gmem_RID;
	input [63:0] qsort_10_m_axi_gmem_RDATA;
	input [1:0] qsort_10_m_axi_gmem_RRESP;
	input qsort_10_m_axi_gmem_RLAST;
	input qsort_10_m_axi_gmem_RUSER;
	input qsort_10_m_axi_gmem_AWREADY;
	output wire qsort_10_m_axi_gmem_AWVALID;
	output wire qsort_10_m_axi_gmem_AWID;
	output wire [63:0] qsort_10_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_10_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_10_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_10_m_axi_gmem_AWBURST;
	output wire qsort_10_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_10_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_10_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_10_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_10_m_axi_gmem_AWREGION;
	output wire qsort_10_m_axi_gmem_AWUSER;
	input qsort_10_m_axi_gmem_WREADY;
	output wire qsort_10_m_axi_gmem_WVALID;
	output wire [63:0] qsort_10_m_axi_gmem_WDATA;
	output wire [7:0] qsort_10_m_axi_gmem_WSTRB;
	output wire qsort_10_m_axi_gmem_WLAST;
	output wire qsort_10_m_axi_gmem_WUSER;
	output wire qsort_10_m_axi_gmem_BREADY;
	input qsort_10_m_axi_gmem_BVALID;
	input qsort_10_m_axi_gmem_BID;
	input [1:0] qsort_10_m_axi_gmem_BRESP;
	input qsort_10_m_axi_gmem_BUSER;
	output wire qsort_10_s_axi_control_ARREADY;
	input qsort_10_s_axi_control_ARVALID;
	input [5:0] qsort_10_s_axi_control_ARADDR;
	input qsort_10_s_axi_control_RREADY;
	output wire qsort_10_s_axi_control_RVALID;
	output wire [31:0] qsort_10_s_axi_control_RDATA;
	output wire [1:0] qsort_10_s_axi_control_RRESP;
	output wire qsort_10_s_axi_control_AWREADY;
	input qsort_10_s_axi_control_AWVALID;
	input [5:0] qsort_10_s_axi_control_AWADDR;
	output wire qsort_10_s_axi_control_WREADY;
	input qsort_10_s_axi_control_WVALID;
	input [31:0] qsort_10_s_axi_control_WDATA;
	input [3:0] qsort_10_s_axi_control_WSTRB;
	input qsort_10_s_axi_control_BREADY;
	output wire qsort_10_s_axi_control_BVALID;
	output wire [1:0] qsort_10_s_axi_control_BRESP;
	input qsort_11_m_axi_gmem_ARREADY;
	output wire qsort_11_m_axi_gmem_ARVALID;
	output wire qsort_11_m_axi_gmem_ARID;
	output wire [63:0] qsort_11_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_11_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_11_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_11_m_axi_gmem_ARBURST;
	output wire qsort_11_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_11_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_11_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_11_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_11_m_axi_gmem_ARREGION;
	output wire qsort_11_m_axi_gmem_ARUSER;
	output wire qsort_11_m_axi_gmem_RREADY;
	input qsort_11_m_axi_gmem_RVALID;
	input qsort_11_m_axi_gmem_RID;
	input [63:0] qsort_11_m_axi_gmem_RDATA;
	input [1:0] qsort_11_m_axi_gmem_RRESP;
	input qsort_11_m_axi_gmem_RLAST;
	input qsort_11_m_axi_gmem_RUSER;
	input qsort_11_m_axi_gmem_AWREADY;
	output wire qsort_11_m_axi_gmem_AWVALID;
	output wire qsort_11_m_axi_gmem_AWID;
	output wire [63:0] qsort_11_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_11_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_11_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_11_m_axi_gmem_AWBURST;
	output wire qsort_11_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_11_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_11_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_11_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_11_m_axi_gmem_AWREGION;
	output wire qsort_11_m_axi_gmem_AWUSER;
	input qsort_11_m_axi_gmem_WREADY;
	output wire qsort_11_m_axi_gmem_WVALID;
	output wire [63:0] qsort_11_m_axi_gmem_WDATA;
	output wire [7:0] qsort_11_m_axi_gmem_WSTRB;
	output wire qsort_11_m_axi_gmem_WLAST;
	output wire qsort_11_m_axi_gmem_WUSER;
	output wire qsort_11_m_axi_gmem_BREADY;
	input qsort_11_m_axi_gmem_BVALID;
	input qsort_11_m_axi_gmem_BID;
	input [1:0] qsort_11_m_axi_gmem_BRESP;
	input qsort_11_m_axi_gmem_BUSER;
	output wire qsort_11_s_axi_control_ARREADY;
	input qsort_11_s_axi_control_ARVALID;
	input [5:0] qsort_11_s_axi_control_ARADDR;
	input qsort_11_s_axi_control_RREADY;
	output wire qsort_11_s_axi_control_RVALID;
	output wire [31:0] qsort_11_s_axi_control_RDATA;
	output wire [1:0] qsort_11_s_axi_control_RRESP;
	output wire qsort_11_s_axi_control_AWREADY;
	input qsort_11_s_axi_control_AWVALID;
	input [5:0] qsort_11_s_axi_control_AWADDR;
	output wire qsort_11_s_axi_control_WREADY;
	input qsort_11_s_axi_control_WVALID;
	input [31:0] qsort_11_s_axi_control_WDATA;
	input [3:0] qsort_11_s_axi_control_WSTRB;
	input qsort_11_s_axi_control_BREADY;
	output wire qsort_11_s_axi_control_BVALID;
	output wire [1:0] qsort_11_s_axi_control_BRESP;
	input qsort_12_m_axi_gmem_ARREADY;
	output wire qsort_12_m_axi_gmem_ARVALID;
	output wire qsort_12_m_axi_gmem_ARID;
	output wire [63:0] qsort_12_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_12_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_12_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_12_m_axi_gmem_ARBURST;
	output wire qsort_12_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_12_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_12_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_12_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_12_m_axi_gmem_ARREGION;
	output wire qsort_12_m_axi_gmem_ARUSER;
	output wire qsort_12_m_axi_gmem_RREADY;
	input qsort_12_m_axi_gmem_RVALID;
	input qsort_12_m_axi_gmem_RID;
	input [63:0] qsort_12_m_axi_gmem_RDATA;
	input [1:0] qsort_12_m_axi_gmem_RRESP;
	input qsort_12_m_axi_gmem_RLAST;
	input qsort_12_m_axi_gmem_RUSER;
	input qsort_12_m_axi_gmem_AWREADY;
	output wire qsort_12_m_axi_gmem_AWVALID;
	output wire qsort_12_m_axi_gmem_AWID;
	output wire [63:0] qsort_12_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_12_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_12_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_12_m_axi_gmem_AWBURST;
	output wire qsort_12_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_12_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_12_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_12_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_12_m_axi_gmem_AWREGION;
	output wire qsort_12_m_axi_gmem_AWUSER;
	input qsort_12_m_axi_gmem_WREADY;
	output wire qsort_12_m_axi_gmem_WVALID;
	output wire [63:0] qsort_12_m_axi_gmem_WDATA;
	output wire [7:0] qsort_12_m_axi_gmem_WSTRB;
	output wire qsort_12_m_axi_gmem_WLAST;
	output wire qsort_12_m_axi_gmem_WUSER;
	output wire qsort_12_m_axi_gmem_BREADY;
	input qsort_12_m_axi_gmem_BVALID;
	input qsort_12_m_axi_gmem_BID;
	input [1:0] qsort_12_m_axi_gmem_BRESP;
	input qsort_12_m_axi_gmem_BUSER;
	output wire qsort_12_s_axi_control_ARREADY;
	input qsort_12_s_axi_control_ARVALID;
	input [5:0] qsort_12_s_axi_control_ARADDR;
	input qsort_12_s_axi_control_RREADY;
	output wire qsort_12_s_axi_control_RVALID;
	output wire [31:0] qsort_12_s_axi_control_RDATA;
	output wire [1:0] qsort_12_s_axi_control_RRESP;
	output wire qsort_12_s_axi_control_AWREADY;
	input qsort_12_s_axi_control_AWVALID;
	input [5:0] qsort_12_s_axi_control_AWADDR;
	output wire qsort_12_s_axi_control_WREADY;
	input qsort_12_s_axi_control_WVALID;
	input [31:0] qsort_12_s_axi_control_WDATA;
	input [3:0] qsort_12_s_axi_control_WSTRB;
	input qsort_12_s_axi_control_BREADY;
	output wire qsort_12_s_axi_control_BVALID;
	output wire [1:0] qsort_12_s_axi_control_BRESP;
	input qsort_13_m_axi_gmem_ARREADY;
	output wire qsort_13_m_axi_gmem_ARVALID;
	output wire qsort_13_m_axi_gmem_ARID;
	output wire [63:0] qsort_13_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_13_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_13_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_13_m_axi_gmem_ARBURST;
	output wire qsort_13_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_13_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_13_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_13_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_13_m_axi_gmem_ARREGION;
	output wire qsort_13_m_axi_gmem_ARUSER;
	output wire qsort_13_m_axi_gmem_RREADY;
	input qsort_13_m_axi_gmem_RVALID;
	input qsort_13_m_axi_gmem_RID;
	input [63:0] qsort_13_m_axi_gmem_RDATA;
	input [1:0] qsort_13_m_axi_gmem_RRESP;
	input qsort_13_m_axi_gmem_RLAST;
	input qsort_13_m_axi_gmem_RUSER;
	input qsort_13_m_axi_gmem_AWREADY;
	output wire qsort_13_m_axi_gmem_AWVALID;
	output wire qsort_13_m_axi_gmem_AWID;
	output wire [63:0] qsort_13_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_13_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_13_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_13_m_axi_gmem_AWBURST;
	output wire qsort_13_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_13_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_13_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_13_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_13_m_axi_gmem_AWREGION;
	output wire qsort_13_m_axi_gmem_AWUSER;
	input qsort_13_m_axi_gmem_WREADY;
	output wire qsort_13_m_axi_gmem_WVALID;
	output wire [63:0] qsort_13_m_axi_gmem_WDATA;
	output wire [7:0] qsort_13_m_axi_gmem_WSTRB;
	output wire qsort_13_m_axi_gmem_WLAST;
	output wire qsort_13_m_axi_gmem_WUSER;
	output wire qsort_13_m_axi_gmem_BREADY;
	input qsort_13_m_axi_gmem_BVALID;
	input qsort_13_m_axi_gmem_BID;
	input [1:0] qsort_13_m_axi_gmem_BRESP;
	input qsort_13_m_axi_gmem_BUSER;
	output wire qsort_13_s_axi_control_ARREADY;
	input qsort_13_s_axi_control_ARVALID;
	input [5:0] qsort_13_s_axi_control_ARADDR;
	input qsort_13_s_axi_control_RREADY;
	output wire qsort_13_s_axi_control_RVALID;
	output wire [31:0] qsort_13_s_axi_control_RDATA;
	output wire [1:0] qsort_13_s_axi_control_RRESP;
	output wire qsort_13_s_axi_control_AWREADY;
	input qsort_13_s_axi_control_AWVALID;
	input [5:0] qsort_13_s_axi_control_AWADDR;
	output wire qsort_13_s_axi_control_WREADY;
	input qsort_13_s_axi_control_WVALID;
	input [31:0] qsort_13_s_axi_control_WDATA;
	input [3:0] qsort_13_s_axi_control_WSTRB;
	input qsort_13_s_axi_control_BREADY;
	output wire qsort_13_s_axi_control_BVALID;
	output wire [1:0] qsort_13_s_axi_control_BRESP;
	input qsort_14_m_axi_gmem_ARREADY;
	output wire qsort_14_m_axi_gmem_ARVALID;
	output wire qsort_14_m_axi_gmem_ARID;
	output wire [63:0] qsort_14_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_14_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_14_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_14_m_axi_gmem_ARBURST;
	output wire qsort_14_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_14_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_14_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_14_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_14_m_axi_gmem_ARREGION;
	output wire qsort_14_m_axi_gmem_ARUSER;
	output wire qsort_14_m_axi_gmem_RREADY;
	input qsort_14_m_axi_gmem_RVALID;
	input qsort_14_m_axi_gmem_RID;
	input [63:0] qsort_14_m_axi_gmem_RDATA;
	input [1:0] qsort_14_m_axi_gmem_RRESP;
	input qsort_14_m_axi_gmem_RLAST;
	input qsort_14_m_axi_gmem_RUSER;
	input qsort_14_m_axi_gmem_AWREADY;
	output wire qsort_14_m_axi_gmem_AWVALID;
	output wire qsort_14_m_axi_gmem_AWID;
	output wire [63:0] qsort_14_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_14_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_14_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_14_m_axi_gmem_AWBURST;
	output wire qsort_14_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_14_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_14_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_14_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_14_m_axi_gmem_AWREGION;
	output wire qsort_14_m_axi_gmem_AWUSER;
	input qsort_14_m_axi_gmem_WREADY;
	output wire qsort_14_m_axi_gmem_WVALID;
	output wire [63:0] qsort_14_m_axi_gmem_WDATA;
	output wire [7:0] qsort_14_m_axi_gmem_WSTRB;
	output wire qsort_14_m_axi_gmem_WLAST;
	output wire qsort_14_m_axi_gmem_WUSER;
	output wire qsort_14_m_axi_gmem_BREADY;
	input qsort_14_m_axi_gmem_BVALID;
	input qsort_14_m_axi_gmem_BID;
	input [1:0] qsort_14_m_axi_gmem_BRESP;
	input qsort_14_m_axi_gmem_BUSER;
	output wire qsort_14_s_axi_control_ARREADY;
	input qsort_14_s_axi_control_ARVALID;
	input [5:0] qsort_14_s_axi_control_ARADDR;
	input qsort_14_s_axi_control_RREADY;
	output wire qsort_14_s_axi_control_RVALID;
	output wire [31:0] qsort_14_s_axi_control_RDATA;
	output wire [1:0] qsort_14_s_axi_control_RRESP;
	output wire qsort_14_s_axi_control_AWREADY;
	input qsort_14_s_axi_control_AWVALID;
	input [5:0] qsort_14_s_axi_control_AWADDR;
	output wire qsort_14_s_axi_control_WREADY;
	input qsort_14_s_axi_control_WVALID;
	input [31:0] qsort_14_s_axi_control_WDATA;
	input [3:0] qsort_14_s_axi_control_WSTRB;
	input qsort_14_s_axi_control_BREADY;
	output wire qsort_14_s_axi_control_BVALID;
	output wire [1:0] qsort_14_s_axi_control_BRESP;
	input qsort_15_m_axi_gmem_ARREADY;
	output wire qsort_15_m_axi_gmem_ARVALID;
	output wire qsort_15_m_axi_gmem_ARID;
	output wire [63:0] qsort_15_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_15_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_15_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_15_m_axi_gmem_ARBURST;
	output wire qsort_15_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_15_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_15_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_15_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_15_m_axi_gmem_ARREGION;
	output wire qsort_15_m_axi_gmem_ARUSER;
	output wire qsort_15_m_axi_gmem_RREADY;
	input qsort_15_m_axi_gmem_RVALID;
	input qsort_15_m_axi_gmem_RID;
	input [63:0] qsort_15_m_axi_gmem_RDATA;
	input [1:0] qsort_15_m_axi_gmem_RRESP;
	input qsort_15_m_axi_gmem_RLAST;
	input qsort_15_m_axi_gmem_RUSER;
	input qsort_15_m_axi_gmem_AWREADY;
	output wire qsort_15_m_axi_gmem_AWVALID;
	output wire qsort_15_m_axi_gmem_AWID;
	output wire [63:0] qsort_15_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_15_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_15_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_15_m_axi_gmem_AWBURST;
	output wire qsort_15_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_15_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_15_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_15_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_15_m_axi_gmem_AWREGION;
	output wire qsort_15_m_axi_gmem_AWUSER;
	input qsort_15_m_axi_gmem_WREADY;
	output wire qsort_15_m_axi_gmem_WVALID;
	output wire [63:0] qsort_15_m_axi_gmem_WDATA;
	output wire [7:0] qsort_15_m_axi_gmem_WSTRB;
	output wire qsort_15_m_axi_gmem_WLAST;
	output wire qsort_15_m_axi_gmem_WUSER;
	output wire qsort_15_m_axi_gmem_BREADY;
	input qsort_15_m_axi_gmem_BVALID;
	input qsort_15_m_axi_gmem_BID;
	input [1:0] qsort_15_m_axi_gmem_BRESP;
	input qsort_15_m_axi_gmem_BUSER;
	output wire qsort_15_s_axi_control_ARREADY;
	input qsort_15_s_axi_control_ARVALID;
	input [5:0] qsort_15_s_axi_control_ARADDR;
	input qsort_15_s_axi_control_RREADY;
	output wire qsort_15_s_axi_control_RVALID;
	output wire [31:0] qsort_15_s_axi_control_RDATA;
	output wire [1:0] qsort_15_s_axi_control_RRESP;
	output wire qsort_15_s_axi_control_AWREADY;
	input qsort_15_s_axi_control_AWVALID;
	input [5:0] qsort_15_s_axi_control_AWADDR;
	output wire qsort_15_s_axi_control_WREADY;
	input qsort_15_s_axi_control_WVALID;
	input [31:0] qsort_15_s_axi_control_WDATA;
	input [3:0] qsort_15_s_axi_control_WSTRB;
	input qsort_15_s_axi_control_BREADY;
	output wire qsort_15_s_axi_control_BVALID;
	output wire [1:0] qsort_15_s_axi_control_BRESP;
	input qsort_16_m_axi_gmem_ARREADY;
	output wire qsort_16_m_axi_gmem_ARVALID;
	output wire qsort_16_m_axi_gmem_ARID;
	output wire [63:0] qsort_16_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_16_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_16_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_16_m_axi_gmem_ARBURST;
	output wire qsort_16_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_16_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_16_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_16_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_16_m_axi_gmem_ARREGION;
	output wire qsort_16_m_axi_gmem_ARUSER;
	output wire qsort_16_m_axi_gmem_RREADY;
	input qsort_16_m_axi_gmem_RVALID;
	input qsort_16_m_axi_gmem_RID;
	input [63:0] qsort_16_m_axi_gmem_RDATA;
	input [1:0] qsort_16_m_axi_gmem_RRESP;
	input qsort_16_m_axi_gmem_RLAST;
	input qsort_16_m_axi_gmem_RUSER;
	input qsort_16_m_axi_gmem_AWREADY;
	output wire qsort_16_m_axi_gmem_AWVALID;
	output wire qsort_16_m_axi_gmem_AWID;
	output wire [63:0] qsort_16_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_16_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_16_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_16_m_axi_gmem_AWBURST;
	output wire qsort_16_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_16_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_16_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_16_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_16_m_axi_gmem_AWREGION;
	output wire qsort_16_m_axi_gmem_AWUSER;
	input qsort_16_m_axi_gmem_WREADY;
	output wire qsort_16_m_axi_gmem_WVALID;
	output wire [63:0] qsort_16_m_axi_gmem_WDATA;
	output wire [7:0] qsort_16_m_axi_gmem_WSTRB;
	output wire qsort_16_m_axi_gmem_WLAST;
	output wire qsort_16_m_axi_gmem_WUSER;
	output wire qsort_16_m_axi_gmem_BREADY;
	input qsort_16_m_axi_gmem_BVALID;
	input qsort_16_m_axi_gmem_BID;
	input [1:0] qsort_16_m_axi_gmem_BRESP;
	input qsort_16_m_axi_gmem_BUSER;
	output wire qsort_16_s_axi_control_ARREADY;
	input qsort_16_s_axi_control_ARVALID;
	input [5:0] qsort_16_s_axi_control_ARADDR;
	input qsort_16_s_axi_control_RREADY;
	output wire qsort_16_s_axi_control_RVALID;
	output wire [31:0] qsort_16_s_axi_control_RDATA;
	output wire [1:0] qsort_16_s_axi_control_RRESP;
	output wire qsort_16_s_axi_control_AWREADY;
	input qsort_16_s_axi_control_AWVALID;
	input [5:0] qsort_16_s_axi_control_AWADDR;
	output wire qsort_16_s_axi_control_WREADY;
	input qsort_16_s_axi_control_WVALID;
	input [31:0] qsort_16_s_axi_control_WDATA;
	input [3:0] qsort_16_s_axi_control_WSTRB;
	input qsort_16_s_axi_control_BREADY;
	output wire qsort_16_s_axi_control_BVALID;
	output wire [1:0] qsort_16_s_axi_control_BRESP;
	input qsort_17_m_axi_gmem_ARREADY;
	output wire qsort_17_m_axi_gmem_ARVALID;
	output wire qsort_17_m_axi_gmem_ARID;
	output wire [63:0] qsort_17_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_17_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_17_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_17_m_axi_gmem_ARBURST;
	output wire qsort_17_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_17_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_17_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_17_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_17_m_axi_gmem_ARREGION;
	output wire qsort_17_m_axi_gmem_ARUSER;
	output wire qsort_17_m_axi_gmem_RREADY;
	input qsort_17_m_axi_gmem_RVALID;
	input qsort_17_m_axi_gmem_RID;
	input [63:0] qsort_17_m_axi_gmem_RDATA;
	input [1:0] qsort_17_m_axi_gmem_RRESP;
	input qsort_17_m_axi_gmem_RLAST;
	input qsort_17_m_axi_gmem_RUSER;
	input qsort_17_m_axi_gmem_AWREADY;
	output wire qsort_17_m_axi_gmem_AWVALID;
	output wire qsort_17_m_axi_gmem_AWID;
	output wire [63:0] qsort_17_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_17_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_17_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_17_m_axi_gmem_AWBURST;
	output wire qsort_17_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_17_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_17_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_17_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_17_m_axi_gmem_AWREGION;
	output wire qsort_17_m_axi_gmem_AWUSER;
	input qsort_17_m_axi_gmem_WREADY;
	output wire qsort_17_m_axi_gmem_WVALID;
	output wire [63:0] qsort_17_m_axi_gmem_WDATA;
	output wire [7:0] qsort_17_m_axi_gmem_WSTRB;
	output wire qsort_17_m_axi_gmem_WLAST;
	output wire qsort_17_m_axi_gmem_WUSER;
	output wire qsort_17_m_axi_gmem_BREADY;
	input qsort_17_m_axi_gmem_BVALID;
	input qsort_17_m_axi_gmem_BID;
	input [1:0] qsort_17_m_axi_gmem_BRESP;
	input qsort_17_m_axi_gmem_BUSER;
	output wire qsort_17_s_axi_control_ARREADY;
	input qsort_17_s_axi_control_ARVALID;
	input [5:0] qsort_17_s_axi_control_ARADDR;
	input qsort_17_s_axi_control_RREADY;
	output wire qsort_17_s_axi_control_RVALID;
	output wire [31:0] qsort_17_s_axi_control_RDATA;
	output wire [1:0] qsort_17_s_axi_control_RRESP;
	output wire qsort_17_s_axi_control_AWREADY;
	input qsort_17_s_axi_control_AWVALID;
	input [5:0] qsort_17_s_axi_control_AWADDR;
	output wire qsort_17_s_axi_control_WREADY;
	input qsort_17_s_axi_control_WVALID;
	input [31:0] qsort_17_s_axi_control_WDATA;
	input [3:0] qsort_17_s_axi_control_WSTRB;
	input qsort_17_s_axi_control_BREADY;
	output wire qsort_17_s_axi_control_BVALID;
	output wire [1:0] qsort_17_s_axi_control_BRESP;
	input qsort_18_m_axi_gmem_ARREADY;
	output wire qsort_18_m_axi_gmem_ARVALID;
	output wire qsort_18_m_axi_gmem_ARID;
	output wire [63:0] qsort_18_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_18_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_18_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_18_m_axi_gmem_ARBURST;
	output wire qsort_18_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_18_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_18_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_18_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_18_m_axi_gmem_ARREGION;
	output wire qsort_18_m_axi_gmem_ARUSER;
	output wire qsort_18_m_axi_gmem_RREADY;
	input qsort_18_m_axi_gmem_RVALID;
	input qsort_18_m_axi_gmem_RID;
	input [63:0] qsort_18_m_axi_gmem_RDATA;
	input [1:0] qsort_18_m_axi_gmem_RRESP;
	input qsort_18_m_axi_gmem_RLAST;
	input qsort_18_m_axi_gmem_RUSER;
	input qsort_18_m_axi_gmem_AWREADY;
	output wire qsort_18_m_axi_gmem_AWVALID;
	output wire qsort_18_m_axi_gmem_AWID;
	output wire [63:0] qsort_18_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_18_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_18_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_18_m_axi_gmem_AWBURST;
	output wire qsort_18_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_18_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_18_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_18_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_18_m_axi_gmem_AWREGION;
	output wire qsort_18_m_axi_gmem_AWUSER;
	input qsort_18_m_axi_gmem_WREADY;
	output wire qsort_18_m_axi_gmem_WVALID;
	output wire [63:0] qsort_18_m_axi_gmem_WDATA;
	output wire [7:0] qsort_18_m_axi_gmem_WSTRB;
	output wire qsort_18_m_axi_gmem_WLAST;
	output wire qsort_18_m_axi_gmem_WUSER;
	output wire qsort_18_m_axi_gmem_BREADY;
	input qsort_18_m_axi_gmem_BVALID;
	input qsort_18_m_axi_gmem_BID;
	input [1:0] qsort_18_m_axi_gmem_BRESP;
	input qsort_18_m_axi_gmem_BUSER;
	output wire qsort_18_s_axi_control_ARREADY;
	input qsort_18_s_axi_control_ARVALID;
	input [5:0] qsort_18_s_axi_control_ARADDR;
	input qsort_18_s_axi_control_RREADY;
	output wire qsort_18_s_axi_control_RVALID;
	output wire [31:0] qsort_18_s_axi_control_RDATA;
	output wire [1:0] qsort_18_s_axi_control_RRESP;
	output wire qsort_18_s_axi_control_AWREADY;
	input qsort_18_s_axi_control_AWVALID;
	input [5:0] qsort_18_s_axi_control_AWADDR;
	output wire qsort_18_s_axi_control_WREADY;
	input qsort_18_s_axi_control_WVALID;
	input [31:0] qsort_18_s_axi_control_WDATA;
	input [3:0] qsort_18_s_axi_control_WSTRB;
	input qsort_18_s_axi_control_BREADY;
	output wire qsort_18_s_axi_control_BVALID;
	output wire [1:0] qsort_18_s_axi_control_BRESP;
	input qsort_19_m_axi_gmem_ARREADY;
	output wire qsort_19_m_axi_gmem_ARVALID;
	output wire qsort_19_m_axi_gmem_ARID;
	output wire [63:0] qsort_19_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_19_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_19_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_19_m_axi_gmem_ARBURST;
	output wire qsort_19_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_19_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_19_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_19_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_19_m_axi_gmem_ARREGION;
	output wire qsort_19_m_axi_gmem_ARUSER;
	output wire qsort_19_m_axi_gmem_RREADY;
	input qsort_19_m_axi_gmem_RVALID;
	input qsort_19_m_axi_gmem_RID;
	input [63:0] qsort_19_m_axi_gmem_RDATA;
	input [1:0] qsort_19_m_axi_gmem_RRESP;
	input qsort_19_m_axi_gmem_RLAST;
	input qsort_19_m_axi_gmem_RUSER;
	input qsort_19_m_axi_gmem_AWREADY;
	output wire qsort_19_m_axi_gmem_AWVALID;
	output wire qsort_19_m_axi_gmem_AWID;
	output wire [63:0] qsort_19_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_19_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_19_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_19_m_axi_gmem_AWBURST;
	output wire qsort_19_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_19_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_19_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_19_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_19_m_axi_gmem_AWREGION;
	output wire qsort_19_m_axi_gmem_AWUSER;
	input qsort_19_m_axi_gmem_WREADY;
	output wire qsort_19_m_axi_gmem_WVALID;
	output wire [63:0] qsort_19_m_axi_gmem_WDATA;
	output wire [7:0] qsort_19_m_axi_gmem_WSTRB;
	output wire qsort_19_m_axi_gmem_WLAST;
	output wire qsort_19_m_axi_gmem_WUSER;
	output wire qsort_19_m_axi_gmem_BREADY;
	input qsort_19_m_axi_gmem_BVALID;
	input qsort_19_m_axi_gmem_BID;
	input [1:0] qsort_19_m_axi_gmem_BRESP;
	input qsort_19_m_axi_gmem_BUSER;
	output wire qsort_19_s_axi_control_ARREADY;
	input qsort_19_s_axi_control_ARVALID;
	input [5:0] qsort_19_s_axi_control_ARADDR;
	input qsort_19_s_axi_control_RREADY;
	output wire qsort_19_s_axi_control_RVALID;
	output wire [31:0] qsort_19_s_axi_control_RDATA;
	output wire [1:0] qsort_19_s_axi_control_RRESP;
	output wire qsort_19_s_axi_control_AWREADY;
	input qsort_19_s_axi_control_AWVALID;
	input [5:0] qsort_19_s_axi_control_AWADDR;
	output wire qsort_19_s_axi_control_WREADY;
	input qsort_19_s_axi_control_WVALID;
	input [31:0] qsort_19_s_axi_control_WDATA;
	input [3:0] qsort_19_s_axi_control_WSTRB;
	input qsort_19_s_axi_control_BREADY;
	output wire qsort_19_s_axi_control_BVALID;
	output wire [1:0] qsort_19_s_axi_control_BRESP;
	input qsort_20_m_axi_gmem_ARREADY;
	output wire qsort_20_m_axi_gmem_ARVALID;
	output wire qsort_20_m_axi_gmem_ARID;
	output wire [63:0] qsort_20_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_20_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_20_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_20_m_axi_gmem_ARBURST;
	output wire qsort_20_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_20_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_20_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_20_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_20_m_axi_gmem_ARREGION;
	output wire qsort_20_m_axi_gmem_ARUSER;
	output wire qsort_20_m_axi_gmem_RREADY;
	input qsort_20_m_axi_gmem_RVALID;
	input qsort_20_m_axi_gmem_RID;
	input [63:0] qsort_20_m_axi_gmem_RDATA;
	input [1:0] qsort_20_m_axi_gmem_RRESP;
	input qsort_20_m_axi_gmem_RLAST;
	input qsort_20_m_axi_gmem_RUSER;
	input qsort_20_m_axi_gmem_AWREADY;
	output wire qsort_20_m_axi_gmem_AWVALID;
	output wire qsort_20_m_axi_gmem_AWID;
	output wire [63:0] qsort_20_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_20_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_20_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_20_m_axi_gmem_AWBURST;
	output wire qsort_20_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_20_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_20_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_20_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_20_m_axi_gmem_AWREGION;
	output wire qsort_20_m_axi_gmem_AWUSER;
	input qsort_20_m_axi_gmem_WREADY;
	output wire qsort_20_m_axi_gmem_WVALID;
	output wire [63:0] qsort_20_m_axi_gmem_WDATA;
	output wire [7:0] qsort_20_m_axi_gmem_WSTRB;
	output wire qsort_20_m_axi_gmem_WLAST;
	output wire qsort_20_m_axi_gmem_WUSER;
	output wire qsort_20_m_axi_gmem_BREADY;
	input qsort_20_m_axi_gmem_BVALID;
	input qsort_20_m_axi_gmem_BID;
	input [1:0] qsort_20_m_axi_gmem_BRESP;
	input qsort_20_m_axi_gmem_BUSER;
	output wire qsort_20_s_axi_control_ARREADY;
	input qsort_20_s_axi_control_ARVALID;
	input [5:0] qsort_20_s_axi_control_ARADDR;
	input qsort_20_s_axi_control_RREADY;
	output wire qsort_20_s_axi_control_RVALID;
	output wire [31:0] qsort_20_s_axi_control_RDATA;
	output wire [1:0] qsort_20_s_axi_control_RRESP;
	output wire qsort_20_s_axi_control_AWREADY;
	input qsort_20_s_axi_control_AWVALID;
	input [5:0] qsort_20_s_axi_control_AWADDR;
	output wire qsort_20_s_axi_control_WREADY;
	input qsort_20_s_axi_control_WVALID;
	input [31:0] qsort_20_s_axi_control_WDATA;
	input [3:0] qsort_20_s_axi_control_WSTRB;
	input qsort_20_s_axi_control_BREADY;
	output wire qsort_20_s_axi_control_BVALID;
	output wire [1:0] qsort_20_s_axi_control_BRESP;
	input qsort_21_m_axi_gmem_ARREADY;
	output wire qsort_21_m_axi_gmem_ARVALID;
	output wire qsort_21_m_axi_gmem_ARID;
	output wire [63:0] qsort_21_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_21_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_21_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_21_m_axi_gmem_ARBURST;
	output wire qsort_21_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_21_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_21_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_21_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_21_m_axi_gmem_ARREGION;
	output wire qsort_21_m_axi_gmem_ARUSER;
	output wire qsort_21_m_axi_gmem_RREADY;
	input qsort_21_m_axi_gmem_RVALID;
	input qsort_21_m_axi_gmem_RID;
	input [63:0] qsort_21_m_axi_gmem_RDATA;
	input [1:0] qsort_21_m_axi_gmem_RRESP;
	input qsort_21_m_axi_gmem_RLAST;
	input qsort_21_m_axi_gmem_RUSER;
	input qsort_21_m_axi_gmem_AWREADY;
	output wire qsort_21_m_axi_gmem_AWVALID;
	output wire qsort_21_m_axi_gmem_AWID;
	output wire [63:0] qsort_21_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_21_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_21_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_21_m_axi_gmem_AWBURST;
	output wire qsort_21_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_21_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_21_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_21_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_21_m_axi_gmem_AWREGION;
	output wire qsort_21_m_axi_gmem_AWUSER;
	input qsort_21_m_axi_gmem_WREADY;
	output wire qsort_21_m_axi_gmem_WVALID;
	output wire [63:0] qsort_21_m_axi_gmem_WDATA;
	output wire [7:0] qsort_21_m_axi_gmem_WSTRB;
	output wire qsort_21_m_axi_gmem_WLAST;
	output wire qsort_21_m_axi_gmem_WUSER;
	output wire qsort_21_m_axi_gmem_BREADY;
	input qsort_21_m_axi_gmem_BVALID;
	input qsort_21_m_axi_gmem_BID;
	input [1:0] qsort_21_m_axi_gmem_BRESP;
	input qsort_21_m_axi_gmem_BUSER;
	output wire qsort_21_s_axi_control_ARREADY;
	input qsort_21_s_axi_control_ARVALID;
	input [5:0] qsort_21_s_axi_control_ARADDR;
	input qsort_21_s_axi_control_RREADY;
	output wire qsort_21_s_axi_control_RVALID;
	output wire [31:0] qsort_21_s_axi_control_RDATA;
	output wire [1:0] qsort_21_s_axi_control_RRESP;
	output wire qsort_21_s_axi_control_AWREADY;
	input qsort_21_s_axi_control_AWVALID;
	input [5:0] qsort_21_s_axi_control_AWADDR;
	output wire qsort_21_s_axi_control_WREADY;
	input qsort_21_s_axi_control_WVALID;
	input [31:0] qsort_21_s_axi_control_WDATA;
	input [3:0] qsort_21_s_axi_control_WSTRB;
	input qsort_21_s_axi_control_BREADY;
	output wire qsort_21_s_axi_control_BVALID;
	output wire [1:0] qsort_21_s_axi_control_BRESP;
	input qsort_22_m_axi_gmem_ARREADY;
	output wire qsort_22_m_axi_gmem_ARVALID;
	output wire qsort_22_m_axi_gmem_ARID;
	output wire [63:0] qsort_22_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_22_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_22_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_22_m_axi_gmem_ARBURST;
	output wire qsort_22_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_22_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_22_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_22_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_22_m_axi_gmem_ARREGION;
	output wire qsort_22_m_axi_gmem_ARUSER;
	output wire qsort_22_m_axi_gmem_RREADY;
	input qsort_22_m_axi_gmem_RVALID;
	input qsort_22_m_axi_gmem_RID;
	input [63:0] qsort_22_m_axi_gmem_RDATA;
	input [1:0] qsort_22_m_axi_gmem_RRESP;
	input qsort_22_m_axi_gmem_RLAST;
	input qsort_22_m_axi_gmem_RUSER;
	input qsort_22_m_axi_gmem_AWREADY;
	output wire qsort_22_m_axi_gmem_AWVALID;
	output wire qsort_22_m_axi_gmem_AWID;
	output wire [63:0] qsort_22_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_22_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_22_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_22_m_axi_gmem_AWBURST;
	output wire qsort_22_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_22_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_22_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_22_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_22_m_axi_gmem_AWREGION;
	output wire qsort_22_m_axi_gmem_AWUSER;
	input qsort_22_m_axi_gmem_WREADY;
	output wire qsort_22_m_axi_gmem_WVALID;
	output wire [63:0] qsort_22_m_axi_gmem_WDATA;
	output wire [7:0] qsort_22_m_axi_gmem_WSTRB;
	output wire qsort_22_m_axi_gmem_WLAST;
	output wire qsort_22_m_axi_gmem_WUSER;
	output wire qsort_22_m_axi_gmem_BREADY;
	input qsort_22_m_axi_gmem_BVALID;
	input qsort_22_m_axi_gmem_BID;
	input [1:0] qsort_22_m_axi_gmem_BRESP;
	input qsort_22_m_axi_gmem_BUSER;
	output wire qsort_22_s_axi_control_ARREADY;
	input qsort_22_s_axi_control_ARVALID;
	input [5:0] qsort_22_s_axi_control_ARADDR;
	input qsort_22_s_axi_control_RREADY;
	output wire qsort_22_s_axi_control_RVALID;
	output wire [31:0] qsort_22_s_axi_control_RDATA;
	output wire [1:0] qsort_22_s_axi_control_RRESP;
	output wire qsort_22_s_axi_control_AWREADY;
	input qsort_22_s_axi_control_AWVALID;
	input [5:0] qsort_22_s_axi_control_AWADDR;
	output wire qsort_22_s_axi_control_WREADY;
	input qsort_22_s_axi_control_WVALID;
	input [31:0] qsort_22_s_axi_control_WDATA;
	input [3:0] qsort_22_s_axi_control_WSTRB;
	input qsort_22_s_axi_control_BREADY;
	output wire qsort_22_s_axi_control_BVALID;
	output wire [1:0] qsort_22_s_axi_control_BRESP;
	input qsort_23_m_axi_gmem_ARREADY;
	output wire qsort_23_m_axi_gmem_ARVALID;
	output wire qsort_23_m_axi_gmem_ARID;
	output wire [63:0] qsort_23_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_23_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_23_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_23_m_axi_gmem_ARBURST;
	output wire qsort_23_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_23_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_23_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_23_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_23_m_axi_gmem_ARREGION;
	output wire qsort_23_m_axi_gmem_ARUSER;
	output wire qsort_23_m_axi_gmem_RREADY;
	input qsort_23_m_axi_gmem_RVALID;
	input qsort_23_m_axi_gmem_RID;
	input [63:0] qsort_23_m_axi_gmem_RDATA;
	input [1:0] qsort_23_m_axi_gmem_RRESP;
	input qsort_23_m_axi_gmem_RLAST;
	input qsort_23_m_axi_gmem_RUSER;
	input qsort_23_m_axi_gmem_AWREADY;
	output wire qsort_23_m_axi_gmem_AWVALID;
	output wire qsort_23_m_axi_gmem_AWID;
	output wire [63:0] qsort_23_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_23_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_23_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_23_m_axi_gmem_AWBURST;
	output wire qsort_23_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_23_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_23_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_23_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_23_m_axi_gmem_AWREGION;
	output wire qsort_23_m_axi_gmem_AWUSER;
	input qsort_23_m_axi_gmem_WREADY;
	output wire qsort_23_m_axi_gmem_WVALID;
	output wire [63:0] qsort_23_m_axi_gmem_WDATA;
	output wire [7:0] qsort_23_m_axi_gmem_WSTRB;
	output wire qsort_23_m_axi_gmem_WLAST;
	output wire qsort_23_m_axi_gmem_WUSER;
	output wire qsort_23_m_axi_gmem_BREADY;
	input qsort_23_m_axi_gmem_BVALID;
	input qsort_23_m_axi_gmem_BID;
	input [1:0] qsort_23_m_axi_gmem_BRESP;
	input qsort_23_m_axi_gmem_BUSER;
	output wire qsort_23_s_axi_control_ARREADY;
	input qsort_23_s_axi_control_ARVALID;
	input [5:0] qsort_23_s_axi_control_ARADDR;
	input qsort_23_s_axi_control_RREADY;
	output wire qsort_23_s_axi_control_RVALID;
	output wire [31:0] qsort_23_s_axi_control_RDATA;
	output wire [1:0] qsort_23_s_axi_control_RRESP;
	output wire qsort_23_s_axi_control_AWREADY;
	input qsort_23_s_axi_control_AWVALID;
	input [5:0] qsort_23_s_axi_control_AWADDR;
	output wire qsort_23_s_axi_control_WREADY;
	input qsort_23_s_axi_control_WVALID;
	input [31:0] qsort_23_s_axi_control_WDATA;
	input [3:0] qsort_23_s_axi_control_WSTRB;
	input qsort_23_s_axi_control_BREADY;
	output wire qsort_23_s_axi_control_BVALID;
	output wire [1:0] qsort_23_s_axi_control_BRESP;
	input qsort_24_m_axi_gmem_ARREADY;
	output wire qsort_24_m_axi_gmem_ARVALID;
	output wire qsort_24_m_axi_gmem_ARID;
	output wire [63:0] qsort_24_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_24_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_24_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_24_m_axi_gmem_ARBURST;
	output wire qsort_24_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_24_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_24_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_24_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_24_m_axi_gmem_ARREGION;
	output wire qsort_24_m_axi_gmem_ARUSER;
	output wire qsort_24_m_axi_gmem_RREADY;
	input qsort_24_m_axi_gmem_RVALID;
	input qsort_24_m_axi_gmem_RID;
	input [63:0] qsort_24_m_axi_gmem_RDATA;
	input [1:0] qsort_24_m_axi_gmem_RRESP;
	input qsort_24_m_axi_gmem_RLAST;
	input qsort_24_m_axi_gmem_RUSER;
	input qsort_24_m_axi_gmem_AWREADY;
	output wire qsort_24_m_axi_gmem_AWVALID;
	output wire qsort_24_m_axi_gmem_AWID;
	output wire [63:0] qsort_24_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_24_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_24_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_24_m_axi_gmem_AWBURST;
	output wire qsort_24_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_24_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_24_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_24_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_24_m_axi_gmem_AWREGION;
	output wire qsort_24_m_axi_gmem_AWUSER;
	input qsort_24_m_axi_gmem_WREADY;
	output wire qsort_24_m_axi_gmem_WVALID;
	output wire [63:0] qsort_24_m_axi_gmem_WDATA;
	output wire [7:0] qsort_24_m_axi_gmem_WSTRB;
	output wire qsort_24_m_axi_gmem_WLAST;
	output wire qsort_24_m_axi_gmem_WUSER;
	output wire qsort_24_m_axi_gmem_BREADY;
	input qsort_24_m_axi_gmem_BVALID;
	input qsort_24_m_axi_gmem_BID;
	input [1:0] qsort_24_m_axi_gmem_BRESP;
	input qsort_24_m_axi_gmem_BUSER;
	output wire qsort_24_s_axi_control_ARREADY;
	input qsort_24_s_axi_control_ARVALID;
	input [5:0] qsort_24_s_axi_control_ARADDR;
	input qsort_24_s_axi_control_RREADY;
	output wire qsort_24_s_axi_control_RVALID;
	output wire [31:0] qsort_24_s_axi_control_RDATA;
	output wire [1:0] qsort_24_s_axi_control_RRESP;
	output wire qsort_24_s_axi_control_AWREADY;
	input qsort_24_s_axi_control_AWVALID;
	input [5:0] qsort_24_s_axi_control_AWADDR;
	output wire qsort_24_s_axi_control_WREADY;
	input qsort_24_s_axi_control_WVALID;
	input [31:0] qsort_24_s_axi_control_WDATA;
	input [3:0] qsort_24_s_axi_control_WSTRB;
	input qsort_24_s_axi_control_BREADY;
	output wire qsort_24_s_axi_control_BVALID;
	output wire [1:0] qsort_24_s_axi_control_BRESP;
	input qsort_25_m_axi_gmem_ARREADY;
	output wire qsort_25_m_axi_gmem_ARVALID;
	output wire qsort_25_m_axi_gmem_ARID;
	output wire [63:0] qsort_25_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_25_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_25_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_25_m_axi_gmem_ARBURST;
	output wire qsort_25_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_25_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_25_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_25_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_25_m_axi_gmem_ARREGION;
	output wire qsort_25_m_axi_gmem_ARUSER;
	output wire qsort_25_m_axi_gmem_RREADY;
	input qsort_25_m_axi_gmem_RVALID;
	input qsort_25_m_axi_gmem_RID;
	input [63:0] qsort_25_m_axi_gmem_RDATA;
	input [1:0] qsort_25_m_axi_gmem_RRESP;
	input qsort_25_m_axi_gmem_RLAST;
	input qsort_25_m_axi_gmem_RUSER;
	input qsort_25_m_axi_gmem_AWREADY;
	output wire qsort_25_m_axi_gmem_AWVALID;
	output wire qsort_25_m_axi_gmem_AWID;
	output wire [63:0] qsort_25_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_25_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_25_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_25_m_axi_gmem_AWBURST;
	output wire qsort_25_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_25_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_25_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_25_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_25_m_axi_gmem_AWREGION;
	output wire qsort_25_m_axi_gmem_AWUSER;
	input qsort_25_m_axi_gmem_WREADY;
	output wire qsort_25_m_axi_gmem_WVALID;
	output wire [63:0] qsort_25_m_axi_gmem_WDATA;
	output wire [7:0] qsort_25_m_axi_gmem_WSTRB;
	output wire qsort_25_m_axi_gmem_WLAST;
	output wire qsort_25_m_axi_gmem_WUSER;
	output wire qsort_25_m_axi_gmem_BREADY;
	input qsort_25_m_axi_gmem_BVALID;
	input qsort_25_m_axi_gmem_BID;
	input [1:0] qsort_25_m_axi_gmem_BRESP;
	input qsort_25_m_axi_gmem_BUSER;
	output wire qsort_25_s_axi_control_ARREADY;
	input qsort_25_s_axi_control_ARVALID;
	input [5:0] qsort_25_s_axi_control_ARADDR;
	input qsort_25_s_axi_control_RREADY;
	output wire qsort_25_s_axi_control_RVALID;
	output wire [31:0] qsort_25_s_axi_control_RDATA;
	output wire [1:0] qsort_25_s_axi_control_RRESP;
	output wire qsort_25_s_axi_control_AWREADY;
	input qsort_25_s_axi_control_AWVALID;
	input [5:0] qsort_25_s_axi_control_AWADDR;
	output wire qsort_25_s_axi_control_WREADY;
	input qsort_25_s_axi_control_WVALID;
	input [31:0] qsort_25_s_axi_control_WDATA;
	input [3:0] qsort_25_s_axi_control_WSTRB;
	input qsort_25_s_axi_control_BREADY;
	output wire qsort_25_s_axi_control_BVALID;
	output wire [1:0] qsort_25_s_axi_control_BRESP;
	input qsort_26_m_axi_gmem_ARREADY;
	output wire qsort_26_m_axi_gmem_ARVALID;
	output wire qsort_26_m_axi_gmem_ARID;
	output wire [63:0] qsort_26_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_26_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_26_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_26_m_axi_gmem_ARBURST;
	output wire qsort_26_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_26_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_26_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_26_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_26_m_axi_gmem_ARREGION;
	output wire qsort_26_m_axi_gmem_ARUSER;
	output wire qsort_26_m_axi_gmem_RREADY;
	input qsort_26_m_axi_gmem_RVALID;
	input qsort_26_m_axi_gmem_RID;
	input [63:0] qsort_26_m_axi_gmem_RDATA;
	input [1:0] qsort_26_m_axi_gmem_RRESP;
	input qsort_26_m_axi_gmem_RLAST;
	input qsort_26_m_axi_gmem_RUSER;
	input qsort_26_m_axi_gmem_AWREADY;
	output wire qsort_26_m_axi_gmem_AWVALID;
	output wire qsort_26_m_axi_gmem_AWID;
	output wire [63:0] qsort_26_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_26_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_26_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_26_m_axi_gmem_AWBURST;
	output wire qsort_26_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_26_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_26_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_26_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_26_m_axi_gmem_AWREGION;
	output wire qsort_26_m_axi_gmem_AWUSER;
	input qsort_26_m_axi_gmem_WREADY;
	output wire qsort_26_m_axi_gmem_WVALID;
	output wire [63:0] qsort_26_m_axi_gmem_WDATA;
	output wire [7:0] qsort_26_m_axi_gmem_WSTRB;
	output wire qsort_26_m_axi_gmem_WLAST;
	output wire qsort_26_m_axi_gmem_WUSER;
	output wire qsort_26_m_axi_gmem_BREADY;
	input qsort_26_m_axi_gmem_BVALID;
	input qsort_26_m_axi_gmem_BID;
	input [1:0] qsort_26_m_axi_gmem_BRESP;
	input qsort_26_m_axi_gmem_BUSER;
	output wire qsort_26_s_axi_control_ARREADY;
	input qsort_26_s_axi_control_ARVALID;
	input [5:0] qsort_26_s_axi_control_ARADDR;
	input qsort_26_s_axi_control_RREADY;
	output wire qsort_26_s_axi_control_RVALID;
	output wire [31:0] qsort_26_s_axi_control_RDATA;
	output wire [1:0] qsort_26_s_axi_control_RRESP;
	output wire qsort_26_s_axi_control_AWREADY;
	input qsort_26_s_axi_control_AWVALID;
	input [5:0] qsort_26_s_axi_control_AWADDR;
	output wire qsort_26_s_axi_control_WREADY;
	input qsort_26_s_axi_control_WVALID;
	input [31:0] qsort_26_s_axi_control_WDATA;
	input [3:0] qsort_26_s_axi_control_WSTRB;
	input qsort_26_s_axi_control_BREADY;
	output wire qsort_26_s_axi_control_BVALID;
	output wire [1:0] qsort_26_s_axi_control_BRESP;
	input qsort_27_m_axi_gmem_ARREADY;
	output wire qsort_27_m_axi_gmem_ARVALID;
	output wire qsort_27_m_axi_gmem_ARID;
	output wire [63:0] qsort_27_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_27_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_27_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_27_m_axi_gmem_ARBURST;
	output wire qsort_27_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_27_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_27_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_27_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_27_m_axi_gmem_ARREGION;
	output wire qsort_27_m_axi_gmem_ARUSER;
	output wire qsort_27_m_axi_gmem_RREADY;
	input qsort_27_m_axi_gmem_RVALID;
	input qsort_27_m_axi_gmem_RID;
	input [63:0] qsort_27_m_axi_gmem_RDATA;
	input [1:0] qsort_27_m_axi_gmem_RRESP;
	input qsort_27_m_axi_gmem_RLAST;
	input qsort_27_m_axi_gmem_RUSER;
	input qsort_27_m_axi_gmem_AWREADY;
	output wire qsort_27_m_axi_gmem_AWVALID;
	output wire qsort_27_m_axi_gmem_AWID;
	output wire [63:0] qsort_27_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_27_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_27_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_27_m_axi_gmem_AWBURST;
	output wire qsort_27_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_27_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_27_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_27_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_27_m_axi_gmem_AWREGION;
	output wire qsort_27_m_axi_gmem_AWUSER;
	input qsort_27_m_axi_gmem_WREADY;
	output wire qsort_27_m_axi_gmem_WVALID;
	output wire [63:0] qsort_27_m_axi_gmem_WDATA;
	output wire [7:0] qsort_27_m_axi_gmem_WSTRB;
	output wire qsort_27_m_axi_gmem_WLAST;
	output wire qsort_27_m_axi_gmem_WUSER;
	output wire qsort_27_m_axi_gmem_BREADY;
	input qsort_27_m_axi_gmem_BVALID;
	input qsort_27_m_axi_gmem_BID;
	input [1:0] qsort_27_m_axi_gmem_BRESP;
	input qsort_27_m_axi_gmem_BUSER;
	output wire qsort_27_s_axi_control_ARREADY;
	input qsort_27_s_axi_control_ARVALID;
	input [5:0] qsort_27_s_axi_control_ARADDR;
	input qsort_27_s_axi_control_RREADY;
	output wire qsort_27_s_axi_control_RVALID;
	output wire [31:0] qsort_27_s_axi_control_RDATA;
	output wire [1:0] qsort_27_s_axi_control_RRESP;
	output wire qsort_27_s_axi_control_AWREADY;
	input qsort_27_s_axi_control_AWVALID;
	input [5:0] qsort_27_s_axi_control_AWADDR;
	output wire qsort_27_s_axi_control_WREADY;
	input qsort_27_s_axi_control_WVALID;
	input [31:0] qsort_27_s_axi_control_WDATA;
	input [3:0] qsort_27_s_axi_control_WSTRB;
	input qsort_27_s_axi_control_BREADY;
	output wire qsort_27_s_axi_control_BVALID;
	output wire [1:0] qsort_27_s_axi_control_BRESP;
	input qsort_28_m_axi_gmem_ARREADY;
	output wire qsort_28_m_axi_gmem_ARVALID;
	output wire qsort_28_m_axi_gmem_ARID;
	output wire [63:0] qsort_28_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_28_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_28_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_28_m_axi_gmem_ARBURST;
	output wire qsort_28_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_28_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_28_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_28_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_28_m_axi_gmem_ARREGION;
	output wire qsort_28_m_axi_gmem_ARUSER;
	output wire qsort_28_m_axi_gmem_RREADY;
	input qsort_28_m_axi_gmem_RVALID;
	input qsort_28_m_axi_gmem_RID;
	input [63:0] qsort_28_m_axi_gmem_RDATA;
	input [1:0] qsort_28_m_axi_gmem_RRESP;
	input qsort_28_m_axi_gmem_RLAST;
	input qsort_28_m_axi_gmem_RUSER;
	input qsort_28_m_axi_gmem_AWREADY;
	output wire qsort_28_m_axi_gmem_AWVALID;
	output wire qsort_28_m_axi_gmem_AWID;
	output wire [63:0] qsort_28_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_28_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_28_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_28_m_axi_gmem_AWBURST;
	output wire qsort_28_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_28_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_28_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_28_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_28_m_axi_gmem_AWREGION;
	output wire qsort_28_m_axi_gmem_AWUSER;
	input qsort_28_m_axi_gmem_WREADY;
	output wire qsort_28_m_axi_gmem_WVALID;
	output wire [63:0] qsort_28_m_axi_gmem_WDATA;
	output wire [7:0] qsort_28_m_axi_gmem_WSTRB;
	output wire qsort_28_m_axi_gmem_WLAST;
	output wire qsort_28_m_axi_gmem_WUSER;
	output wire qsort_28_m_axi_gmem_BREADY;
	input qsort_28_m_axi_gmem_BVALID;
	input qsort_28_m_axi_gmem_BID;
	input [1:0] qsort_28_m_axi_gmem_BRESP;
	input qsort_28_m_axi_gmem_BUSER;
	output wire qsort_28_s_axi_control_ARREADY;
	input qsort_28_s_axi_control_ARVALID;
	input [5:0] qsort_28_s_axi_control_ARADDR;
	input qsort_28_s_axi_control_RREADY;
	output wire qsort_28_s_axi_control_RVALID;
	output wire [31:0] qsort_28_s_axi_control_RDATA;
	output wire [1:0] qsort_28_s_axi_control_RRESP;
	output wire qsort_28_s_axi_control_AWREADY;
	input qsort_28_s_axi_control_AWVALID;
	input [5:0] qsort_28_s_axi_control_AWADDR;
	output wire qsort_28_s_axi_control_WREADY;
	input qsort_28_s_axi_control_WVALID;
	input [31:0] qsort_28_s_axi_control_WDATA;
	input [3:0] qsort_28_s_axi_control_WSTRB;
	input qsort_28_s_axi_control_BREADY;
	output wire qsort_28_s_axi_control_BVALID;
	output wire [1:0] qsort_28_s_axi_control_BRESP;
	input qsort_29_m_axi_gmem_ARREADY;
	output wire qsort_29_m_axi_gmem_ARVALID;
	output wire qsort_29_m_axi_gmem_ARID;
	output wire [63:0] qsort_29_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_29_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_29_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_29_m_axi_gmem_ARBURST;
	output wire qsort_29_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_29_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_29_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_29_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_29_m_axi_gmem_ARREGION;
	output wire qsort_29_m_axi_gmem_ARUSER;
	output wire qsort_29_m_axi_gmem_RREADY;
	input qsort_29_m_axi_gmem_RVALID;
	input qsort_29_m_axi_gmem_RID;
	input [63:0] qsort_29_m_axi_gmem_RDATA;
	input [1:0] qsort_29_m_axi_gmem_RRESP;
	input qsort_29_m_axi_gmem_RLAST;
	input qsort_29_m_axi_gmem_RUSER;
	input qsort_29_m_axi_gmem_AWREADY;
	output wire qsort_29_m_axi_gmem_AWVALID;
	output wire qsort_29_m_axi_gmem_AWID;
	output wire [63:0] qsort_29_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_29_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_29_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_29_m_axi_gmem_AWBURST;
	output wire qsort_29_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_29_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_29_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_29_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_29_m_axi_gmem_AWREGION;
	output wire qsort_29_m_axi_gmem_AWUSER;
	input qsort_29_m_axi_gmem_WREADY;
	output wire qsort_29_m_axi_gmem_WVALID;
	output wire [63:0] qsort_29_m_axi_gmem_WDATA;
	output wire [7:0] qsort_29_m_axi_gmem_WSTRB;
	output wire qsort_29_m_axi_gmem_WLAST;
	output wire qsort_29_m_axi_gmem_WUSER;
	output wire qsort_29_m_axi_gmem_BREADY;
	input qsort_29_m_axi_gmem_BVALID;
	input qsort_29_m_axi_gmem_BID;
	input [1:0] qsort_29_m_axi_gmem_BRESP;
	input qsort_29_m_axi_gmem_BUSER;
	output wire qsort_29_s_axi_control_ARREADY;
	input qsort_29_s_axi_control_ARVALID;
	input [5:0] qsort_29_s_axi_control_ARADDR;
	input qsort_29_s_axi_control_RREADY;
	output wire qsort_29_s_axi_control_RVALID;
	output wire [31:0] qsort_29_s_axi_control_RDATA;
	output wire [1:0] qsort_29_s_axi_control_RRESP;
	output wire qsort_29_s_axi_control_AWREADY;
	input qsort_29_s_axi_control_AWVALID;
	input [5:0] qsort_29_s_axi_control_AWADDR;
	output wire qsort_29_s_axi_control_WREADY;
	input qsort_29_s_axi_control_WVALID;
	input [31:0] qsort_29_s_axi_control_WDATA;
	input [3:0] qsort_29_s_axi_control_WSTRB;
	input qsort_29_s_axi_control_BREADY;
	output wire qsort_29_s_axi_control_BVALID;
	output wire [1:0] qsort_29_s_axi_control_BRESP;
	input qsort_30_m_axi_gmem_ARREADY;
	output wire qsort_30_m_axi_gmem_ARVALID;
	output wire qsort_30_m_axi_gmem_ARID;
	output wire [63:0] qsort_30_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_30_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_30_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_30_m_axi_gmem_ARBURST;
	output wire qsort_30_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_30_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_30_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_30_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_30_m_axi_gmem_ARREGION;
	output wire qsort_30_m_axi_gmem_ARUSER;
	output wire qsort_30_m_axi_gmem_RREADY;
	input qsort_30_m_axi_gmem_RVALID;
	input qsort_30_m_axi_gmem_RID;
	input [63:0] qsort_30_m_axi_gmem_RDATA;
	input [1:0] qsort_30_m_axi_gmem_RRESP;
	input qsort_30_m_axi_gmem_RLAST;
	input qsort_30_m_axi_gmem_RUSER;
	input qsort_30_m_axi_gmem_AWREADY;
	output wire qsort_30_m_axi_gmem_AWVALID;
	output wire qsort_30_m_axi_gmem_AWID;
	output wire [63:0] qsort_30_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_30_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_30_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_30_m_axi_gmem_AWBURST;
	output wire qsort_30_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_30_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_30_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_30_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_30_m_axi_gmem_AWREGION;
	output wire qsort_30_m_axi_gmem_AWUSER;
	input qsort_30_m_axi_gmem_WREADY;
	output wire qsort_30_m_axi_gmem_WVALID;
	output wire [63:0] qsort_30_m_axi_gmem_WDATA;
	output wire [7:0] qsort_30_m_axi_gmem_WSTRB;
	output wire qsort_30_m_axi_gmem_WLAST;
	output wire qsort_30_m_axi_gmem_WUSER;
	output wire qsort_30_m_axi_gmem_BREADY;
	input qsort_30_m_axi_gmem_BVALID;
	input qsort_30_m_axi_gmem_BID;
	input [1:0] qsort_30_m_axi_gmem_BRESP;
	input qsort_30_m_axi_gmem_BUSER;
	output wire qsort_30_s_axi_control_ARREADY;
	input qsort_30_s_axi_control_ARVALID;
	input [5:0] qsort_30_s_axi_control_ARADDR;
	input qsort_30_s_axi_control_RREADY;
	output wire qsort_30_s_axi_control_RVALID;
	output wire [31:0] qsort_30_s_axi_control_RDATA;
	output wire [1:0] qsort_30_s_axi_control_RRESP;
	output wire qsort_30_s_axi_control_AWREADY;
	input qsort_30_s_axi_control_AWVALID;
	input [5:0] qsort_30_s_axi_control_AWADDR;
	output wire qsort_30_s_axi_control_WREADY;
	input qsort_30_s_axi_control_WVALID;
	input [31:0] qsort_30_s_axi_control_WDATA;
	input [3:0] qsort_30_s_axi_control_WSTRB;
	input qsort_30_s_axi_control_BREADY;
	output wire qsort_30_s_axi_control_BVALID;
	output wire [1:0] qsort_30_s_axi_control_BRESP;
	input qsort_31_m_axi_gmem_ARREADY;
	output wire qsort_31_m_axi_gmem_ARVALID;
	output wire qsort_31_m_axi_gmem_ARID;
	output wire [63:0] qsort_31_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_31_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_31_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_31_m_axi_gmem_ARBURST;
	output wire qsort_31_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_31_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_31_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_31_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_31_m_axi_gmem_ARREGION;
	output wire qsort_31_m_axi_gmem_ARUSER;
	output wire qsort_31_m_axi_gmem_RREADY;
	input qsort_31_m_axi_gmem_RVALID;
	input qsort_31_m_axi_gmem_RID;
	input [63:0] qsort_31_m_axi_gmem_RDATA;
	input [1:0] qsort_31_m_axi_gmem_RRESP;
	input qsort_31_m_axi_gmem_RLAST;
	input qsort_31_m_axi_gmem_RUSER;
	input qsort_31_m_axi_gmem_AWREADY;
	output wire qsort_31_m_axi_gmem_AWVALID;
	output wire qsort_31_m_axi_gmem_AWID;
	output wire [63:0] qsort_31_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_31_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_31_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_31_m_axi_gmem_AWBURST;
	output wire qsort_31_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_31_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_31_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_31_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_31_m_axi_gmem_AWREGION;
	output wire qsort_31_m_axi_gmem_AWUSER;
	input qsort_31_m_axi_gmem_WREADY;
	output wire qsort_31_m_axi_gmem_WVALID;
	output wire [63:0] qsort_31_m_axi_gmem_WDATA;
	output wire [7:0] qsort_31_m_axi_gmem_WSTRB;
	output wire qsort_31_m_axi_gmem_WLAST;
	output wire qsort_31_m_axi_gmem_WUSER;
	output wire qsort_31_m_axi_gmem_BREADY;
	input qsort_31_m_axi_gmem_BVALID;
	input qsort_31_m_axi_gmem_BID;
	input [1:0] qsort_31_m_axi_gmem_BRESP;
	input qsort_31_m_axi_gmem_BUSER;
	output wire qsort_31_s_axi_control_ARREADY;
	input qsort_31_s_axi_control_ARVALID;
	input [5:0] qsort_31_s_axi_control_ARADDR;
	input qsort_31_s_axi_control_RREADY;
	output wire qsort_31_s_axi_control_RVALID;
	output wire [31:0] qsort_31_s_axi_control_RDATA;
	output wire [1:0] qsort_31_s_axi_control_RRESP;
	output wire qsort_31_s_axi_control_AWREADY;
	input qsort_31_s_axi_control_AWVALID;
	input [5:0] qsort_31_s_axi_control_AWADDR;
	output wire qsort_31_s_axi_control_WREADY;
	input qsort_31_s_axi_control_WVALID;
	input [31:0] qsort_31_s_axi_control_WDATA;
	input [3:0] qsort_31_s_axi_control_WSTRB;
	input qsort_31_s_axi_control_BREADY;
	output wire qsort_31_s_axi_control_BVALID;
	output wire [1:0] qsort_31_s_axi_control_BRESP;
	input qsort_32_m_axi_gmem_ARREADY;
	output wire qsort_32_m_axi_gmem_ARVALID;
	output wire qsort_32_m_axi_gmem_ARID;
	output wire [63:0] qsort_32_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_32_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_32_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_32_m_axi_gmem_ARBURST;
	output wire qsort_32_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_32_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_32_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_32_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_32_m_axi_gmem_ARREGION;
	output wire qsort_32_m_axi_gmem_ARUSER;
	output wire qsort_32_m_axi_gmem_RREADY;
	input qsort_32_m_axi_gmem_RVALID;
	input qsort_32_m_axi_gmem_RID;
	input [63:0] qsort_32_m_axi_gmem_RDATA;
	input [1:0] qsort_32_m_axi_gmem_RRESP;
	input qsort_32_m_axi_gmem_RLAST;
	input qsort_32_m_axi_gmem_RUSER;
	input qsort_32_m_axi_gmem_AWREADY;
	output wire qsort_32_m_axi_gmem_AWVALID;
	output wire qsort_32_m_axi_gmem_AWID;
	output wire [63:0] qsort_32_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_32_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_32_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_32_m_axi_gmem_AWBURST;
	output wire qsort_32_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_32_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_32_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_32_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_32_m_axi_gmem_AWREGION;
	output wire qsort_32_m_axi_gmem_AWUSER;
	input qsort_32_m_axi_gmem_WREADY;
	output wire qsort_32_m_axi_gmem_WVALID;
	output wire [63:0] qsort_32_m_axi_gmem_WDATA;
	output wire [7:0] qsort_32_m_axi_gmem_WSTRB;
	output wire qsort_32_m_axi_gmem_WLAST;
	output wire qsort_32_m_axi_gmem_WUSER;
	output wire qsort_32_m_axi_gmem_BREADY;
	input qsort_32_m_axi_gmem_BVALID;
	input qsort_32_m_axi_gmem_BID;
	input [1:0] qsort_32_m_axi_gmem_BRESP;
	input qsort_32_m_axi_gmem_BUSER;
	output wire qsort_32_s_axi_control_ARREADY;
	input qsort_32_s_axi_control_ARVALID;
	input [5:0] qsort_32_s_axi_control_ARADDR;
	input qsort_32_s_axi_control_RREADY;
	output wire qsort_32_s_axi_control_RVALID;
	output wire [31:0] qsort_32_s_axi_control_RDATA;
	output wire [1:0] qsort_32_s_axi_control_RRESP;
	output wire qsort_32_s_axi_control_AWREADY;
	input qsort_32_s_axi_control_AWVALID;
	input [5:0] qsort_32_s_axi_control_AWADDR;
	output wire qsort_32_s_axi_control_WREADY;
	input qsort_32_s_axi_control_WVALID;
	input [31:0] qsort_32_s_axi_control_WDATA;
	input [3:0] qsort_32_s_axi_control_WSTRB;
	input qsort_32_s_axi_control_BREADY;
	output wire qsort_32_s_axi_control_BVALID;
	output wire [1:0] qsort_32_s_axi_control_BRESP;
	input qsort_33_m_axi_gmem_ARREADY;
	output wire qsort_33_m_axi_gmem_ARVALID;
	output wire qsort_33_m_axi_gmem_ARID;
	output wire [63:0] qsort_33_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_33_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_33_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_33_m_axi_gmem_ARBURST;
	output wire qsort_33_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_33_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_33_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_33_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_33_m_axi_gmem_ARREGION;
	output wire qsort_33_m_axi_gmem_ARUSER;
	output wire qsort_33_m_axi_gmem_RREADY;
	input qsort_33_m_axi_gmem_RVALID;
	input qsort_33_m_axi_gmem_RID;
	input [63:0] qsort_33_m_axi_gmem_RDATA;
	input [1:0] qsort_33_m_axi_gmem_RRESP;
	input qsort_33_m_axi_gmem_RLAST;
	input qsort_33_m_axi_gmem_RUSER;
	input qsort_33_m_axi_gmem_AWREADY;
	output wire qsort_33_m_axi_gmem_AWVALID;
	output wire qsort_33_m_axi_gmem_AWID;
	output wire [63:0] qsort_33_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_33_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_33_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_33_m_axi_gmem_AWBURST;
	output wire qsort_33_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_33_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_33_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_33_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_33_m_axi_gmem_AWREGION;
	output wire qsort_33_m_axi_gmem_AWUSER;
	input qsort_33_m_axi_gmem_WREADY;
	output wire qsort_33_m_axi_gmem_WVALID;
	output wire [63:0] qsort_33_m_axi_gmem_WDATA;
	output wire [7:0] qsort_33_m_axi_gmem_WSTRB;
	output wire qsort_33_m_axi_gmem_WLAST;
	output wire qsort_33_m_axi_gmem_WUSER;
	output wire qsort_33_m_axi_gmem_BREADY;
	input qsort_33_m_axi_gmem_BVALID;
	input qsort_33_m_axi_gmem_BID;
	input [1:0] qsort_33_m_axi_gmem_BRESP;
	input qsort_33_m_axi_gmem_BUSER;
	output wire qsort_33_s_axi_control_ARREADY;
	input qsort_33_s_axi_control_ARVALID;
	input [5:0] qsort_33_s_axi_control_ARADDR;
	input qsort_33_s_axi_control_RREADY;
	output wire qsort_33_s_axi_control_RVALID;
	output wire [31:0] qsort_33_s_axi_control_RDATA;
	output wire [1:0] qsort_33_s_axi_control_RRESP;
	output wire qsort_33_s_axi_control_AWREADY;
	input qsort_33_s_axi_control_AWVALID;
	input [5:0] qsort_33_s_axi_control_AWADDR;
	output wire qsort_33_s_axi_control_WREADY;
	input qsort_33_s_axi_control_WVALID;
	input [31:0] qsort_33_s_axi_control_WDATA;
	input [3:0] qsort_33_s_axi_control_WSTRB;
	input qsort_33_s_axi_control_BREADY;
	output wire qsort_33_s_axi_control_BVALID;
	output wire [1:0] qsort_33_s_axi_control_BRESP;
	input qsort_34_m_axi_gmem_ARREADY;
	output wire qsort_34_m_axi_gmem_ARVALID;
	output wire qsort_34_m_axi_gmem_ARID;
	output wire [63:0] qsort_34_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_34_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_34_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_34_m_axi_gmem_ARBURST;
	output wire qsort_34_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_34_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_34_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_34_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_34_m_axi_gmem_ARREGION;
	output wire qsort_34_m_axi_gmem_ARUSER;
	output wire qsort_34_m_axi_gmem_RREADY;
	input qsort_34_m_axi_gmem_RVALID;
	input qsort_34_m_axi_gmem_RID;
	input [63:0] qsort_34_m_axi_gmem_RDATA;
	input [1:0] qsort_34_m_axi_gmem_RRESP;
	input qsort_34_m_axi_gmem_RLAST;
	input qsort_34_m_axi_gmem_RUSER;
	input qsort_34_m_axi_gmem_AWREADY;
	output wire qsort_34_m_axi_gmem_AWVALID;
	output wire qsort_34_m_axi_gmem_AWID;
	output wire [63:0] qsort_34_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_34_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_34_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_34_m_axi_gmem_AWBURST;
	output wire qsort_34_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_34_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_34_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_34_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_34_m_axi_gmem_AWREGION;
	output wire qsort_34_m_axi_gmem_AWUSER;
	input qsort_34_m_axi_gmem_WREADY;
	output wire qsort_34_m_axi_gmem_WVALID;
	output wire [63:0] qsort_34_m_axi_gmem_WDATA;
	output wire [7:0] qsort_34_m_axi_gmem_WSTRB;
	output wire qsort_34_m_axi_gmem_WLAST;
	output wire qsort_34_m_axi_gmem_WUSER;
	output wire qsort_34_m_axi_gmem_BREADY;
	input qsort_34_m_axi_gmem_BVALID;
	input qsort_34_m_axi_gmem_BID;
	input [1:0] qsort_34_m_axi_gmem_BRESP;
	input qsort_34_m_axi_gmem_BUSER;
	output wire qsort_34_s_axi_control_ARREADY;
	input qsort_34_s_axi_control_ARVALID;
	input [5:0] qsort_34_s_axi_control_ARADDR;
	input qsort_34_s_axi_control_RREADY;
	output wire qsort_34_s_axi_control_RVALID;
	output wire [31:0] qsort_34_s_axi_control_RDATA;
	output wire [1:0] qsort_34_s_axi_control_RRESP;
	output wire qsort_34_s_axi_control_AWREADY;
	input qsort_34_s_axi_control_AWVALID;
	input [5:0] qsort_34_s_axi_control_AWADDR;
	output wire qsort_34_s_axi_control_WREADY;
	input qsort_34_s_axi_control_WVALID;
	input [31:0] qsort_34_s_axi_control_WDATA;
	input [3:0] qsort_34_s_axi_control_WSTRB;
	input qsort_34_s_axi_control_BREADY;
	output wire qsort_34_s_axi_control_BVALID;
	output wire [1:0] qsort_34_s_axi_control_BRESP;
	input qsort_35_m_axi_gmem_ARREADY;
	output wire qsort_35_m_axi_gmem_ARVALID;
	output wire qsort_35_m_axi_gmem_ARID;
	output wire [63:0] qsort_35_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_35_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_35_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_35_m_axi_gmem_ARBURST;
	output wire qsort_35_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_35_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_35_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_35_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_35_m_axi_gmem_ARREGION;
	output wire qsort_35_m_axi_gmem_ARUSER;
	output wire qsort_35_m_axi_gmem_RREADY;
	input qsort_35_m_axi_gmem_RVALID;
	input qsort_35_m_axi_gmem_RID;
	input [63:0] qsort_35_m_axi_gmem_RDATA;
	input [1:0] qsort_35_m_axi_gmem_RRESP;
	input qsort_35_m_axi_gmem_RLAST;
	input qsort_35_m_axi_gmem_RUSER;
	input qsort_35_m_axi_gmem_AWREADY;
	output wire qsort_35_m_axi_gmem_AWVALID;
	output wire qsort_35_m_axi_gmem_AWID;
	output wire [63:0] qsort_35_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_35_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_35_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_35_m_axi_gmem_AWBURST;
	output wire qsort_35_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_35_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_35_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_35_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_35_m_axi_gmem_AWREGION;
	output wire qsort_35_m_axi_gmem_AWUSER;
	input qsort_35_m_axi_gmem_WREADY;
	output wire qsort_35_m_axi_gmem_WVALID;
	output wire [63:0] qsort_35_m_axi_gmem_WDATA;
	output wire [7:0] qsort_35_m_axi_gmem_WSTRB;
	output wire qsort_35_m_axi_gmem_WLAST;
	output wire qsort_35_m_axi_gmem_WUSER;
	output wire qsort_35_m_axi_gmem_BREADY;
	input qsort_35_m_axi_gmem_BVALID;
	input qsort_35_m_axi_gmem_BID;
	input [1:0] qsort_35_m_axi_gmem_BRESP;
	input qsort_35_m_axi_gmem_BUSER;
	output wire qsort_35_s_axi_control_ARREADY;
	input qsort_35_s_axi_control_ARVALID;
	input [5:0] qsort_35_s_axi_control_ARADDR;
	input qsort_35_s_axi_control_RREADY;
	output wire qsort_35_s_axi_control_RVALID;
	output wire [31:0] qsort_35_s_axi_control_RDATA;
	output wire [1:0] qsort_35_s_axi_control_RRESP;
	output wire qsort_35_s_axi_control_AWREADY;
	input qsort_35_s_axi_control_AWVALID;
	input [5:0] qsort_35_s_axi_control_AWADDR;
	output wire qsort_35_s_axi_control_WREADY;
	input qsort_35_s_axi_control_WVALID;
	input [31:0] qsort_35_s_axi_control_WDATA;
	input [3:0] qsort_35_s_axi_control_WSTRB;
	input qsort_35_s_axi_control_BREADY;
	output wire qsort_35_s_axi_control_BVALID;
	output wire [1:0] qsort_35_s_axi_control_BRESP;
	input qsort_36_m_axi_gmem_ARREADY;
	output wire qsort_36_m_axi_gmem_ARVALID;
	output wire qsort_36_m_axi_gmem_ARID;
	output wire [63:0] qsort_36_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_36_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_36_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_36_m_axi_gmem_ARBURST;
	output wire qsort_36_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_36_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_36_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_36_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_36_m_axi_gmem_ARREGION;
	output wire qsort_36_m_axi_gmem_ARUSER;
	output wire qsort_36_m_axi_gmem_RREADY;
	input qsort_36_m_axi_gmem_RVALID;
	input qsort_36_m_axi_gmem_RID;
	input [63:0] qsort_36_m_axi_gmem_RDATA;
	input [1:0] qsort_36_m_axi_gmem_RRESP;
	input qsort_36_m_axi_gmem_RLAST;
	input qsort_36_m_axi_gmem_RUSER;
	input qsort_36_m_axi_gmem_AWREADY;
	output wire qsort_36_m_axi_gmem_AWVALID;
	output wire qsort_36_m_axi_gmem_AWID;
	output wire [63:0] qsort_36_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_36_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_36_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_36_m_axi_gmem_AWBURST;
	output wire qsort_36_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_36_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_36_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_36_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_36_m_axi_gmem_AWREGION;
	output wire qsort_36_m_axi_gmem_AWUSER;
	input qsort_36_m_axi_gmem_WREADY;
	output wire qsort_36_m_axi_gmem_WVALID;
	output wire [63:0] qsort_36_m_axi_gmem_WDATA;
	output wire [7:0] qsort_36_m_axi_gmem_WSTRB;
	output wire qsort_36_m_axi_gmem_WLAST;
	output wire qsort_36_m_axi_gmem_WUSER;
	output wire qsort_36_m_axi_gmem_BREADY;
	input qsort_36_m_axi_gmem_BVALID;
	input qsort_36_m_axi_gmem_BID;
	input [1:0] qsort_36_m_axi_gmem_BRESP;
	input qsort_36_m_axi_gmem_BUSER;
	output wire qsort_36_s_axi_control_ARREADY;
	input qsort_36_s_axi_control_ARVALID;
	input [5:0] qsort_36_s_axi_control_ARADDR;
	input qsort_36_s_axi_control_RREADY;
	output wire qsort_36_s_axi_control_RVALID;
	output wire [31:0] qsort_36_s_axi_control_RDATA;
	output wire [1:0] qsort_36_s_axi_control_RRESP;
	output wire qsort_36_s_axi_control_AWREADY;
	input qsort_36_s_axi_control_AWVALID;
	input [5:0] qsort_36_s_axi_control_AWADDR;
	output wire qsort_36_s_axi_control_WREADY;
	input qsort_36_s_axi_control_WVALID;
	input [31:0] qsort_36_s_axi_control_WDATA;
	input [3:0] qsort_36_s_axi_control_WSTRB;
	input qsort_36_s_axi_control_BREADY;
	output wire qsort_36_s_axi_control_BVALID;
	output wire [1:0] qsort_36_s_axi_control_BRESP;
	input qsort_37_m_axi_gmem_ARREADY;
	output wire qsort_37_m_axi_gmem_ARVALID;
	output wire qsort_37_m_axi_gmem_ARID;
	output wire [63:0] qsort_37_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_37_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_37_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_37_m_axi_gmem_ARBURST;
	output wire qsort_37_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_37_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_37_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_37_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_37_m_axi_gmem_ARREGION;
	output wire qsort_37_m_axi_gmem_ARUSER;
	output wire qsort_37_m_axi_gmem_RREADY;
	input qsort_37_m_axi_gmem_RVALID;
	input qsort_37_m_axi_gmem_RID;
	input [63:0] qsort_37_m_axi_gmem_RDATA;
	input [1:0] qsort_37_m_axi_gmem_RRESP;
	input qsort_37_m_axi_gmem_RLAST;
	input qsort_37_m_axi_gmem_RUSER;
	input qsort_37_m_axi_gmem_AWREADY;
	output wire qsort_37_m_axi_gmem_AWVALID;
	output wire qsort_37_m_axi_gmem_AWID;
	output wire [63:0] qsort_37_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_37_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_37_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_37_m_axi_gmem_AWBURST;
	output wire qsort_37_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_37_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_37_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_37_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_37_m_axi_gmem_AWREGION;
	output wire qsort_37_m_axi_gmem_AWUSER;
	input qsort_37_m_axi_gmem_WREADY;
	output wire qsort_37_m_axi_gmem_WVALID;
	output wire [63:0] qsort_37_m_axi_gmem_WDATA;
	output wire [7:0] qsort_37_m_axi_gmem_WSTRB;
	output wire qsort_37_m_axi_gmem_WLAST;
	output wire qsort_37_m_axi_gmem_WUSER;
	output wire qsort_37_m_axi_gmem_BREADY;
	input qsort_37_m_axi_gmem_BVALID;
	input qsort_37_m_axi_gmem_BID;
	input [1:0] qsort_37_m_axi_gmem_BRESP;
	input qsort_37_m_axi_gmem_BUSER;
	output wire qsort_37_s_axi_control_ARREADY;
	input qsort_37_s_axi_control_ARVALID;
	input [5:0] qsort_37_s_axi_control_ARADDR;
	input qsort_37_s_axi_control_RREADY;
	output wire qsort_37_s_axi_control_RVALID;
	output wire [31:0] qsort_37_s_axi_control_RDATA;
	output wire [1:0] qsort_37_s_axi_control_RRESP;
	output wire qsort_37_s_axi_control_AWREADY;
	input qsort_37_s_axi_control_AWVALID;
	input [5:0] qsort_37_s_axi_control_AWADDR;
	output wire qsort_37_s_axi_control_WREADY;
	input qsort_37_s_axi_control_WVALID;
	input [31:0] qsort_37_s_axi_control_WDATA;
	input [3:0] qsort_37_s_axi_control_WSTRB;
	input qsort_37_s_axi_control_BREADY;
	output wire qsort_37_s_axi_control_BVALID;
	output wire [1:0] qsort_37_s_axi_control_BRESP;
	input qsort_38_m_axi_gmem_ARREADY;
	output wire qsort_38_m_axi_gmem_ARVALID;
	output wire qsort_38_m_axi_gmem_ARID;
	output wire [63:0] qsort_38_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_38_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_38_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_38_m_axi_gmem_ARBURST;
	output wire qsort_38_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_38_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_38_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_38_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_38_m_axi_gmem_ARREGION;
	output wire qsort_38_m_axi_gmem_ARUSER;
	output wire qsort_38_m_axi_gmem_RREADY;
	input qsort_38_m_axi_gmem_RVALID;
	input qsort_38_m_axi_gmem_RID;
	input [63:0] qsort_38_m_axi_gmem_RDATA;
	input [1:0] qsort_38_m_axi_gmem_RRESP;
	input qsort_38_m_axi_gmem_RLAST;
	input qsort_38_m_axi_gmem_RUSER;
	input qsort_38_m_axi_gmem_AWREADY;
	output wire qsort_38_m_axi_gmem_AWVALID;
	output wire qsort_38_m_axi_gmem_AWID;
	output wire [63:0] qsort_38_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_38_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_38_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_38_m_axi_gmem_AWBURST;
	output wire qsort_38_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_38_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_38_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_38_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_38_m_axi_gmem_AWREGION;
	output wire qsort_38_m_axi_gmem_AWUSER;
	input qsort_38_m_axi_gmem_WREADY;
	output wire qsort_38_m_axi_gmem_WVALID;
	output wire [63:0] qsort_38_m_axi_gmem_WDATA;
	output wire [7:0] qsort_38_m_axi_gmem_WSTRB;
	output wire qsort_38_m_axi_gmem_WLAST;
	output wire qsort_38_m_axi_gmem_WUSER;
	output wire qsort_38_m_axi_gmem_BREADY;
	input qsort_38_m_axi_gmem_BVALID;
	input qsort_38_m_axi_gmem_BID;
	input [1:0] qsort_38_m_axi_gmem_BRESP;
	input qsort_38_m_axi_gmem_BUSER;
	output wire qsort_38_s_axi_control_ARREADY;
	input qsort_38_s_axi_control_ARVALID;
	input [5:0] qsort_38_s_axi_control_ARADDR;
	input qsort_38_s_axi_control_RREADY;
	output wire qsort_38_s_axi_control_RVALID;
	output wire [31:0] qsort_38_s_axi_control_RDATA;
	output wire [1:0] qsort_38_s_axi_control_RRESP;
	output wire qsort_38_s_axi_control_AWREADY;
	input qsort_38_s_axi_control_AWVALID;
	input [5:0] qsort_38_s_axi_control_AWADDR;
	output wire qsort_38_s_axi_control_WREADY;
	input qsort_38_s_axi_control_WVALID;
	input [31:0] qsort_38_s_axi_control_WDATA;
	input [3:0] qsort_38_s_axi_control_WSTRB;
	input qsort_38_s_axi_control_BREADY;
	output wire qsort_38_s_axi_control_BVALID;
	output wire [1:0] qsort_38_s_axi_control_BRESP;
	input qsort_39_m_axi_gmem_ARREADY;
	output wire qsort_39_m_axi_gmem_ARVALID;
	output wire qsort_39_m_axi_gmem_ARID;
	output wire [63:0] qsort_39_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_39_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_39_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_39_m_axi_gmem_ARBURST;
	output wire qsort_39_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_39_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_39_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_39_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_39_m_axi_gmem_ARREGION;
	output wire qsort_39_m_axi_gmem_ARUSER;
	output wire qsort_39_m_axi_gmem_RREADY;
	input qsort_39_m_axi_gmem_RVALID;
	input qsort_39_m_axi_gmem_RID;
	input [63:0] qsort_39_m_axi_gmem_RDATA;
	input [1:0] qsort_39_m_axi_gmem_RRESP;
	input qsort_39_m_axi_gmem_RLAST;
	input qsort_39_m_axi_gmem_RUSER;
	input qsort_39_m_axi_gmem_AWREADY;
	output wire qsort_39_m_axi_gmem_AWVALID;
	output wire qsort_39_m_axi_gmem_AWID;
	output wire [63:0] qsort_39_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_39_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_39_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_39_m_axi_gmem_AWBURST;
	output wire qsort_39_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_39_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_39_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_39_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_39_m_axi_gmem_AWREGION;
	output wire qsort_39_m_axi_gmem_AWUSER;
	input qsort_39_m_axi_gmem_WREADY;
	output wire qsort_39_m_axi_gmem_WVALID;
	output wire [63:0] qsort_39_m_axi_gmem_WDATA;
	output wire [7:0] qsort_39_m_axi_gmem_WSTRB;
	output wire qsort_39_m_axi_gmem_WLAST;
	output wire qsort_39_m_axi_gmem_WUSER;
	output wire qsort_39_m_axi_gmem_BREADY;
	input qsort_39_m_axi_gmem_BVALID;
	input qsort_39_m_axi_gmem_BID;
	input [1:0] qsort_39_m_axi_gmem_BRESP;
	input qsort_39_m_axi_gmem_BUSER;
	output wire qsort_39_s_axi_control_ARREADY;
	input qsort_39_s_axi_control_ARVALID;
	input [5:0] qsort_39_s_axi_control_ARADDR;
	input qsort_39_s_axi_control_RREADY;
	output wire qsort_39_s_axi_control_RVALID;
	output wire [31:0] qsort_39_s_axi_control_RDATA;
	output wire [1:0] qsort_39_s_axi_control_RRESP;
	output wire qsort_39_s_axi_control_AWREADY;
	input qsort_39_s_axi_control_AWVALID;
	input [5:0] qsort_39_s_axi_control_AWADDR;
	output wire qsort_39_s_axi_control_WREADY;
	input qsort_39_s_axi_control_WVALID;
	input [31:0] qsort_39_s_axi_control_WDATA;
	input [3:0] qsort_39_s_axi_control_WSTRB;
	input qsort_39_s_axi_control_BREADY;
	output wire qsort_39_s_axi_control_BVALID;
	output wire [1:0] qsort_39_s_axi_control_BRESP;
	input qsort_40_m_axi_gmem_ARREADY;
	output wire qsort_40_m_axi_gmem_ARVALID;
	output wire qsort_40_m_axi_gmem_ARID;
	output wire [63:0] qsort_40_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_40_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_40_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_40_m_axi_gmem_ARBURST;
	output wire qsort_40_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_40_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_40_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_40_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_40_m_axi_gmem_ARREGION;
	output wire qsort_40_m_axi_gmem_ARUSER;
	output wire qsort_40_m_axi_gmem_RREADY;
	input qsort_40_m_axi_gmem_RVALID;
	input qsort_40_m_axi_gmem_RID;
	input [63:0] qsort_40_m_axi_gmem_RDATA;
	input [1:0] qsort_40_m_axi_gmem_RRESP;
	input qsort_40_m_axi_gmem_RLAST;
	input qsort_40_m_axi_gmem_RUSER;
	input qsort_40_m_axi_gmem_AWREADY;
	output wire qsort_40_m_axi_gmem_AWVALID;
	output wire qsort_40_m_axi_gmem_AWID;
	output wire [63:0] qsort_40_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_40_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_40_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_40_m_axi_gmem_AWBURST;
	output wire qsort_40_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_40_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_40_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_40_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_40_m_axi_gmem_AWREGION;
	output wire qsort_40_m_axi_gmem_AWUSER;
	input qsort_40_m_axi_gmem_WREADY;
	output wire qsort_40_m_axi_gmem_WVALID;
	output wire [63:0] qsort_40_m_axi_gmem_WDATA;
	output wire [7:0] qsort_40_m_axi_gmem_WSTRB;
	output wire qsort_40_m_axi_gmem_WLAST;
	output wire qsort_40_m_axi_gmem_WUSER;
	output wire qsort_40_m_axi_gmem_BREADY;
	input qsort_40_m_axi_gmem_BVALID;
	input qsort_40_m_axi_gmem_BID;
	input [1:0] qsort_40_m_axi_gmem_BRESP;
	input qsort_40_m_axi_gmem_BUSER;
	output wire qsort_40_s_axi_control_ARREADY;
	input qsort_40_s_axi_control_ARVALID;
	input [5:0] qsort_40_s_axi_control_ARADDR;
	input qsort_40_s_axi_control_RREADY;
	output wire qsort_40_s_axi_control_RVALID;
	output wire [31:0] qsort_40_s_axi_control_RDATA;
	output wire [1:0] qsort_40_s_axi_control_RRESP;
	output wire qsort_40_s_axi_control_AWREADY;
	input qsort_40_s_axi_control_AWVALID;
	input [5:0] qsort_40_s_axi_control_AWADDR;
	output wire qsort_40_s_axi_control_WREADY;
	input qsort_40_s_axi_control_WVALID;
	input [31:0] qsort_40_s_axi_control_WDATA;
	input [3:0] qsort_40_s_axi_control_WSTRB;
	input qsort_40_s_axi_control_BREADY;
	output wire qsort_40_s_axi_control_BVALID;
	output wire [1:0] qsort_40_s_axi_control_BRESP;
	input qsort_41_m_axi_gmem_ARREADY;
	output wire qsort_41_m_axi_gmem_ARVALID;
	output wire qsort_41_m_axi_gmem_ARID;
	output wire [63:0] qsort_41_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_41_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_41_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_41_m_axi_gmem_ARBURST;
	output wire qsort_41_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_41_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_41_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_41_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_41_m_axi_gmem_ARREGION;
	output wire qsort_41_m_axi_gmem_ARUSER;
	output wire qsort_41_m_axi_gmem_RREADY;
	input qsort_41_m_axi_gmem_RVALID;
	input qsort_41_m_axi_gmem_RID;
	input [63:0] qsort_41_m_axi_gmem_RDATA;
	input [1:0] qsort_41_m_axi_gmem_RRESP;
	input qsort_41_m_axi_gmem_RLAST;
	input qsort_41_m_axi_gmem_RUSER;
	input qsort_41_m_axi_gmem_AWREADY;
	output wire qsort_41_m_axi_gmem_AWVALID;
	output wire qsort_41_m_axi_gmem_AWID;
	output wire [63:0] qsort_41_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_41_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_41_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_41_m_axi_gmem_AWBURST;
	output wire qsort_41_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_41_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_41_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_41_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_41_m_axi_gmem_AWREGION;
	output wire qsort_41_m_axi_gmem_AWUSER;
	input qsort_41_m_axi_gmem_WREADY;
	output wire qsort_41_m_axi_gmem_WVALID;
	output wire [63:0] qsort_41_m_axi_gmem_WDATA;
	output wire [7:0] qsort_41_m_axi_gmem_WSTRB;
	output wire qsort_41_m_axi_gmem_WLAST;
	output wire qsort_41_m_axi_gmem_WUSER;
	output wire qsort_41_m_axi_gmem_BREADY;
	input qsort_41_m_axi_gmem_BVALID;
	input qsort_41_m_axi_gmem_BID;
	input [1:0] qsort_41_m_axi_gmem_BRESP;
	input qsort_41_m_axi_gmem_BUSER;
	output wire qsort_41_s_axi_control_ARREADY;
	input qsort_41_s_axi_control_ARVALID;
	input [5:0] qsort_41_s_axi_control_ARADDR;
	input qsort_41_s_axi_control_RREADY;
	output wire qsort_41_s_axi_control_RVALID;
	output wire [31:0] qsort_41_s_axi_control_RDATA;
	output wire [1:0] qsort_41_s_axi_control_RRESP;
	output wire qsort_41_s_axi_control_AWREADY;
	input qsort_41_s_axi_control_AWVALID;
	input [5:0] qsort_41_s_axi_control_AWADDR;
	output wire qsort_41_s_axi_control_WREADY;
	input qsort_41_s_axi_control_WVALID;
	input [31:0] qsort_41_s_axi_control_WDATA;
	input [3:0] qsort_41_s_axi_control_WSTRB;
	input qsort_41_s_axi_control_BREADY;
	output wire qsort_41_s_axi_control_BVALID;
	output wire [1:0] qsort_41_s_axi_control_BRESP;
	input qsort_42_m_axi_gmem_ARREADY;
	output wire qsort_42_m_axi_gmem_ARVALID;
	output wire qsort_42_m_axi_gmem_ARID;
	output wire [63:0] qsort_42_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_42_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_42_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_42_m_axi_gmem_ARBURST;
	output wire qsort_42_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_42_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_42_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_42_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_42_m_axi_gmem_ARREGION;
	output wire qsort_42_m_axi_gmem_ARUSER;
	output wire qsort_42_m_axi_gmem_RREADY;
	input qsort_42_m_axi_gmem_RVALID;
	input qsort_42_m_axi_gmem_RID;
	input [63:0] qsort_42_m_axi_gmem_RDATA;
	input [1:0] qsort_42_m_axi_gmem_RRESP;
	input qsort_42_m_axi_gmem_RLAST;
	input qsort_42_m_axi_gmem_RUSER;
	input qsort_42_m_axi_gmem_AWREADY;
	output wire qsort_42_m_axi_gmem_AWVALID;
	output wire qsort_42_m_axi_gmem_AWID;
	output wire [63:0] qsort_42_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_42_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_42_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_42_m_axi_gmem_AWBURST;
	output wire qsort_42_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_42_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_42_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_42_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_42_m_axi_gmem_AWREGION;
	output wire qsort_42_m_axi_gmem_AWUSER;
	input qsort_42_m_axi_gmem_WREADY;
	output wire qsort_42_m_axi_gmem_WVALID;
	output wire [63:0] qsort_42_m_axi_gmem_WDATA;
	output wire [7:0] qsort_42_m_axi_gmem_WSTRB;
	output wire qsort_42_m_axi_gmem_WLAST;
	output wire qsort_42_m_axi_gmem_WUSER;
	output wire qsort_42_m_axi_gmem_BREADY;
	input qsort_42_m_axi_gmem_BVALID;
	input qsort_42_m_axi_gmem_BID;
	input [1:0] qsort_42_m_axi_gmem_BRESP;
	input qsort_42_m_axi_gmem_BUSER;
	output wire qsort_42_s_axi_control_ARREADY;
	input qsort_42_s_axi_control_ARVALID;
	input [5:0] qsort_42_s_axi_control_ARADDR;
	input qsort_42_s_axi_control_RREADY;
	output wire qsort_42_s_axi_control_RVALID;
	output wire [31:0] qsort_42_s_axi_control_RDATA;
	output wire [1:0] qsort_42_s_axi_control_RRESP;
	output wire qsort_42_s_axi_control_AWREADY;
	input qsort_42_s_axi_control_AWVALID;
	input [5:0] qsort_42_s_axi_control_AWADDR;
	output wire qsort_42_s_axi_control_WREADY;
	input qsort_42_s_axi_control_WVALID;
	input [31:0] qsort_42_s_axi_control_WDATA;
	input [3:0] qsort_42_s_axi_control_WSTRB;
	input qsort_42_s_axi_control_BREADY;
	output wire qsort_42_s_axi_control_BVALID;
	output wire [1:0] qsort_42_s_axi_control_BRESP;
	input qsort_43_m_axi_gmem_ARREADY;
	output wire qsort_43_m_axi_gmem_ARVALID;
	output wire qsort_43_m_axi_gmem_ARID;
	output wire [63:0] qsort_43_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_43_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_43_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_43_m_axi_gmem_ARBURST;
	output wire qsort_43_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_43_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_43_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_43_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_43_m_axi_gmem_ARREGION;
	output wire qsort_43_m_axi_gmem_ARUSER;
	output wire qsort_43_m_axi_gmem_RREADY;
	input qsort_43_m_axi_gmem_RVALID;
	input qsort_43_m_axi_gmem_RID;
	input [63:0] qsort_43_m_axi_gmem_RDATA;
	input [1:0] qsort_43_m_axi_gmem_RRESP;
	input qsort_43_m_axi_gmem_RLAST;
	input qsort_43_m_axi_gmem_RUSER;
	input qsort_43_m_axi_gmem_AWREADY;
	output wire qsort_43_m_axi_gmem_AWVALID;
	output wire qsort_43_m_axi_gmem_AWID;
	output wire [63:0] qsort_43_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_43_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_43_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_43_m_axi_gmem_AWBURST;
	output wire qsort_43_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_43_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_43_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_43_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_43_m_axi_gmem_AWREGION;
	output wire qsort_43_m_axi_gmem_AWUSER;
	input qsort_43_m_axi_gmem_WREADY;
	output wire qsort_43_m_axi_gmem_WVALID;
	output wire [63:0] qsort_43_m_axi_gmem_WDATA;
	output wire [7:0] qsort_43_m_axi_gmem_WSTRB;
	output wire qsort_43_m_axi_gmem_WLAST;
	output wire qsort_43_m_axi_gmem_WUSER;
	output wire qsort_43_m_axi_gmem_BREADY;
	input qsort_43_m_axi_gmem_BVALID;
	input qsort_43_m_axi_gmem_BID;
	input [1:0] qsort_43_m_axi_gmem_BRESP;
	input qsort_43_m_axi_gmem_BUSER;
	output wire qsort_43_s_axi_control_ARREADY;
	input qsort_43_s_axi_control_ARVALID;
	input [5:0] qsort_43_s_axi_control_ARADDR;
	input qsort_43_s_axi_control_RREADY;
	output wire qsort_43_s_axi_control_RVALID;
	output wire [31:0] qsort_43_s_axi_control_RDATA;
	output wire [1:0] qsort_43_s_axi_control_RRESP;
	output wire qsort_43_s_axi_control_AWREADY;
	input qsort_43_s_axi_control_AWVALID;
	input [5:0] qsort_43_s_axi_control_AWADDR;
	output wire qsort_43_s_axi_control_WREADY;
	input qsort_43_s_axi_control_WVALID;
	input [31:0] qsort_43_s_axi_control_WDATA;
	input [3:0] qsort_43_s_axi_control_WSTRB;
	input qsort_43_s_axi_control_BREADY;
	output wire qsort_43_s_axi_control_BVALID;
	output wire [1:0] qsort_43_s_axi_control_BRESP;
	input qsort_44_m_axi_gmem_ARREADY;
	output wire qsort_44_m_axi_gmem_ARVALID;
	output wire qsort_44_m_axi_gmem_ARID;
	output wire [63:0] qsort_44_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_44_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_44_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_44_m_axi_gmem_ARBURST;
	output wire qsort_44_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_44_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_44_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_44_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_44_m_axi_gmem_ARREGION;
	output wire qsort_44_m_axi_gmem_ARUSER;
	output wire qsort_44_m_axi_gmem_RREADY;
	input qsort_44_m_axi_gmem_RVALID;
	input qsort_44_m_axi_gmem_RID;
	input [63:0] qsort_44_m_axi_gmem_RDATA;
	input [1:0] qsort_44_m_axi_gmem_RRESP;
	input qsort_44_m_axi_gmem_RLAST;
	input qsort_44_m_axi_gmem_RUSER;
	input qsort_44_m_axi_gmem_AWREADY;
	output wire qsort_44_m_axi_gmem_AWVALID;
	output wire qsort_44_m_axi_gmem_AWID;
	output wire [63:0] qsort_44_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_44_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_44_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_44_m_axi_gmem_AWBURST;
	output wire qsort_44_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_44_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_44_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_44_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_44_m_axi_gmem_AWREGION;
	output wire qsort_44_m_axi_gmem_AWUSER;
	input qsort_44_m_axi_gmem_WREADY;
	output wire qsort_44_m_axi_gmem_WVALID;
	output wire [63:0] qsort_44_m_axi_gmem_WDATA;
	output wire [7:0] qsort_44_m_axi_gmem_WSTRB;
	output wire qsort_44_m_axi_gmem_WLAST;
	output wire qsort_44_m_axi_gmem_WUSER;
	output wire qsort_44_m_axi_gmem_BREADY;
	input qsort_44_m_axi_gmem_BVALID;
	input qsort_44_m_axi_gmem_BID;
	input [1:0] qsort_44_m_axi_gmem_BRESP;
	input qsort_44_m_axi_gmem_BUSER;
	output wire qsort_44_s_axi_control_ARREADY;
	input qsort_44_s_axi_control_ARVALID;
	input [5:0] qsort_44_s_axi_control_ARADDR;
	input qsort_44_s_axi_control_RREADY;
	output wire qsort_44_s_axi_control_RVALID;
	output wire [31:0] qsort_44_s_axi_control_RDATA;
	output wire [1:0] qsort_44_s_axi_control_RRESP;
	output wire qsort_44_s_axi_control_AWREADY;
	input qsort_44_s_axi_control_AWVALID;
	input [5:0] qsort_44_s_axi_control_AWADDR;
	output wire qsort_44_s_axi_control_WREADY;
	input qsort_44_s_axi_control_WVALID;
	input [31:0] qsort_44_s_axi_control_WDATA;
	input [3:0] qsort_44_s_axi_control_WSTRB;
	input qsort_44_s_axi_control_BREADY;
	output wire qsort_44_s_axi_control_BVALID;
	output wire [1:0] qsort_44_s_axi_control_BRESP;
	input qsort_45_m_axi_gmem_ARREADY;
	output wire qsort_45_m_axi_gmem_ARVALID;
	output wire qsort_45_m_axi_gmem_ARID;
	output wire [63:0] qsort_45_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_45_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_45_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_45_m_axi_gmem_ARBURST;
	output wire qsort_45_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_45_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_45_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_45_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_45_m_axi_gmem_ARREGION;
	output wire qsort_45_m_axi_gmem_ARUSER;
	output wire qsort_45_m_axi_gmem_RREADY;
	input qsort_45_m_axi_gmem_RVALID;
	input qsort_45_m_axi_gmem_RID;
	input [63:0] qsort_45_m_axi_gmem_RDATA;
	input [1:0] qsort_45_m_axi_gmem_RRESP;
	input qsort_45_m_axi_gmem_RLAST;
	input qsort_45_m_axi_gmem_RUSER;
	input qsort_45_m_axi_gmem_AWREADY;
	output wire qsort_45_m_axi_gmem_AWVALID;
	output wire qsort_45_m_axi_gmem_AWID;
	output wire [63:0] qsort_45_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_45_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_45_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_45_m_axi_gmem_AWBURST;
	output wire qsort_45_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_45_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_45_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_45_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_45_m_axi_gmem_AWREGION;
	output wire qsort_45_m_axi_gmem_AWUSER;
	input qsort_45_m_axi_gmem_WREADY;
	output wire qsort_45_m_axi_gmem_WVALID;
	output wire [63:0] qsort_45_m_axi_gmem_WDATA;
	output wire [7:0] qsort_45_m_axi_gmem_WSTRB;
	output wire qsort_45_m_axi_gmem_WLAST;
	output wire qsort_45_m_axi_gmem_WUSER;
	output wire qsort_45_m_axi_gmem_BREADY;
	input qsort_45_m_axi_gmem_BVALID;
	input qsort_45_m_axi_gmem_BID;
	input [1:0] qsort_45_m_axi_gmem_BRESP;
	input qsort_45_m_axi_gmem_BUSER;
	output wire qsort_45_s_axi_control_ARREADY;
	input qsort_45_s_axi_control_ARVALID;
	input [5:0] qsort_45_s_axi_control_ARADDR;
	input qsort_45_s_axi_control_RREADY;
	output wire qsort_45_s_axi_control_RVALID;
	output wire [31:0] qsort_45_s_axi_control_RDATA;
	output wire [1:0] qsort_45_s_axi_control_RRESP;
	output wire qsort_45_s_axi_control_AWREADY;
	input qsort_45_s_axi_control_AWVALID;
	input [5:0] qsort_45_s_axi_control_AWADDR;
	output wire qsort_45_s_axi_control_WREADY;
	input qsort_45_s_axi_control_WVALID;
	input [31:0] qsort_45_s_axi_control_WDATA;
	input [3:0] qsort_45_s_axi_control_WSTRB;
	input qsort_45_s_axi_control_BREADY;
	output wire qsort_45_s_axi_control_BVALID;
	output wire [1:0] qsort_45_s_axi_control_BRESP;
	input qsort_46_m_axi_gmem_ARREADY;
	output wire qsort_46_m_axi_gmem_ARVALID;
	output wire qsort_46_m_axi_gmem_ARID;
	output wire [63:0] qsort_46_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_46_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_46_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_46_m_axi_gmem_ARBURST;
	output wire qsort_46_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_46_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_46_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_46_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_46_m_axi_gmem_ARREGION;
	output wire qsort_46_m_axi_gmem_ARUSER;
	output wire qsort_46_m_axi_gmem_RREADY;
	input qsort_46_m_axi_gmem_RVALID;
	input qsort_46_m_axi_gmem_RID;
	input [63:0] qsort_46_m_axi_gmem_RDATA;
	input [1:0] qsort_46_m_axi_gmem_RRESP;
	input qsort_46_m_axi_gmem_RLAST;
	input qsort_46_m_axi_gmem_RUSER;
	input qsort_46_m_axi_gmem_AWREADY;
	output wire qsort_46_m_axi_gmem_AWVALID;
	output wire qsort_46_m_axi_gmem_AWID;
	output wire [63:0] qsort_46_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_46_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_46_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_46_m_axi_gmem_AWBURST;
	output wire qsort_46_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_46_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_46_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_46_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_46_m_axi_gmem_AWREGION;
	output wire qsort_46_m_axi_gmem_AWUSER;
	input qsort_46_m_axi_gmem_WREADY;
	output wire qsort_46_m_axi_gmem_WVALID;
	output wire [63:0] qsort_46_m_axi_gmem_WDATA;
	output wire [7:0] qsort_46_m_axi_gmem_WSTRB;
	output wire qsort_46_m_axi_gmem_WLAST;
	output wire qsort_46_m_axi_gmem_WUSER;
	output wire qsort_46_m_axi_gmem_BREADY;
	input qsort_46_m_axi_gmem_BVALID;
	input qsort_46_m_axi_gmem_BID;
	input [1:0] qsort_46_m_axi_gmem_BRESP;
	input qsort_46_m_axi_gmem_BUSER;
	output wire qsort_46_s_axi_control_ARREADY;
	input qsort_46_s_axi_control_ARVALID;
	input [5:0] qsort_46_s_axi_control_ARADDR;
	input qsort_46_s_axi_control_RREADY;
	output wire qsort_46_s_axi_control_RVALID;
	output wire [31:0] qsort_46_s_axi_control_RDATA;
	output wire [1:0] qsort_46_s_axi_control_RRESP;
	output wire qsort_46_s_axi_control_AWREADY;
	input qsort_46_s_axi_control_AWVALID;
	input [5:0] qsort_46_s_axi_control_AWADDR;
	output wire qsort_46_s_axi_control_WREADY;
	input qsort_46_s_axi_control_WVALID;
	input [31:0] qsort_46_s_axi_control_WDATA;
	input [3:0] qsort_46_s_axi_control_WSTRB;
	input qsort_46_s_axi_control_BREADY;
	output wire qsort_46_s_axi_control_BVALID;
	output wire [1:0] qsort_46_s_axi_control_BRESP;
	input qsort_47_m_axi_gmem_ARREADY;
	output wire qsort_47_m_axi_gmem_ARVALID;
	output wire qsort_47_m_axi_gmem_ARID;
	output wire [63:0] qsort_47_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_47_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_47_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_47_m_axi_gmem_ARBURST;
	output wire qsort_47_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_47_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_47_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_47_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_47_m_axi_gmem_ARREGION;
	output wire qsort_47_m_axi_gmem_ARUSER;
	output wire qsort_47_m_axi_gmem_RREADY;
	input qsort_47_m_axi_gmem_RVALID;
	input qsort_47_m_axi_gmem_RID;
	input [63:0] qsort_47_m_axi_gmem_RDATA;
	input [1:0] qsort_47_m_axi_gmem_RRESP;
	input qsort_47_m_axi_gmem_RLAST;
	input qsort_47_m_axi_gmem_RUSER;
	input qsort_47_m_axi_gmem_AWREADY;
	output wire qsort_47_m_axi_gmem_AWVALID;
	output wire qsort_47_m_axi_gmem_AWID;
	output wire [63:0] qsort_47_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_47_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_47_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_47_m_axi_gmem_AWBURST;
	output wire qsort_47_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_47_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_47_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_47_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_47_m_axi_gmem_AWREGION;
	output wire qsort_47_m_axi_gmem_AWUSER;
	input qsort_47_m_axi_gmem_WREADY;
	output wire qsort_47_m_axi_gmem_WVALID;
	output wire [63:0] qsort_47_m_axi_gmem_WDATA;
	output wire [7:0] qsort_47_m_axi_gmem_WSTRB;
	output wire qsort_47_m_axi_gmem_WLAST;
	output wire qsort_47_m_axi_gmem_WUSER;
	output wire qsort_47_m_axi_gmem_BREADY;
	input qsort_47_m_axi_gmem_BVALID;
	input qsort_47_m_axi_gmem_BID;
	input [1:0] qsort_47_m_axi_gmem_BRESP;
	input qsort_47_m_axi_gmem_BUSER;
	output wire qsort_47_s_axi_control_ARREADY;
	input qsort_47_s_axi_control_ARVALID;
	input [5:0] qsort_47_s_axi_control_ARADDR;
	input qsort_47_s_axi_control_RREADY;
	output wire qsort_47_s_axi_control_RVALID;
	output wire [31:0] qsort_47_s_axi_control_RDATA;
	output wire [1:0] qsort_47_s_axi_control_RRESP;
	output wire qsort_47_s_axi_control_AWREADY;
	input qsort_47_s_axi_control_AWVALID;
	input [5:0] qsort_47_s_axi_control_AWADDR;
	output wire qsort_47_s_axi_control_WREADY;
	input qsort_47_s_axi_control_WVALID;
	input [31:0] qsort_47_s_axi_control_WDATA;
	input [3:0] qsort_47_s_axi_control_WSTRB;
	input qsort_47_s_axi_control_BREADY;
	output wire qsort_47_s_axi_control_BVALID;
	output wire [1:0] qsort_47_s_axi_control_BRESP;
	input qsort_48_m_axi_gmem_ARREADY;
	output wire qsort_48_m_axi_gmem_ARVALID;
	output wire qsort_48_m_axi_gmem_ARID;
	output wire [63:0] qsort_48_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_48_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_48_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_48_m_axi_gmem_ARBURST;
	output wire qsort_48_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_48_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_48_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_48_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_48_m_axi_gmem_ARREGION;
	output wire qsort_48_m_axi_gmem_ARUSER;
	output wire qsort_48_m_axi_gmem_RREADY;
	input qsort_48_m_axi_gmem_RVALID;
	input qsort_48_m_axi_gmem_RID;
	input [63:0] qsort_48_m_axi_gmem_RDATA;
	input [1:0] qsort_48_m_axi_gmem_RRESP;
	input qsort_48_m_axi_gmem_RLAST;
	input qsort_48_m_axi_gmem_RUSER;
	input qsort_48_m_axi_gmem_AWREADY;
	output wire qsort_48_m_axi_gmem_AWVALID;
	output wire qsort_48_m_axi_gmem_AWID;
	output wire [63:0] qsort_48_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_48_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_48_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_48_m_axi_gmem_AWBURST;
	output wire qsort_48_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_48_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_48_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_48_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_48_m_axi_gmem_AWREGION;
	output wire qsort_48_m_axi_gmem_AWUSER;
	input qsort_48_m_axi_gmem_WREADY;
	output wire qsort_48_m_axi_gmem_WVALID;
	output wire [63:0] qsort_48_m_axi_gmem_WDATA;
	output wire [7:0] qsort_48_m_axi_gmem_WSTRB;
	output wire qsort_48_m_axi_gmem_WLAST;
	output wire qsort_48_m_axi_gmem_WUSER;
	output wire qsort_48_m_axi_gmem_BREADY;
	input qsort_48_m_axi_gmem_BVALID;
	input qsort_48_m_axi_gmem_BID;
	input [1:0] qsort_48_m_axi_gmem_BRESP;
	input qsort_48_m_axi_gmem_BUSER;
	output wire qsort_48_s_axi_control_ARREADY;
	input qsort_48_s_axi_control_ARVALID;
	input [5:0] qsort_48_s_axi_control_ARADDR;
	input qsort_48_s_axi_control_RREADY;
	output wire qsort_48_s_axi_control_RVALID;
	output wire [31:0] qsort_48_s_axi_control_RDATA;
	output wire [1:0] qsort_48_s_axi_control_RRESP;
	output wire qsort_48_s_axi_control_AWREADY;
	input qsort_48_s_axi_control_AWVALID;
	input [5:0] qsort_48_s_axi_control_AWADDR;
	output wire qsort_48_s_axi_control_WREADY;
	input qsort_48_s_axi_control_WVALID;
	input [31:0] qsort_48_s_axi_control_WDATA;
	input [3:0] qsort_48_s_axi_control_WSTRB;
	input qsort_48_s_axi_control_BREADY;
	output wire qsort_48_s_axi_control_BVALID;
	output wire [1:0] qsort_48_s_axi_control_BRESP;
	input qsort_49_m_axi_gmem_ARREADY;
	output wire qsort_49_m_axi_gmem_ARVALID;
	output wire qsort_49_m_axi_gmem_ARID;
	output wire [63:0] qsort_49_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_49_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_49_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_49_m_axi_gmem_ARBURST;
	output wire qsort_49_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_49_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_49_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_49_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_49_m_axi_gmem_ARREGION;
	output wire qsort_49_m_axi_gmem_ARUSER;
	output wire qsort_49_m_axi_gmem_RREADY;
	input qsort_49_m_axi_gmem_RVALID;
	input qsort_49_m_axi_gmem_RID;
	input [63:0] qsort_49_m_axi_gmem_RDATA;
	input [1:0] qsort_49_m_axi_gmem_RRESP;
	input qsort_49_m_axi_gmem_RLAST;
	input qsort_49_m_axi_gmem_RUSER;
	input qsort_49_m_axi_gmem_AWREADY;
	output wire qsort_49_m_axi_gmem_AWVALID;
	output wire qsort_49_m_axi_gmem_AWID;
	output wire [63:0] qsort_49_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_49_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_49_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_49_m_axi_gmem_AWBURST;
	output wire qsort_49_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_49_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_49_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_49_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_49_m_axi_gmem_AWREGION;
	output wire qsort_49_m_axi_gmem_AWUSER;
	input qsort_49_m_axi_gmem_WREADY;
	output wire qsort_49_m_axi_gmem_WVALID;
	output wire [63:0] qsort_49_m_axi_gmem_WDATA;
	output wire [7:0] qsort_49_m_axi_gmem_WSTRB;
	output wire qsort_49_m_axi_gmem_WLAST;
	output wire qsort_49_m_axi_gmem_WUSER;
	output wire qsort_49_m_axi_gmem_BREADY;
	input qsort_49_m_axi_gmem_BVALID;
	input qsort_49_m_axi_gmem_BID;
	input [1:0] qsort_49_m_axi_gmem_BRESP;
	input qsort_49_m_axi_gmem_BUSER;
	output wire qsort_49_s_axi_control_ARREADY;
	input qsort_49_s_axi_control_ARVALID;
	input [5:0] qsort_49_s_axi_control_ARADDR;
	input qsort_49_s_axi_control_RREADY;
	output wire qsort_49_s_axi_control_RVALID;
	output wire [31:0] qsort_49_s_axi_control_RDATA;
	output wire [1:0] qsort_49_s_axi_control_RRESP;
	output wire qsort_49_s_axi_control_AWREADY;
	input qsort_49_s_axi_control_AWVALID;
	input [5:0] qsort_49_s_axi_control_AWADDR;
	output wire qsort_49_s_axi_control_WREADY;
	input qsort_49_s_axi_control_WVALID;
	input [31:0] qsort_49_s_axi_control_WDATA;
	input [3:0] qsort_49_s_axi_control_WSTRB;
	input qsort_49_s_axi_control_BREADY;
	output wire qsort_49_s_axi_control_BVALID;
	output wire [1:0] qsort_49_s_axi_control_BRESP;
	input qsort_50_m_axi_gmem_ARREADY;
	output wire qsort_50_m_axi_gmem_ARVALID;
	output wire qsort_50_m_axi_gmem_ARID;
	output wire [63:0] qsort_50_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_50_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_50_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_50_m_axi_gmem_ARBURST;
	output wire qsort_50_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_50_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_50_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_50_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_50_m_axi_gmem_ARREGION;
	output wire qsort_50_m_axi_gmem_ARUSER;
	output wire qsort_50_m_axi_gmem_RREADY;
	input qsort_50_m_axi_gmem_RVALID;
	input qsort_50_m_axi_gmem_RID;
	input [63:0] qsort_50_m_axi_gmem_RDATA;
	input [1:0] qsort_50_m_axi_gmem_RRESP;
	input qsort_50_m_axi_gmem_RLAST;
	input qsort_50_m_axi_gmem_RUSER;
	input qsort_50_m_axi_gmem_AWREADY;
	output wire qsort_50_m_axi_gmem_AWVALID;
	output wire qsort_50_m_axi_gmem_AWID;
	output wire [63:0] qsort_50_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_50_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_50_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_50_m_axi_gmem_AWBURST;
	output wire qsort_50_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_50_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_50_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_50_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_50_m_axi_gmem_AWREGION;
	output wire qsort_50_m_axi_gmem_AWUSER;
	input qsort_50_m_axi_gmem_WREADY;
	output wire qsort_50_m_axi_gmem_WVALID;
	output wire [63:0] qsort_50_m_axi_gmem_WDATA;
	output wire [7:0] qsort_50_m_axi_gmem_WSTRB;
	output wire qsort_50_m_axi_gmem_WLAST;
	output wire qsort_50_m_axi_gmem_WUSER;
	output wire qsort_50_m_axi_gmem_BREADY;
	input qsort_50_m_axi_gmem_BVALID;
	input qsort_50_m_axi_gmem_BID;
	input [1:0] qsort_50_m_axi_gmem_BRESP;
	input qsort_50_m_axi_gmem_BUSER;
	output wire qsort_50_s_axi_control_ARREADY;
	input qsort_50_s_axi_control_ARVALID;
	input [5:0] qsort_50_s_axi_control_ARADDR;
	input qsort_50_s_axi_control_RREADY;
	output wire qsort_50_s_axi_control_RVALID;
	output wire [31:0] qsort_50_s_axi_control_RDATA;
	output wire [1:0] qsort_50_s_axi_control_RRESP;
	output wire qsort_50_s_axi_control_AWREADY;
	input qsort_50_s_axi_control_AWVALID;
	input [5:0] qsort_50_s_axi_control_AWADDR;
	output wire qsort_50_s_axi_control_WREADY;
	input qsort_50_s_axi_control_WVALID;
	input [31:0] qsort_50_s_axi_control_WDATA;
	input [3:0] qsort_50_s_axi_control_WSTRB;
	input qsort_50_s_axi_control_BREADY;
	output wire qsort_50_s_axi_control_BVALID;
	output wire [1:0] qsort_50_s_axi_control_BRESP;
	input qsort_51_m_axi_gmem_ARREADY;
	output wire qsort_51_m_axi_gmem_ARVALID;
	output wire qsort_51_m_axi_gmem_ARID;
	output wire [63:0] qsort_51_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_51_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_51_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_51_m_axi_gmem_ARBURST;
	output wire qsort_51_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_51_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_51_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_51_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_51_m_axi_gmem_ARREGION;
	output wire qsort_51_m_axi_gmem_ARUSER;
	output wire qsort_51_m_axi_gmem_RREADY;
	input qsort_51_m_axi_gmem_RVALID;
	input qsort_51_m_axi_gmem_RID;
	input [63:0] qsort_51_m_axi_gmem_RDATA;
	input [1:0] qsort_51_m_axi_gmem_RRESP;
	input qsort_51_m_axi_gmem_RLAST;
	input qsort_51_m_axi_gmem_RUSER;
	input qsort_51_m_axi_gmem_AWREADY;
	output wire qsort_51_m_axi_gmem_AWVALID;
	output wire qsort_51_m_axi_gmem_AWID;
	output wire [63:0] qsort_51_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_51_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_51_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_51_m_axi_gmem_AWBURST;
	output wire qsort_51_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_51_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_51_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_51_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_51_m_axi_gmem_AWREGION;
	output wire qsort_51_m_axi_gmem_AWUSER;
	input qsort_51_m_axi_gmem_WREADY;
	output wire qsort_51_m_axi_gmem_WVALID;
	output wire [63:0] qsort_51_m_axi_gmem_WDATA;
	output wire [7:0] qsort_51_m_axi_gmem_WSTRB;
	output wire qsort_51_m_axi_gmem_WLAST;
	output wire qsort_51_m_axi_gmem_WUSER;
	output wire qsort_51_m_axi_gmem_BREADY;
	input qsort_51_m_axi_gmem_BVALID;
	input qsort_51_m_axi_gmem_BID;
	input [1:0] qsort_51_m_axi_gmem_BRESP;
	input qsort_51_m_axi_gmem_BUSER;
	output wire qsort_51_s_axi_control_ARREADY;
	input qsort_51_s_axi_control_ARVALID;
	input [5:0] qsort_51_s_axi_control_ARADDR;
	input qsort_51_s_axi_control_RREADY;
	output wire qsort_51_s_axi_control_RVALID;
	output wire [31:0] qsort_51_s_axi_control_RDATA;
	output wire [1:0] qsort_51_s_axi_control_RRESP;
	output wire qsort_51_s_axi_control_AWREADY;
	input qsort_51_s_axi_control_AWVALID;
	input [5:0] qsort_51_s_axi_control_AWADDR;
	output wire qsort_51_s_axi_control_WREADY;
	input qsort_51_s_axi_control_WVALID;
	input [31:0] qsort_51_s_axi_control_WDATA;
	input [3:0] qsort_51_s_axi_control_WSTRB;
	input qsort_51_s_axi_control_BREADY;
	output wire qsort_51_s_axi_control_BVALID;
	output wire [1:0] qsort_51_s_axi_control_BRESP;
	input qsort_52_m_axi_gmem_ARREADY;
	output wire qsort_52_m_axi_gmem_ARVALID;
	output wire qsort_52_m_axi_gmem_ARID;
	output wire [63:0] qsort_52_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_52_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_52_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_52_m_axi_gmem_ARBURST;
	output wire qsort_52_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_52_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_52_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_52_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_52_m_axi_gmem_ARREGION;
	output wire qsort_52_m_axi_gmem_ARUSER;
	output wire qsort_52_m_axi_gmem_RREADY;
	input qsort_52_m_axi_gmem_RVALID;
	input qsort_52_m_axi_gmem_RID;
	input [63:0] qsort_52_m_axi_gmem_RDATA;
	input [1:0] qsort_52_m_axi_gmem_RRESP;
	input qsort_52_m_axi_gmem_RLAST;
	input qsort_52_m_axi_gmem_RUSER;
	input qsort_52_m_axi_gmem_AWREADY;
	output wire qsort_52_m_axi_gmem_AWVALID;
	output wire qsort_52_m_axi_gmem_AWID;
	output wire [63:0] qsort_52_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_52_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_52_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_52_m_axi_gmem_AWBURST;
	output wire qsort_52_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_52_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_52_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_52_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_52_m_axi_gmem_AWREGION;
	output wire qsort_52_m_axi_gmem_AWUSER;
	input qsort_52_m_axi_gmem_WREADY;
	output wire qsort_52_m_axi_gmem_WVALID;
	output wire [63:0] qsort_52_m_axi_gmem_WDATA;
	output wire [7:0] qsort_52_m_axi_gmem_WSTRB;
	output wire qsort_52_m_axi_gmem_WLAST;
	output wire qsort_52_m_axi_gmem_WUSER;
	output wire qsort_52_m_axi_gmem_BREADY;
	input qsort_52_m_axi_gmem_BVALID;
	input qsort_52_m_axi_gmem_BID;
	input [1:0] qsort_52_m_axi_gmem_BRESP;
	input qsort_52_m_axi_gmem_BUSER;
	output wire qsort_52_s_axi_control_ARREADY;
	input qsort_52_s_axi_control_ARVALID;
	input [5:0] qsort_52_s_axi_control_ARADDR;
	input qsort_52_s_axi_control_RREADY;
	output wire qsort_52_s_axi_control_RVALID;
	output wire [31:0] qsort_52_s_axi_control_RDATA;
	output wire [1:0] qsort_52_s_axi_control_RRESP;
	output wire qsort_52_s_axi_control_AWREADY;
	input qsort_52_s_axi_control_AWVALID;
	input [5:0] qsort_52_s_axi_control_AWADDR;
	output wire qsort_52_s_axi_control_WREADY;
	input qsort_52_s_axi_control_WVALID;
	input [31:0] qsort_52_s_axi_control_WDATA;
	input [3:0] qsort_52_s_axi_control_WSTRB;
	input qsort_52_s_axi_control_BREADY;
	output wire qsort_52_s_axi_control_BVALID;
	output wire [1:0] qsort_52_s_axi_control_BRESP;
	input qsort_53_m_axi_gmem_ARREADY;
	output wire qsort_53_m_axi_gmem_ARVALID;
	output wire qsort_53_m_axi_gmem_ARID;
	output wire [63:0] qsort_53_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_53_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_53_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_53_m_axi_gmem_ARBURST;
	output wire qsort_53_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_53_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_53_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_53_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_53_m_axi_gmem_ARREGION;
	output wire qsort_53_m_axi_gmem_ARUSER;
	output wire qsort_53_m_axi_gmem_RREADY;
	input qsort_53_m_axi_gmem_RVALID;
	input qsort_53_m_axi_gmem_RID;
	input [63:0] qsort_53_m_axi_gmem_RDATA;
	input [1:0] qsort_53_m_axi_gmem_RRESP;
	input qsort_53_m_axi_gmem_RLAST;
	input qsort_53_m_axi_gmem_RUSER;
	input qsort_53_m_axi_gmem_AWREADY;
	output wire qsort_53_m_axi_gmem_AWVALID;
	output wire qsort_53_m_axi_gmem_AWID;
	output wire [63:0] qsort_53_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_53_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_53_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_53_m_axi_gmem_AWBURST;
	output wire qsort_53_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_53_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_53_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_53_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_53_m_axi_gmem_AWREGION;
	output wire qsort_53_m_axi_gmem_AWUSER;
	input qsort_53_m_axi_gmem_WREADY;
	output wire qsort_53_m_axi_gmem_WVALID;
	output wire [63:0] qsort_53_m_axi_gmem_WDATA;
	output wire [7:0] qsort_53_m_axi_gmem_WSTRB;
	output wire qsort_53_m_axi_gmem_WLAST;
	output wire qsort_53_m_axi_gmem_WUSER;
	output wire qsort_53_m_axi_gmem_BREADY;
	input qsort_53_m_axi_gmem_BVALID;
	input qsort_53_m_axi_gmem_BID;
	input [1:0] qsort_53_m_axi_gmem_BRESP;
	input qsort_53_m_axi_gmem_BUSER;
	output wire qsort_53_s_axi_control_ARREADY;
	input qsort_53_s_axi_control_ARVALID;
	input [5:0] qsort_53_s_axi_control_ARADDR;
	input qsort_53_s_axi_control_RREADY;
	output wire qsort_53_s_axi_control_RVALID;
	output wire [31:0] qsort_53_s_axi_control_RDATA;
	output wire [1:0] qsort_53_s_axi_control_RRESP;
	output wire qsort_53_s_axi_control_AWREADY;
	input qsort_53_s_axi_control_AWVALID;
	input [5:0] qsort_53_s_axi_control_AWADDR;
	output wire qsort_53_s_axi_control_WREADY;
	input qsort_53_s_axi_control_WVALID;
	input [31:0] qsort_53_s_axi_control_WDATA;
	input [3:0] qsort_53_s_axi_control_WSTRB;
	input qsort_53_s_axi_control_BREADY;
	output wire qsort_53_s_axi_control_BVALID;
	output wire [1:0] qsort_53_s_axi_control_BRESP;
	input qsort_54_m_axi_gmem_ARREADY;
	output wire qsort_54_m_axi_gmem_ARVALID;
	output wire qsort_54_m_axi_gmem_ARID;
	output wire [63:0] qsort_54_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_54_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_54_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_54_m_axi_gmem_ARBURST;
	output wire qsort_54_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_54_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_54_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_54_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_54_m_axi_gmem_ARREGION;
	output wire qsort_54_m_axi_gmem_ARUSER;
	output wire qsort_54_m_axi_gmem_RREADY;
	input qsort_54_m_axi_gmem_RVALID;
	input qsort_54_m_axi_gmem_RID;
	input [63:0] qsort_54_m_axi_gmem_RDATA;
	input [1:0] qsort_54_m_axi_gmem_RRESP;
	input qsort_54_m_axi_gmem_RLAST;
	input qsort_54_m_axi_gmem_RUSER;
	input qsort_54_m_axi_gmem_AWREADY;
	output wire qsort_54_m_axi_gmem_AWVALID;
	output wire qsort_54_m_axi_gmem_AWID;
	output wire [63:0] qsort_54_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_54_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_54_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_54_m_axi_gmem_AWBURST;
	output wire qsort_54_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_54_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_54_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_54_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_54_m_axi_gmem_AWREGION;
	output wire qsort_54_m_axi_gmem_AWUSER;
	input qsort_54_m_axi_gmem_WREADY;
	output wire qsort_54_m_axi_gmem_WVALID;
	output wire [63:0] qsort_54_m_axi_gmem_WDATA;
	output wire [7:0] qsort_54_m_axi_gmem_WSTRB;
	output wire qsort_54_m_axi_gmem_WLAST;
	output wire qsort_54_m_axi_gmem_WUSER;
	output wire qsort_54_m_axi_gmem_BREADY;
	input qsort_54_m_axi_gmem_BVALID;
	input qsort_54_m_axi_gmem_BID;
	input [1:0] qsort_54_m_axi_gmem_BRESP;
	input qsort_54_m_axi_gmem_BUSER;
	output wire qsort_54_s_axi_control_ARREADY;
	input qsort_54_s_axi_control_ARVALID;
	input [5:0] qsort_54_s_axi_control_ARADDR;
	input qsort_54_s_axi_control_RREADY;
	output wire qsort_54_s_axi_control_RVALID;
	output wire [31:0] qsort_54_s_axi_control_RDATA;
	output wire [1:0] qsort_54_s_axi_control_RRESP;
	output wire qsort_54_s_axi_control_AWREADY;
	input qsort_54_s_axi_control_AWVALID;
	input [5:0] qsort_54_s_axi_control_AWADDR;
	output wire qsort_54_s_axi_control_WREADY;
	input qsort_54_s_axi_control_WVALID;
	input [31:0] qsort_54_s_axi_control_WDATA;
	input [3:0] qsort_54_s_axi_control_WSTRB;
	input qsort_54_s_axi_control_BREADY;
	output wire qsort_54_s_axi_control_BVALID;
	output wire [1:0] qsort_54_s_axi_control_BRESP;
	input qsort_55_m_axi_gmem_ARREADY;
	output wire qsort_55_m_axi_gmem_ARVALID;
	output wire qsort_55_m_axi_gmem_ARID;
	output wire [63:0] qsort_55_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_55_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_55_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_55_m_axi_gmem_ARBURST;
	output wire qsort_55_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_55_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_55_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_55_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_55_m_axi_gmem_ARREGION;
	output wire qsort_55_m_axi_gmem_ARUSER;
	output wire qsort_55_m_axi_gmem_RREADY;
	input qsort_55_m_axi_gmem_RVALID;
	input qsort_55_m_axi_gmem_RID;
	input [63:0] qsort_55_m_axi_gmem_RDATA;
	input [1:0] qsort_55_m_axi_gmem_RRESP;
	input qsort_55_m_axi_gmem_RLAST;
	input qsort_55_m_axi_gmem_RUSER;
	input qsort_55_m_axi_gmem_AWREADY;
	output wire qsort_55_m_axi_gmem_AWVALID;
	output wire qsort_55_m_axi_gmem_AWID;
	output wire [63:0] qsort_55_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_55_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_55_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_55_m_axi_gmem_AWBURST;
	output wire qsort_55_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_55_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_55_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_55_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_55_m_axi_gmem_AWREGION;
	output wire qsort_55_m_axi_gmem_AWUSER;
	input qsort_55_m_axi_gmem_WREADY;
	output wire qsort_55_m_axi_gmem_WVALID;
	output wire [63:0] qsort_55_m_axi_gmem_WDATA;
	output wire [7:0] qsort_55_m_axi_gmem_WSTRB;
	output wire qsort_55_m_axi_gmem_WLAST;
	output wire qsort_55_m_axi_gmem_WUSER;
	output wire qsort_55_m_axi_gmem_BREADY;
	input qsort_55_m_axi_gmem_BVALID;
	input qsort_55_m_axi_gmem_BID;
	input [1:0] qsort_55_m_axi_gmem_BRESP;
	input qsort_55_m_axi_gmem_BUSER;
	output wire qsort_55_s_axi_control_ARREADY;
	input qsort_55_s_axi_control_ARVALID;
	input [5:0] qsort_55_s_axi_control_ARADDR;
	input qsort_55_s_axi_control_RREADY;
	output wire qsort_55_s_axi_control_RVALID;
	output wire [31:0] qsort_55_s_axi_control_RDATA;
	output wire [1:0] qsort_55_s_axi_control_RRESP;
	output wire qsort_55_s_axi_control_AWREADY;
	input qsort_55_s_axi_control_AWVALID;
	input [5:0] qsort_55_s_axi_control_AWADDR;
	output wire qsort_55_s_axi_control_WREADY;
	input qsort_55_s_axi_control_WVALID;
	input [31:0] qsort_55_s_axi_control_WDATA;
	input [3:0] qsort_55_s_axi_control_WSTRB;
	input qsort_55_s_axi_control_BREADY;
	output wire qsort_55_s_axi_control_BVALID;
	output wire [1:0] qsort_55_s_axi_control_BRESP;
	input qsort_56_m_axi_gmem_ARREADY;
	output wire qsort_56_m_axi_gmem_ARVALID;
	output wire qsort_56_m_axi_gmem_ARID;
	output wire [63:0] qsort_56_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_56_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_56_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_56_m_axi_gmem_ARBURST;
	output wire qsort_56_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_56_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_56_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_56_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_56_m_axi_gmem_ARREGION;
	output wire qsort_56_m_axi_gmem_ARUSER;
	output wire qsort_56_m_axi_gmem_RREADY;
	input qsort_56_m_axi_gmem_RVALID;
	input qsort_56_m_axi_gmem_RID;
	input [63:0] qsort_56_m_axi_gmem_RDATA;
	input [1:0] qsort_56_m_axi_gmem_RRESP;
	input qsort_56_m_axi_gmem_RLAST;
	input qsort_56_m_axi_gmem_RUSER;
	input qsort_56_m_axi_gmem_AWREADY;
	output wire qsort_56_m_axi_gmem_AWVALID;
	output wire qsort_56_m_axi_gmem_AWID;
	output wire [63:0] qsort_56_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_56_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_56_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_56_m_axi_gmem_AWBURST;
	output wire qsort_56_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_56_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_56_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_56_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_56_m_axi_gmem_AWREGION;
	output wire qsort_56_m_axi_gmem_AWUSER;
	input qsort_56_m_axi_gmem_WREADY;
	output wire qsort_56_m_axi_gmem_WVALID;
	output wire [63:0] qsort_56_m_axi_gmem_WDATA;
	output wire [7:0] qsort_56_m_axi_gmem_WSTRB;
	output wire qsort_56_m_axi_gmem_WLAST;
	output wire qsort_56_m_axi_gmem_WUSER;
	output wire qsort_56_m_axi_gmem_BREADY;
	input qsort_56_m_axi_gmem_BVALID;
	input qsort_56_m_axi_gmem_BID;
	input [1:0] qsort_56_m_axi_gmem_BRESP;
	input qsort_56_m_axi_gmem_BUSER;
	output wire qsort_56_s_axi_control_ARREADY;
	input qsort_56_s_axi_control_ARVALID;
	input [5:0] qsort_56_s_axi_control_ARADDR;
	input qsort_56_s_axi_control_RREADY;
	output wire qsort_56_s_axi_control_RVALID;
	output wire [31:0] qsort_56_s_axi_control_RDATA;
	output wire [1:0] qsort_56_s_axi_control_RRESP;
	output wire qsort_56_s_axi_control_AWREADY;
	input qsort_56_s_axi_control_AWVALID;
	input [5:0] qsort_56_s_axi_control_AWADDR;
	output wire qsort_56_s_axi_control_WREADY;
	input qsort_56_s_axi_control_WVALID;
	input [31:0] qsort_56_s_axi_control_WDATA;
	input [3:0] qsort_56_s_axi_control_WSTRB;
	input qsort_56_s_axi_control_BREADY;
	output wire qsort_56_s_axi_control_BVALID;
	output wire [1:0] qsort_56_s_axi_control_BRESP;
	input qsort_57_m_axi_gmem_ARREADY;
	output wire qsort_57_m_axi_gmem_ARVALID;
	output wire qsort_57_m_axi_gmem_ARID;
	output wire [63:0] qsort_57_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_57_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_57_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_57_m_axi_gmem_ARBURST;
	output wire qsort_57_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_57_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_57_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_57_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_57_m_axi_gmem_ARREGION;
	output wire qsort_57_m_axi_gmem_ARUSER;
	output wire qsort_57_m_axi_gmem_RREADY;
	input qsort_57_m_axi_gmem_RVALID;
	input qsort_57_m_axi_gmem_RID;
	input [63:0] qsort_57_m_axi_gmem_RDATA;
	input [1:0] qsort_57_m_axi_gmem_RRESP;
	input qsort_57_m_axi_gmem_RLAST;
	input qsort_57_m_axi_gmem_RUSER;
	input qsort_57_m_axi_gmem_AWREADY;
	output wire qsort_57_m_axi_gmem_AWVALID;
	output wire qsort_57_m_axi_gmem_AWID;
	output wire [63:0] qsort_57_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_57_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_57_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_57_m_axi_gmem_AWBURST;
	output wire qsort_57_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_57_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_57_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_57_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_57_m_axi_gmem_AWREGION;
	output wire qsort_57_m_axi_gmem_AWUSER;
	input qsort_57_m_axi_gmem_WREADY;
	output wire qsort_57_m_axi_gmem_WVALID;
	output wire [63:0] qsort_57_m_axi_gmem_WDATA;
	output wire [7:0] qsort_57_m_axi_gmem_WSTRB;
	output wire qsort_57_m_axi_gmem_WLAST;
	output wire qsort_57_m_axi_gmem_WUSER;
	output wire qsort_57_m_axi_gmem_BREADY;
	input qsort_57_m_axi_gmem_BVALID;
	input qsort_57_m_axi_gmem_BID;
	input [1:0] qsort_57_m_axi_gmem_BRESP;
	input qsort_57_m_axi_gmem_BUSER;
	output wire qsort_57_s_axi_control_ARREADY;
	input qsort_57_s_axi_control_ARVALID;
	input [5:0] qsort_57_s_axi_control_ARADDR;
	input qsort_57_s_axi_control_RREADY;
	output wire qsort_57_s_axi_control_RVALID;
	output wire [31:0] qsort_57_s_axi_control_RDATA;
	output wire [1:0] qsort_57_s_axi_control_RRESP;
	output wire qsort_57_s_axi_control_AWREADY;
	input qsort_57_s_axi_control_AWVALID;
	input [5:0] qsort_57_s_axi_control_AWADDR;
	output wire qsort_57_s_axi_control_WREADY;
	input qsort_57_s_axi_control_WVALID;
	input [31:0] qsort_57_s_axi_control_WDATA;
	input [3:0] qsort_57_s_axi_control_WSTRB;
	input qsort_57_s_axi_control_BREADY;
	output wire qsort_57_s_axi_control_BVALID;
	output wire [1:0] qsort_57_s_axi_control_BRESP;
	input qsort_58_m_axi_gmem_ARREADY;
	output wire qsort_58_m_axi_gmem_ARVALID;
	output wire qsort_58_m_axi_gmem_ARID;
	output wire [63:0] qsort_58_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_58_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_58_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_58_m_axi_gmem_ARBURST;
	output wire qsort_58_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_58_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_58_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_58_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_58_m_axi_gmem_ARREGION;
	output wire qsort_58_m_axi_gmem_ARUSER;
	output wire qsort_58_m_axi_gmem_RREADY;
	input qsort_58_m_axi_gmem_RVALID;
	input qsort_58_m_axi_gmem_RID;
	input [63:0] qsort_58_m_axi_gmem_RDATA;
	input [1:0] qsort_58_m_axi_gmem_RRESP;
	input qsort_58_m_axi_gmem_RLAST;
	input qsort_58_m_axi_gmem_RUSER;
	input qsort_58_m_axi_gmem_AWREADY;
	output wire qsort_58_m_axi_gmem_AWVALID;
	output wire qsort_58_m_axi_gmem_AWID;
	output wire [63:0] qsort_58_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_58_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_58_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_58_m_axi_gmem_AWBURST;
	output wire qsort_58_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_58_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_58_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_58_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_58_m_axi_gmem_AWREGION;
	output wire qsort_58_m_axi_gmem_AWUSER;
	input qsort_58_m_axi_gmem_WREADY;
	output wire qsort_58_m_axi_gmem_WVALID;
	output wire [63:0] qsort_58_m_axi_gmem_WDATA;
	output wire [7:0] qsort_58_m_axi_gmem_WSTRB;
	output wire qsort_58_m_axi_gmem_WLAST;
	output wire qsort_58_m_axi_gmem_WUSER;
	output wire qsort_58_m_axi_gmem_BREADY;
	input qsort_58_m_axi_gmem_BVALID;
	input qsort_58_m_axi_gmem_BID;
	input [1:0] qsort_58_m_axi_gmem_BRESP;
	input qsort_58_m_axi_gmem_BUSER;
	output wire qsort_58_s_axi_control_ARREADY;
	input qsort_58_s_axi_control_ARVALID;
	input [5:0] qsort_58_s_axi_control_ARADDR;
	input qsort_58_s_axi_control_RREADY;
	output wire qsort_58_s_axi_control_RVALID;
	output wire [31:0] qsort_58_s_axi_control_RDATA;
	output wire [1:0] qsort_58_s_axi_control_RRESP;
	output wire qsort_58_s_axi_control_AWREADY;
	input qsort_58_s_axi_control_AWVALID;
	input [5:0] qsort_58_s_axi_control_AWADDR;
	output wire qsort_58_s_axi_control_WREADY;
	input qsort_58_s_axi_control_WVALID;
	input [31:0] qsort_58_s_axi_control_WDATA;
	input [3:0] qsort_58_s_axi_control_WSTRB;
	input qsort_58_s_axi_control_BREADY;
	output wire qsort_58_s_axi_control_BVALID;
	output wire [1:0] qsort_58_s_axi_control_BRESP;
	input qsort_59_m_axi_gmem_ARREADY;
	output wire qsort_59_m_axi_gmem_ARVALID;
	output wire qsort_59_m_axi_gmem_ARID;
	output wire [63:0] qsort_59_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_59_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_59_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_59_m_axi_gmem_ARBURST;
	output wire qsort_59_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_59_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_59_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_59_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_59_m_axi_gmem_ARREGION;
	output wire qsort_59_m_axi_gmem_ARUSER;
	output wire qsort_59_m_axi_gmem_RREADY;
	input qsort_59_m_axi_gmem_RVALID;
	input qsort_59_m_axi_gmem_RID;
	input [63:0] qsort_59_m_axi_gmem_RDATA;
	input [1:0] qsort_59_m_axi_gmem_RRESP;
	input qsort_59_m_axi_gmem_RLAST;
	input qsort_59_m_axi_gmem_RUSER;
	input qsort_59_m_axi_gmem_AWREADY;
	output wire qsort_59_m_axi_gmem_AWVALID;
	output wire qsort_59_m_axi_gmem_AWID;
	output wire [63:0] qsort_59_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_59_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_59_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_59_m_axi_gmem_AWBURST;
	output wire qsort_59_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_59_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_59_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_59_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_59_m_axi_gmem_AWREGION;
	output wire qsort_59_m_axi_gmem_AWUSER;
	input qsort_59_m_axi_gmem_WREADY;
	output wire qsort_59_m_axi_gmem_WVALID;
	output wire [63:0] qsort_59_m_axi_gmem_WDATA;
	output wire [7:0] qsort_59_m_axi_gmem_WSTRB;
	output wire qsort_59_m_axi_gmem_WLAST;
	output wire qsort_59_m_axi_gmem_WUSER;
	output wire qsort_59_m_axi_gmem_BREADY;
	input qsort_59_m_axi_gmem_BVALID;
	input qsort_59_m_axi_gmem_BID;
	input [1:0] qsort_59_m_axi_gmem_BRESP;
	input qsort_59_m_axi_gmem_BUSER;
	output wire qsort_59_s_axi_control_ARREADY;
	input qsort_59_s_axi_control_ARVALID;
	input [5:0] qsort_59_s_axi_control_ARADDR;
	input qsort_59_s_axi_control_RREADY;
	output wire qsort_59_s_axi_control_RVALID;
	output wire [31:0] qsort_59_s_axi_control_RDATA;
	output wire [1:0] qsort_59_s_axi_control_RRESP;
	output wire qsort_59_s_axi_control_AWREADY;
	input qsort_59_s_axi_control_AWVALID;
	input [5:0] qsort_59_s_axi_control_AWADDR;
	output wire qsort_59_s_axi_control_WREADY;
	input qsort_59_s_axi_control_WVALID;
	input [31:0] qsort_59_s_axi_control_WDATA;
	input [3:0] qsort_59_s_axi_control_WSTRB;
	input qsort_59_s_axi_control_BREADY;
	output wire qsort_59_s_axi_control_BVALID;
	output wire [1:0] qsort_59_s_axi_control_BRESP;
	input qsort_60_m_axi_gmem_ARREADY;
	output wire qsort_60_m_axi_gmem_ARVALID;
	output wire qsort_60_m_axi_gmem_ARID;
	output wire [63:0] qsort_60_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_60_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_60_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_60_m_axi_gmem_ARBURST;
	output wire qsort_60_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_60_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_60_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_60_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_60_m_axi_gmem_ARREGION;
	output wire qsort_60_m_axi_gmem_ARUSER;
	output wire qsort_60_m_axi_gmem_RREADY;
	input qsort_60_m_axi_gmem_RVALID;
	input qsort_60_m_axi_gmem_RID;
	input [63:0] qsort_60_m_axi_gmem_RDATA;
	input [1:0] qsort_60_m_axi_gmem_RRESP;
	input qsort_60_m_axi_gmem_RLAST;
	input qsort_60_m_axi_gmem_RUSER;
	input qsort_60_m_axi_gmem_AWREADY;
	output wire qsort_60_m_axi_gmem_AWVALID;
	output wire qsort_60_m_axi_gmem_AWID;
	output wire [63:0] qsort_60_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_60_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_60_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_60_m_axi_gmem_AWBURST;
	output wire qsort_60_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_60_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_60_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_60_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_60_m_axi_gmem_AWREGION;
	output wire qsort_60_m_axi_gmem_AWUSER;
	input qsort_60_m_axi_gmem_WREADY;
	output wire qsort_60_m_axi_gmem_WVALID;
	output wire [63:0] qsort_60_m_axi_gmem_WDATA;
	output wire [7:0] qsort_60_m_axi_gmem_WSTRB;
	output wire qsort_60_m_axi_gmem_WLAST;
	output wire qsort_60_m_axi_gmem_WUSER;
	output wire qsort_60_m_axi_gmem_BREADY;
	input qsort_60_m_axi_gmem_BVALID;
	input qsort_60_m_axi_gmem_BID;
	input [1:0] qsort_60_m_axi_gmem_BRESP;
	input qsort_60_m_axi_gmem_BUSER;
	output wire qsort_60_s_axi_control_ARREADY;
	input qsort_60_s_axi_control_ARVALID;
	input [5:0] qsort_60_s_axi_control_ARADDR;
	input qsort_60_s_axi_control_RREADY;
	output wire qsort_60_s_axi_control_RVALID;
	output wire [31:0] qsort_60_s_axi_control_RDATA;
	output wire [1:0] qsort_60_s_axi_control_RRESP;
	output wire qsort_60_s_axi_control_AWREADY;
	input qsort_60_s_axi_control_AWVALID;
	input [5:0] qsort_60_s_axi_control_AWADDR;
	output wire qsort_60_s_axi_control_WREADY;
	input qsort_60_s_axi_control_WVALID;
	input [31:0] qsort_60_s_axi_control_WDATA;
	input [3:0] qsort_60_s_axi_control_WSTRB;
	input qsort_60_s_axi_control_BREADY;
	output wire qsort_60_s_axi_control_BVALID;
	output wire [1:0] qsort_60_s_axi_control_BRESP;
	input qsort_61_m_axi_gmem_ARREADY;
	output wire qsort_61_m_axi_gmem_ARVALID;
	output wire qsort_61_m_axi_gmem_ARID;
	output wire [63:0] qsort_61_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_61_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_61_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_61_m_axi_gmem_ARBURST;
	output wire qsort_61_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_61_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_61_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_61_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_61_m_axi_gmem_ARREGION;
	output wire qsort_61_m_axi_gmem_ARUSER;
	output wire qsort_61_m_axi_gmem_RREADY;
	input qsort_61_m_axi_gmem_RVALID;
	input qsort_61_m_axi_gmem_RID;
	input [63:0] qsort_61_m_axi_gmem_RDATA;
	input [1:0] qsort_61_m_axi_gmem_RRESP;
	input qsort_61_m_axi_gmem_RLAST;
	input qsort_61_m_axi_gmem_RUSER;
	input qsort_61_m_axi_gmem_AWREADY;
	output wire qsort_61_m_axi_gmem_AWVALID;
	output wire qsort_61_m_axi_gmem_AWID;
	output wire [63:0] qsort_61_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_61_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_61_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_61_m_axi_gmem_AWBURST;
	output wire qsort_61_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_61_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_61_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_61_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_61_m_axi_gmem_AWREGION;
	output wire qsort_61_m_axi_gmem_AWUSER;
	input qsort_61_m_axi_gmem_WREADY;
	output wire qsort_61_m_axi_gmem_WVALID;
	output wire [63:0] qsort_61_m_axi_gmem_WDATA;
	output wire [7:0] qsort_61_m_axi_gmem_WSTRB;
	output wire qsort_61_m_axi_gmem_WLAST;
	output wire qsort_61_m_axi_gmem_WUSER;
	output wire qsort_61_m_axi_gmem_BREADY;
	input qsort_61_m_axi_gmem_BVALID;
	input qsort_61_m_axi_gmem_BID;
	input [1:0] qsort_61_m_axi_gmem_BRESP;
	input qsort_61_m_axi_gmem_BUSER;
	output wire qsort_61_s_axi_control_ARREADY;
	input qsort_61_s_axi_control_ARVALID;
	input [5:0] qsort_61_s_axi_control_ARADDR;
	input qsort_61_s_axi_control_RREADY;
	output wire qsort_61_s_axi_control_RVALID;
	output wire [31:0] qsort_61_s_axi_control_RDATA;
	output wire [1:0] qsort_61_s_axi_control_RRESP;
	output wire qsort_61_s_axi_control_AWREADY;
	input qsort_61_s_axi_control_AWVALID;
	input [5:0] qsort_61_s_axi_control_AWADDR;
	output wire qsort_61_s_axi_control_WREADY;
	input qsort_61_s_axi_control_WVALID;
	input [31:0] qsort_61_s_axi_control_WDATA;
	input [3:0] qsort_61_s_axi_control_WSTRB;
	input qsort_61_s_axi_control_BREADY;
	output wire qsort_61_s_axi_control_BVALID;
	output wire [1:0] qsort_61_s_axi_control_BRESP;
	input qsort_62_m_axi_gmem_ARREADY;
	output wire qsort_62_m_axi_gmem_ARVALID;
	output wire qsort_62_m_axi_gmem_ARID;
	output wire [63:0] qsort_62_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_62_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_62_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_62_m_axi_gmem_ARBURST;
	output wire qsort_62_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_62_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_62_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_62_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_62_m_axi_gmem_ARREGION;
	output wire qsort_62_m_axi_gmem_ARUSER;
	output wire qsort_62_m_axi_gmem_RREADY;
	input qsort_62_m_axi_gmem_RVALID;
	input qsort_62_m_axi_gmem_RID;
	input [63:0] qsort_62_m_axi_gmem_RDATA;
	input [1:0] qsort_62_m_axi_gmem_RRESP;
	input qsort_62_m_axi_gmem_RLAST;
	input qsort_62_m_axi_gmem_RUSER;
	input qsort_62_m_axi_gmem_AWREADY;
	output wire qsort_62_m_axi_gmem_AWVALID;
	output wire qsort_62_m_axi_gmem_AWID;
	output wire [63:0] qsort_62_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_62_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_62_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_62_m_axi_gmem_AWBURST;
	output wire qsort_62_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_62_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_62_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_62_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_62_m_axi_gmem_AWREGION;
	output wire qsort_62_m_axi_gmem_AWUSER;
	input qsort_62_m_axi_gmem_WREADY;
	output wire qsort_62_m_axi_gmem_WVALID;
	output wire [63:0] qsort_62_m_axi_gmem_WDATA;
	output wire [7:0] qsort_62_m_axi_gmem_WSTRB;
	output wire qsort_62_m_axi_gmem_WLAST;
	output wire qsort_62_m_axi_gmem_WUSER;
	output wire qsort_62_m_axi_gmem_BREADY;
	input qsort_62_m_axi_gmem_BVALID;
	input qsort_62_m_axi_gmem_BID;
	input [1:0] qsort_62_m_axi_gmem_BRESP;
	input qsort_62_m_axi_gmem_BUSER;
	output wire qsort_62_s_axi_control_ARREADY;
	input qsort_62_s_axi_control_ARVALID;
	input [5:0] qsort_62_s_axi_control_ARADDR;
	input qsort_62_s_axi_control_RREADY;
	output wire qsort_62_s_axi_control_RVALID;
	output wire [31:0] qsort_62_s_axi_control_RDATA;
	output wire [1:0] qsort_62_s_axi_control_RRESP;
	output wire qsort_62_s_axi_control_AWREADY;
	input qsort_62_s_axi_control_AWVALID;
	input [5:0] qsort_62_s_axi_control_AWADDR;
	output wire qsort_62_s_axi_control_WREADY;
	input qsort_62_s_axi_control_WVALID;
	input [31:0] qsort_62_s_axi_control_WDATA;
	input [3:0] qsort_62_s_axi_control_WSTRB;
	input qsort_62_s_axi_control_BREADY;
	output wire qsort_62_s_axi_control_BVALID;
	output wire [1:0] qsort_62_s_axi_control_BRESP;
	input qsort_63_m_axi_gmem_ARREADY;
	output wire qsort_63_m_axi_gmem_ARVALID;
	output wire qsort_63_m_axi_gmem_ARID;
	output wire [63:0] qsort_63_m_axi_gmem_ARADDR;
	output wire [7:0] qsort_63_m_axi_gmem_ARLEN;
	output wire [2:0] qsort_63_m_axi_gmem_ARSIZE;
	output wire [1:0] qsort_63_m_axi_gmem_ARBURST;
	output wire qsort_63_m_axi_gmem_ARLOCK;
	output wire [3:0] qsort_63_m_axi_gmem_ARCACHE;
	output wire [2:0] qsort_63_m_axi_gmem_ARPROT;
	output wire [3:0] qsort_63_m_axi_gmem_ARQOS;
	output wire [3:0] qsort_63_m_axi_gmem_ARREGION;
	output wire qsort_63_m_axi_gmem_ARUSER;
	output wire qsort_63_m_axi_gmem_RREADY;
	input qsort_63_m_axi_gmem_RVALID;
	input qsort_63_m_axi_gmem_RID;
	input [63:0] qsort_63_m_axi_gmem_RDATA;
	input [1:0] qsort_63_m_axi_gmem_RRESP;
	input qsort_63_m_axi_gmem_RLAST;
	input qsort_63_m_axi_gmem_RUSER;
	input qsort_63_m_axi_gmem_AWREADY;
	output wire qsort_63_m_axi_gmem_AWVALID;
	output wire qsort_63_m_axi_gmem_AWID;
	output wire [63:0] qsort_63_m_axi_gmem_AWADDR;
	output wire [7:0] qsort_63_m_axi_gmem_AWLEN;
	output wire [2:0] qsort_63_m_axi_gmem_AWSIZE;
	output wire [1:0] qsort_63_m_axi_gmem_AWBURST;
	output wire qsort_63_m_axi_gmem_AWLOCK;
	output wire [3:0] qsort_63_m_axi_gmem_AWCACHE;
	output wire [2:0] qsort_63_m_axi_gmem_AWPROT;
	output wire [3:0] qsort_63_m_axi_gmem_AWQOS;
	output wire [3:0] qsort_63_m_axi_gmem_AWREGION;
	output wire qsort_63_m_axi_gmem_AWUSER;
	input qsort_63_m_axi_gmem_WREADY;
	output wire qsort_63_m_axi_gmem_WVALID;
	output wire [63:0] qsort_63_m_axi_gmem_WDATA;
	output wire [7:0] qsort_63_m_axi_gmem_WSTRB;
	output wire qsort_63_m_axi_gmem_WLAST;
	output wire qsort_63_m_axi_gmem_WUSER;
	output wire qsort_63_m_axi_gmem_BREADY;
	input qsort_63_m_axi_gmem_BVALID;
	input qsort_63_m_axi_gmem_BID;
	input [1:0] qsort_63_m_axi_gmem_BRESP;
	input qsort_63_m_axi_gmem_BUSER;
	output wire qsort_63_s_axi_control_ARREADY;
	input qsort_63_s_axi_control_ARVALID;
	input [5:0] qsort_63_s_axi_control_ARADDR;
	input qsort_63_s_axi_control_RREADY;
	output wire qsort_63_s_axi_control_RVALID;
	output wire [31:0] qsort_63_s_axi_control_RDATA;
	output wire [1:0] qsort_63_s_axi_control_RRESP;
	output wire qsort_63_s_axi_control_AWREADY;
	input qsort_63_s_axi_control_AWVALID;
	input [5:0] qsort_63_s_axi_control_AWADDR;
	output wire qsort_63_s_axi_control_WREADY;
	input qsort_63_s_axi_control_WVALID;
	input [31:0] qsort_63_s_axi_control_WDATA;
	input [3:0] qsort_63_s_axi_control_WSTRB;
	input qsort_63_s_axi_control_BREADY;
	output wire qsort_63_s_axi_control_BVALID;
	output wire [1:0] qsort_63_s_axi_control_BRESP;
	input qsort_schedulerAXI_0_ARREADY;
	output wire qsort_schedulerAXI_0_ARVALID;
	output wire qsort_schedulerAXI_0_ARID;
	output wire [63:0] qsort_schedulerAXI_0_ARADDR;
	output wire [7:0] qsort_schedulerAXI_0_ARLEN;
	output wire [2:0] qsort_schedulerAXI_0_ARSIZE;
	output wire [1:0] qsort_schedulerAXI_0_ARBURST;
	output wire qsort_schedulerAXI_0_ARLOCK;
	output wire [3:0] qsort_schedulerAXI_0_ARCACHE;
	output wire [2:0] qsort_schedulerAXI_0_ARPROT;
	output wire [3:0] qsort_schedulerAXI_0_ARQOS;
	output wire [3:0] qsort_schedulerAXI_0_ARREGION;
	output wire qsort_schedulerAXI_0_RREADY;
	input qsort_schedulerAXI_0_RVALID;
	input qsort_schedulerAXI_0_RID;
	input [255:0] qsort_schedulerAXI_0_RDATA;
	input [1:0] qsort_schedulerAXI_0_RRESP;
	input qsort_schedulerAXI_0_RLAST;
	input qsort_schedulerAXI_0_AWREADY;
	output wire qsort_schedulerAXI_0_AWVALID;
	output wire qsort_schedulerAXI_0_AWID;
	output wire [63:0] qsort_schedulerAXI_0_AWADDR;
	output wire [7:0] qsort_schedulerAXI_0_AWLEN;
	output wire [2:0] qsort_schedulerAXI_0_AWSIZE;
	output wire [1:0] qsort_schedulerAXI_0_AWBURST;
	output wire qsort_schedulerAXI_0_AWLOCK;
	output wire [3:0] qsort_schedulerAXI_0_AWCACHE;
	output wire [2:0] qsort_schedulerAXI_0_AWPROT;
	output wire [3:0] qsort_schedulerAXI_0_AWQOS;
	output wire [3:0] qsort_schedulerAXI_0_AWREGION;
	input qsort_schedulerAXI_0_WREADY;
	output wire qsort_schedulerAXI_0_WVALID;
	output wire [255:0] qsort_schedulerAXI_0_WDATA;
	output wire [31:0] qsort_schedulerAXI_0_WSTRB;
	output wire qsort_schedulerAXI_0_WLAST;
	output wire qsort_schedulerAXI_0_BREADY;
	input qsort_schedulerAXI_0_BVALID;
	input qsort_schedulerAXI_0_BID;
	input [1:0] qsort_schedulerAXI_0_BRESP;
	input sync_schedulerAXI_0_ARREADY;
	output wire sync_schedulerAXI_0_ARVALID;
	output wire sync_schedulerAXI_0_ARID;
	output wire [63:0] sync_schedulerAXI_0_ARADDR;
	output wire [7:0] sync_schedulerAXI_0_ARLEN;
	output wire [2:0] sync_schedulerAXI_0_ARSIZE;
	output wire [1:0] sync_schedulerAXI_0_ARBURST;
	output wire sync_schedulerAXI_0_ARLOCK;
	output wire [3:0] sync_schedulerAXI_0_ARCACHE;
	output wire [2:0] sync_schedulerAXI_0_ARPROT;
	output wire [3:0] sync_schedulerAXI_0_ARQOS;
	output wire [3:0] sync_schedulerAXI_0_ARREGION;
	output wire sync_schedulerAXI_0_RREADY;
	input sync_schedulerAXI_0_RVALID;
	input sync_schedulerAXI_0_RID;
	input [127:0] sync_schedulerAXI_0_RDATA;
	input [1:0] sync_schedulerAXI_0_RRESP;
	input sync_schedulerAXI_0_RLAST;
	input sync_schedulerAXI_0_AWREADY;
	output wire sync_schedulerAXI_0_AWVALID;
	output wire sync_schedulerAXI_0_AWID;
	output wire [63:0] sync_schedulerAXI_0_AWADDR;
	output wire [7:0] sync_schedulerAXI_0_AWLEN;
	output wire [2:0] sync_schedulerAXI_0_AWSIZE;
	output wire [1:0] sync_schedulerAXI_0_AWBURST;
	output wire sync_schedulerAXI_0_AWLOCK;
	output wire [3:0] sync_schedulerAXI_0_AWCACHE;
	output wire [2:0] sync_schedulerAXI_0_AWPROT;
	output wire [3:0] sync_schedulerAXI_0_AWQOS;
	output wire [3:0] sync_schedulerAXI_0_AWREGION;
	input sync_schedulerAXI_0_WREADY;
	output wire sync_schedulerAXI_0_WVALID;
	output wire [127:0] sync_schedulerAXI_0_WDATA;
	output wire [15:0] sync_schedulerAXI_0_WSTRB;
	output wire sync_schedulerAXI_0_WLAST;
	output wire sync_schedulerAXI_0_BREADY;
	input sync_schedulerAXI_0_BVALID;
	input sync_schedulerAXI_0_BID;
	input [1:0] sync_schedulerAXI_0_BRESP;
	input sync_closureAllocatorAXI_0_ARREADY;
	output wire sync_closureAllocatorAXI_0_ARVALID;
	output wire [4:0] sync_closureAllocatorAXI_0_ARID;
	output wire [63:0] sync_closureAllocatorAXI_0_ARADDR;
	output wire [7:0] sync_closureAllocatorAXI_0_ARLEN;
	output wire [2:0] sync_closureAllocatorAXI_0_ARSIZE;
	output wire [1:0] sync_closureAllocatorAXI_0_ARBURST;
	output wire sync_closureAllocatorAXI_0_ARLOCK;
	output wire [3:0] sync_closureAllocatorAXI_0_ARCACHE;
	output wire [2:0] sync_closureAllocatorAXI_0_ARPROT;
	output wire [3:0] sync_closureAllocatorAXI_0_ARQOS;
	output wire [3:0] sync_closureAllocatorAXI_0_ARREGION;
	output wire sync_closureAllocatorAXI_0_RREADY;
	input sync_closureAllocatorAXI_0_RVALID;
	input [4:0] sync_closureAllocatorAXI_0_RID;
	input [63:0] sync_closureAllocatorAXI_0_RDATA;
	input [1:0] sync_closureAllocatorAXI_0_RRESP;
	input sync_closureAllocatorAXI_0_RLAST;
	input sync_closureAllocatorAXI_0_AWREADY;
	output wire sync_closureAllocatorAXI_0_AWVALID;
	output wire [4:0] sync_closureAllocatorAXI_0_AWID;
	output wire [63:0] sync_closureAllocatorAXI_0_AWADDR;
	output wire [7:0] sync_closureAllocatorAXI_0_AWLEN;
	output wire [2:0] sync_closureAllocatorAXI_0_AWSIZE;
	output wire [1:0] sync_closureAllocatorAXI_0_AWBURST;
	output wire sync_closureAllocatorAXI_0_AWLOCK;
	output wire [3:0] sync_closureAllocatorAXI_0_AWCACHE;
	output wire [2:0] sync_closureAllocatorAXI_0_AWPROT;
	output wire [3:0] sync_closureAllocatorAXI_0_AWQOS;
	output wire [3:0] sync_closureAllocatorAXI_0_AWREGION;
	input sync_closureAllocatorAXI_0_WREADY;
	output wire sync_closureAllocatorAXI_0_WVALID;
	output wire [63:0] sync_closureAllocatorAXI_0_WDATA;
	output wire [7:0] sync_closureAllocatorAXI_0_WSTRB;
	output wire sync_closureAllocatorAXI_0_WLAST;
	output wire sync_closureAllocatorAXI_0_BREADY;
	input sync_closureAllocatorAXI_0_BVALID;
	input [4:0] sync_closureAllocatorAXI_0_BID;
	input [1:0] sync_closureAllocatorAXI_0_BRESP;
	input sync_closureAllocatorAXI_1_ARREADY;
	output wire sync_closureAllocatorAXI_1_ARVALID;
	output wire [4:0] sync_closureAllocatorAXI_1_ARID;
	output wire [63:0] sync_closureAllocatorAXI_1_ARADDR;
	output wire [7:0] sync_closureAllocatorAXI_1_ARLEN;
	output wire [2:0] sync_closureAllocatorAXI_1_ARSIZE;
	output wire [1:0] sync_closureAllocatorAXI_1_ARBURST;
	output wire sync_closureAllocatorAXI_1_ARLOCK;
	output wire [3:0] sync_closureAllocatorAXI_1_ARCACHE;
	output wire [2:0] sync_closureAllocatorAXI_1_ARPROT;
	output wire [3:0] sync_closureAllocatorAXI_1_ARQOS;
	output wire [3:0] sync_closureAllocatorAXI_1_ARREGION;
	output wire sync_closureAllocatorAXI_1_RREADY;
	input sync_closureAllocatorAXI_1_RVALID;
	input [4:0] sync_closureAllocatorAXI_1_RID;
	input [63:0] sync_closureAllocatorAXI_1_RDATA;
	input [1:0] sync_closureAllocatorAXI_1_RRESP;
	input sync_closureAllocatorAXI_1_RLAST;
	input sync_closureAllocatorAXI_1_AWREADY;
	output wire sync_closureAllocatorAXI_1_AWVALID;
	output wire [4:0] sync_closureAllocatorAXI_1_AWID;
	output wire [63:0] sync_closureAllocatorAXI_1_AWADDR;
	output wire [7:0] sync_closureAllocatorAXI_1_AWLEN;
	output wire [2:0] sync_closureAllocatorAXI_1_AWSIZE;
	output wire [1:0] sync_closureAllocatorAXI_1_AWBURST;
	output wire sync_closureAllocatorAXI_1_AWLOCK;
	output wire [3:0] sync_closureAllocatorAXI_1_AWCACHE;
	output wire [2:0] sync_closureAllocatorAXI_1_AWPROT;
	output wire [3:0] sync_closureAllocatorAXI_1_AWQOS;
	output wire [3:0] sync_closureAllocatorAXI_1_AWREGION;
	input sync_closureAllocatorAXI_1_WREADY;
	output wire sync_closureAllocatorAXI_1_WVALID;
	output wire [63:0] sync_closureAllocatorAXI_1_WDATA;
	output wire [7:0] sync_closureAllocatorAXI_1_WSTRB;
	output wire sync_closureAllocatorAXI_1_WLAST;
	output wire sync_closureAllocatorAXI_1_BREADY;
	input sync_closureAllocatorAXI_1_BVALID;
	input [4:0] sync_closureAllocatorAXI_1_BID;
	input [1:0] sync_closureAllocatorAXI_1_BRESP;
	input sync_closureAllocatorAXI_2_ARREADY;
	output wire sync_closureAllocatorAXI_2_ARVALID;
	output wire [4:0] sync_closureAllocatorAXI_2_ARID;
	output wire [63:0] sync_closureAllocatorAXI_2_ARADDR;
	output wire [7:0] sync_closureAllocatorAXI_2_ARLEN;
	output wire [2:0] sync_closureAllocatorAXI_2_ARSIZE;
	output wire [1:0] sync_closureAllocatorAXI_2_ARBURST;
	output wire sync_closureAllocatorAXI_2_ARLOCK;
	output wire [3:0] sync_closureAllocatorAXI_2_ARCACHE;
	output wire [2:0] sync_closureAllocatorAXI_2_ARPROT;
	output wire [3:0] sync_closureAllocatorAXI_2_ARQOS;
	output wire [3:0] sync_closureAllocatorAXI_2_ARREGION;
	output wire sync_closureAllocatorAXI_2_RREADY;
	input sync_closureAllocatorAXI_2_RVALID;
	input [4:0] sync_closureAllocatorAXI_2_RID;
	input [63:0] sync_closureAllocatorAXI_2_RDATA;
	input [1:0] sync_closureAllocatorAXI_2_RRESP;
	input sync_closureAllocatorAXI_2_RLAST;
	input sync_closureAllocatorAXI_2_AWREADY;
	output wire sync_closureAllocatorAXI_2_AWVALID;
	output wire [4:0] sync_closureAllocatorAXI_2_AWID;
	output wire [63:0] sync_closureAllocatorAXI_2_AWADDR;
	output wire [7:0] sync_closureAllocatorAXI_2_AWLEN;
	output wire [2:0] sync_closureAllocatorAXI_2_AWSIZE;
	output wire [1:0] sync_closureAllocatorAXI_2_AWBURST;
	output wire sync_closureAllocatorAXI_2_AWLOCK;
	output wire [3:0] sync_closureAllocatorAXI_2_AWCACHE;
	output wire [2:0] sync_closureAllocatorAXI_2_AWPROT;
	output wire [3:0] sync_closureAllocatorAXI_2_AWQOS;
	output wire [3:0] sync_closureAllocatorAXI_2_AWREGION;
	input sync_closureAllocatorAXI_2_WREADY;
	output wire sync_closureAllocatorAXI_2_WVALID;
	output wire [63:0] sync_closureAllocatorAXI_2_WDATA;
	output wire [7:0] sync_closureAllocatorAXI_2_WSTRB;
	output wire sync_closureAllocatorAXI_2_WLAST;
	output wire sync_closureAllocatorAXI_2_BREADY;
	input sync_closureAllocatorAXI_2_BVALID;
	input [4:0] sync_closureAllocatorAXI_2_BID;
	input [1:0] sync_closureAllocatorAXI_2_BRESP;
	input sync_closureAllocatorAXI_3_ARREADY;
	output wire sync_closureAllocatorAXI_3_ARVALID;
	output wire [4:0] sync_closureAllocatorAXI_3_ARID;
	output wire [63:0] sync_closureAllocatorAXI_3_ARADDR;
	output wire [7:0] sync_closureAllocatorAXI_3_ARLEN;
	output wire [2:0] sync_closureAllocatorAXI_3_ARSIZE;
	output wire [1:0] sync_closureAllocatorAXI_3_ARBURST;
	output wire sync_closureAllocatorAXI_3_ARLOCK;
	output wire [3:0] sync_closureAllocatorAXI_3_ARCACHE;
	output wire [2:0] sync_closureAllocatorAXI_3_ARPROT;
	output wire [3:0] sync_closureAllocatorAXI_3_ARQOS;
	output wire [3:0] sync_closureAllocatorAXI_3_ARREGION;
	output wire sync_closureAllocatorAXI_3_RREADY;
	input sync_closureAllocatorAXI_3_RVALID;
	input [4:0] sync_closureAllocatorAXI_3_RID;
	input [63:0] sync_closureAllocatorAXI_3_RDATA;
	input [1:0] sync_closureAllocatorAXI_3_RRESP;
	input sync_closureAllocatorAXI_3_RLAST;
	input sync_closureAllocatorAXI_3_AWREADY;
	output wire sync_closureAllocatorAXI_3_AWVALID;
	output wire [4:0] sync_closureAllocatorAXI_3_AWID;
	output wire [63:0] sync_closureAllocatorAXI_3_AWADDR;
	output wire [7:0] sync_closureAllocatorAXI_3_AWLEN;
	output wire [2:0] sync_closureAllocatorAXI_3_AWSIZE;
	output wire [1:0] sync_closureAllocatorAXI_3_AWBURST;
	output wire sync_closureAllocatorAXI_3_AWLOCK;
	output wire [3:0] sync_closureAllocatorAXI_3_AWCACHE;
	output wire [2:0] sync_closureAllocatorAXI_3_AWPROT;
	output wire [3:0] sync_closureAllocatorAXI_3_AWQOS;
	output wire [3:0] sync_closureAllocatorAXI_3_AWREGION;
	input sync_closureAllocatorAXI_3_WREADY;
	output wire sync_closureAllocatorAXI_3_WVALID;
	output wire [63:0] sync_closureAllocatorAXI_3_WDATA;
	output wire [7:0] sync_closureAllocatorAXI_3_WSTRB;
	output wire sync_closureAllocatorAXI_3_WLAST;
	output wire sync_closureAllocatorAXI_3_BREADY;
	input sync_closureAllocatorAXI_3_BVALID;
	input [4:0] sync_closureAllocatorAXI_3_BID;
	input [1:0] sync_closureAllocatorAXI_3_BRESP;
	input sync_argumentNotifierAXI_0_ARREADY;
	output wire sync_argumentNotifierAXI_0_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_0_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_0_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_0_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_0_ARBURST;
	output wire sync_argumentNotifierAXI_0_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_0_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_0_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_0_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_0_ARREGION;
	output wire sync_argumentNotifierAXI_0_RREADY;
	input sync_argumentNotifierAXI_0_RVALID;
	input [31:0] sync_argumentNotifierAXI_0_RDATA;
	input [1:0] sync_argumentNotifierAXI_0_RRESP;
	input sync_argumentNotifierAXI_0_RLAST;
	input sync_argumentNotifierAXI_0_AWREADY;
	output wire sync_argumentNotifierAXI_0_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_0_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_0_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_0_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_0_AWBURST;
	output wire sync_argumentNotifierAXI_0_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_0_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_0_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_0_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_0_AWREGION;
	input sync_argumentNotifierAXI_0_WREADY;
	output wire sync_argumentNotifierAXI_0_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_0_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_0_WSTRB;
	output wire sync_argumentNotifierAXI_0_WLAST;
	output wire sync_argumentNotifierAXI_0_BREADY;
	input sync_argumentNotifierAXI_0_BVALID;
	input [1:0] sync_argumentNotifierAXI_0_BRESP;
	input sync_argumentNotifierAXI_1_ARREADY;
	output wire sync_argumentNotifierAXI_1_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_1_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_1_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_1_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_1_ARBURST;
	output wire sync_argumentNotifierAXI_1_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_1_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_1_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_1_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_1_ARREGION;
	output wire sync_argumentNotifierAXI_1_RREADY;
	input sync_argumentNotifierAXI_1_RVALID;
	input [31:0] sync_argumentNotifierAXI_1_RDATA;
	input [1:0] sync_argumentNotifierAXI_1_RRESP;
	input sync_argumentNotifierAXI_1_RLAST;
	input sync_argumentNotifierAXI_1_AWREADY;
	output wire sync_argumentNotifierAXI_1_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_1_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_1_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_1_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_1_AWBURST;
	output wire sync_argumentNotifierAXI_1_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_1_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_1_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_1_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_1_AWREGION;
	input sync_argumentNotifierAXI_1_WREADY;
	output wire sync_argumentNotifierAXI_1_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_1_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_1_WSTRB;
	output wire sync_argumentNotifierAXI_1_WLAST;
	output wire sync_argumentNotifierAXI_1_BREADY;
	input sync_argumentNotifierAXI_1_BVALID;
	input [1:0] sync_argumentNotifierAXI_1_BRESP;
	input sync_argumentNotifierAXI_2_ARREADY;
	output wire sync_argumentNotifierAXI_2_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_2_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_2_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_2_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_2_ARBURST;
	output wire sync_argumentNotifierAXI_2_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_2_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_2_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_2_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_2_ARREGION;
	output wire sync_argumentNotifierAXI_2_RREADY;
	input sync_argumentNotifierAXI_2_RVALID;
	input [31:0] sync_argumentNotifierAXI_2_RDATA;
	input [1:0] sync_argumentNotifierAXI_2_RRESP;
	input sync_argumentNotifierAXI_2_RLAST;
	input sync_argumentNotifierAXI_2_AWREADY;
	output wire sync_argumentNotifierAXI_2_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_2_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_2_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_2_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_2_AWBURST;
	output wire sync_argumentNotifierAXI_2_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_2_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_2_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_2_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_2_AWREGION;
	input sync_argumentNotifierAXI_2_WREADY;
	output wire sync_argumentNotifierAXI_2_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_2_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_2_WSTRB;
	output wire sync_argumentNotifierAXI_2_WLAST;
	output wire sync_argumentNotifierAXI_2_BREADY;
	input sync_argumentNotifierAXI_2_BVALID;
	input [1:0] sync_argumentNotifierAXI_2_BRESP;
	input sync_argumentNotifierAXI_3_ARREADY;
	output wire sync_argumentNotifierAXI_3_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_3_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_3_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_3_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_3_ARBURST;
	output wire sync_argumentNotifierAXI_3_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_3_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_3_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_3_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_3_ARREGION;
	output wire sync_argumentNotifierAXI_3_RREADY;
	input sync_argumentNotifierAXI_3_RVALID;
	input [31:0] sync_argumentNotifierAXI_3_RDATA;
	input [1:0] sync_argumentNotifierAXI_3_RRESP;
	input sync_argumentNotifierAXI_3_RLAST;
	input sync_argumentNotifierAXI_3_AWREADY;
	output wire sync_argumentNotifierAXI_3_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_3_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_3_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_3_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_3_AWBURST;
	output wire sync_argumentNotifierAXI_3_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_3_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_3_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_3_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_3_AWREGION;
	input sync_argumentNotifierAXI_3_WREADY;
	output wire sync_argumentNotifierAXI_3_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_3_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_3_WSTRB;
	output wire sync_argumentNotifierAXI_3_WLAST;
	output wire sync_argumentNotifierAXI_3_BREADY;
	input sync_argumentNotifierAXI_3_BVALID;
	input [1:0] sync_argumentNotifierAXI_3_BRESP;
	input sync_argumentNotifierAXI_4_ARREADY;
	output wire sync_argumentNotifierAXI_4_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_4_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_4_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_4_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_4_ARBURST;
	output wire sync_argumentNotifierAXI_4_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_4_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_4_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_4_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_4_ARREGION;
	output wire sync_argumentNotifierAXI_4_RREADY;
	input sync_argumentNotifierAXI_4_RVALID;
	input [31:0] sync_argumentNotifierAXI_4_RDATA;
	input [1:0] sync_argumentNotifierAXI_4_RRESP;
	input sync_argumentNotifierAXI_4_RLAST;
	input sync_argumentNotifierAXI_4_AWREADY;
	output wire sync_argumentNotifierAXI_4_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_4_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_4_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_4_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_4_AWBURST;
	output wire sync_argumentNotifierAXI_4_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_4_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_4_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_4_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_4_AWREGION;
	input sync_argumentNotifierAXI_4_WREADY;
	output wire sync_argumentNotifierAXI_4_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_4_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_4_WSTRB;
	output wire sync_argumentNotifierAXI_4_WLAST;
	output wire sync_argumentNotifierAXI_4_BREADY;
	input sync_argumentNotifierAXI_4_BVALID;
	input [1:0] sync_argumentNotifierAXI_4_BRESP;
	input sync_argumentNotifierAXI_5_ARREADY;
	output wire sync_argumentNotifierAXI_5_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_5_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_5_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_5_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_5_ARBURST;
	output wire sync_argumentNotifierAXI_5_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_5_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_5_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_5_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_5_ARREGION;
	output wire sync_argumentNotifierAXI_5_RREADY;
	input sync_argumentNotifierAXI_5_RVALID;
	input [31:0] sync_argumentNotifierAXI_5_RDATA;
	input [1:0] sync_argumentNotifierAXI_5_RRESP;
	input sync_argumentNotifierAXI_5_RLAST;
	input sync_argumentNotifierAXI_5_AWREADY;
	output wire sync_argumentNotifierAXI_5_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_5_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_5_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_5_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_5_AWBURST;
	output wire sync_argumentNotifierAXI_5_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_5_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_5_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_5_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_5_AWREGION;
	input sync_argumentNotifierAXI_5_WREADY;
	output wire sync_argumentNotifierAXI_5_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_5_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_5_WSTRB;
	output wire sync_argumentNotifierAXI_5_WLAST;
	output wire sync_argumentNotifierAXI_5_BREADY;
	input sync_argumentNotifierAXI_5_BVALID;
	input [1:0] sync_argumentNotifierAXI_5_BRESP;
	input sync_argumentNotifierAXI_6_ARREADY;
	output wire sync_argumentNotifierAXI_6_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_6_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_6_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_6_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_6_ARBURST;
	output wire sync_argumentNotifierAXI_6_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_6_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_6_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_6_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_6_ARREGION;
	output wire sync_argumentNotifierAXI_6_RREADY;
	input sync_argumentNotifierAXI_6_RVALID;
	input [31:0] sync_argumentNotifierAXI_6_RDATA;
	input [1:0] sync_argumentNotifierAXI_6_RRESP;
	input sync_argumentNotifierAXI_6_RLAST;
	input sync_argumentNotifierAXI_6_AWREADY;
	output wire sync_argumentNotifierAXI_6_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_6_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_6_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_6_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_6_AWBURST;
	output wire sync_argumentNotifierAXI_6_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_6_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_6_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_6_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_6_AWREGION;
	input sync_argumentNotifierAXI_6_WREADY;
	output wire sync_argumentNotifierAXI_6_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_6_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_6_WSTRB;
	output wire sync_argumentNotifierAXI_6_WLAST;
	output wire sync_argumentNotifierAXI_6_BREADY;
	input sync_argumentNotifierAXI_6_BVALID;
	input [1:0] sync_argumentNotifierAXI_6_BRESP;
	input sync_argumentNotifierAXI_7_ARREADY;
	output wire sync_argumentNotifierAXI_7_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_7_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_7_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_7_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_7_ARBURST;
	output wire sync_argumentNotifierAXI_7_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_7_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_7_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_7_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_7_ARREGION;
	output wire sync_argumentNotifierAXI_7_RREADY;
	input sync_argumentNotifierAXI_7_RVALID;
	input [31:0] sync_argumentNotifierAXI_7_RDATA;
	input [1:0] sync_argumentNotifierAXI_7_RRESP;
	input sync_argumentNotifierAXI_7_RLAST;
	input sync_argumentNotifierAXI_7_AWREADY;
	output wire sync_argumentNotifierAXI_7_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_7_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_7_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_7_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_7_AWBURST;
	output wire sync_argumentNotifierAXI_7_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_7_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_7_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_7_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_7_AWREGION;
	input sync_argumentNotifierAXI_7_WREADY;
	output wire sync_argumentNotifierAXI_7_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_7_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_7_WSTRB;
	output wire sync_argumentNotifierAXI_7_WLAST;
	output wire sync_argumentNotifierAXI_7_BREADY;
	input sync_argumentNotifierAXI_7_BVALID;
	input [1:0] sync_argumentNotifierAXI_7_BRESP;
	input sync_argumentNotifierAXI_8_ARREADY;
	output wire sync_argumentNotifierAXI_8_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_8_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_8_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_8_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_8_ARBURST;
	output wire sync_argumentNotifierAXI_8_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_8_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_8_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_8_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_8_ARREGION;
	output wire sync_argumentNotifierAXI_8_RREADY;
	input sync_argumentNotifierAXI_8_RVALID;
	input [31:0] sync_argumentNotifierAXI_8_RDATA;
	input [1:0] sync_argumentNotifierAXI_8_RRESP;
	input sync_argumentNotifierAXI_8_RLAST;
	input sync_argumentNotifierAXI_8_AWREADY;
	output wire sync_argumentNotifierAXI_8_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_8_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_8_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_8_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_8_AWBURST;
	output wire sync_argumentNotifierAXI_8_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_8_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_8_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_8_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_8_AWREGION;
	input sync_argumentNotifierAXI_8_WREADY;
	output wire sync_argumentNotifierAXI_8_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_8_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_8_WSTRB;
	output wire sync_argumentNotifierAXI_8_WLAST;
	output wire sync_argumentNotifierAXI_8_BREADY;
	input sync_argumentNotifierAXI_8_BVALID;
	input [1:0] sync_argumentNotifierAXI_8_BRESP;
	input sync_argumentNotifierAXI_9_ARREADY;
	output wire sync_argumentNotifierAXI_9_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_9_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_9_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_9_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_9_ARBURST;
	output wire sync_argumentNotifierAXI_9_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_9_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_9_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_9_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_9_ARREGION;
	output wire sync_argumentNotifierAXI_9_RREADY;
	input sync_argumentNotifierAXI_9_RVALID;
	input [31:0] sync_argumentNotifierAXI_9_RDATA;
	input [1:0] sync_argumentNotifierAXI_9_RRESP;
	input sync_argumentNotifierAXI_9_RLAST;
	input sync_argumentNotifierAXI_9_AWREADY;
	output wire sync_argumentNotifierAXI_9_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_9_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_9_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_9_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_9_AWBURST;
	output wire sync_argumentNotifierAXI_9_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_9_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_9_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_9_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_9_AWREGION;
	input sync_argumentNotifierAXI_9_WREADY;
	output wire sync_argumentNotifierAXI_9_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_9_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_9_WSTRB;
	output wire sync_argumentNotifierAXI_9_WLAST;
	output wire sync_argumentNotifierAXI_9_BREADY;
	input sync_argumentNotifierAXI_9_BVALID;
	input [1:0] sync_argumentNotifierAXI_9_BRESP;
	input sync_argumentNotifierAXI_10_ARREADY;
	output wire sync_argumentNotifierAXI_10_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_10_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_10_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_10_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_10_ARBURST;
	output wire sync_argumentNotifierAXI_10_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_10_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_10_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_10_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_10_ARREGION;
	output wire sync_argumentNotifierAXI_10_RREADY;
	input sync_argumentNotifierAXI_10_RVALID;
	input [31:0] sync_argumentNotifierAXI_10_RDATA;
	input [1:0] sync_argumentNotifierAXI_10_RRESP;
	input sync_argumentNotifierAXI_10_RLAST;
	input sync_argumentNotifierAXI_10_AWREADY;
	output wire sync_argumentNotifierAXI_10_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_10_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_10_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_10_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_10_AWBURST;
	output wire sync_argumentNotifierAXI_10_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_10_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_10_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_10_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_10_AWREGION;
	input sync_argumentNotifierAXI_10_WREADY;
	output wire sync_argumentNotifierAXI_10_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_10_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_10_WSTRB;
	output wire sync_argumentNotifierAXI_10_WLAST;
	output wire sync_argumentNotifierAXI_10_BREADY;
	input sync_argumentNotifierAXI_10_BVALID;
	input [1:0] sync_argumentNotifierAXI_10_BRESP;
	input sync_argumentNotifierAXI_11_ARREADY;
	output wire sync_argumentNotifierAXI_11_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_11_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_11_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_11_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_11_ARBURST;
	output wire sync_argumentNotifierAXI_11_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_11_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_11_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_11_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_11_ARREGION;
	output wire sync_argumentNotifierAXI_11_RREADY;
	input sync_argumentNotifierAXI_11_RVALID;
	input [31:0] sync_argumentNotifierAXI_11_RDATA;
	input [1:0] sync_argumentNotifierAXI_11_RRESP;
	input sync_argumentNotifierAXI_11_RLAST;
	input sync_argumentNotifierAXI_11_AWREADY;
	output wire sync_argumentNotifierAXI_11_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_11_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_11_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_11_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_11_AWBURST;
	output wire sync_argumentNotifierAXI_11_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_11_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_11_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_11_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_11_AWREGION;
	input sync_argumentNotifierAXI_11_WREADY;
	output wire sync_argumentNotifierAXI_11_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_11_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_11_WSTRB;
	output wire sync_argumentNotifierAXI_11_WLAST;
	output wire sync_argumentNotifierAXI_11_BREADY;
	input sync_argumentNotifierAXI_11_BVALID;
	input [1:0] sync_argumentNotifierAXI_11_BRESP;
	input sync_argumentNotifierAXI_12_ARREADY;
	output wire sync_argumentNotifierAXI_12_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_12_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_12_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_12_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_12_ARBURST;
	output wire sync_argumentNotifierAXI_12_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_12_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_12_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_12_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_12_ARREGION;
	output wire sync_argumentNotifierAXI_12_RREADY;
	input sync_argumentNotifierAXI_12_RVALID;
	input [31:0] sync_argumentNotifierAXI_12_RDATA;
	input [1:0] sync_argumentNotifierAXI_12_RRESP;
	input sync_argumentNotifierAXI_12_RLAST;
	input sync_argumentNotifierAXI_12_AWREADY;
	output wire sync_argumentNotifierAXI_12_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_12_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_12_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_12_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_12_AWBURST;
	output wire sync_argumentNotifierAXI_12_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_12_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_12_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_12_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_12_AWREGION;
	input sync_argumentNotifierAXI_12_WREADY;
	output wire sync_argumentNotifierAXI_12_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_12_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_12_WSTRB;
	output wire sync_argumentNotifierAXI_12_WLAST;
	output wire sync_argumentNotifierAXI_12_BREADY;
	input sync_argumentNotifierAXI_12_BVALID;
	input [1:0] sync_argumentNotifierAXI_12_BRESP;
	input sync_argumentNotifierAXI_13_ARREADY;
	output wire sync_argumentNotifierAXI_13_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_13_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_13_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_13_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_13_ARBURST;
	output wire sync_argumentNotifierAXI_13_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_13_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_13_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_13_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_13_ARREGION;
	output wire sync_argumentNotifierAXI_13_RREADY;
	input sync_argumentNotifierAXI_13_RVALID;
	input [31:0] sync_argumentNotifierAXI_13_RDATA;
	input [1:0] sync_argumentNotifierAXI_13_RRESP;
	input sync_argumentNotifierAXI_13_RLAST;
	input sync_argumentNotifierAXI_13_AWREADY;
	output wire sync_argumentNotifierAXI_13_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_13_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_13_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_13_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_13_AWBURST;
	output wire sync_argumentNotifierAXI_13_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_13_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_13_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_13_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_13_AWREGION;
	input sync_argumentNotifierAXI_13_WREADY;
	output wire sync_argumentNotifierAXI_13_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_13_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_13_WSTRB;
	output wire sync_argumentNotifierAXI_13_WLAST;
	output wire sync_argumentNotifierAXI_13_BREADY;
	input sync_argumentNotifierAXI_13_BVALID;
	input [1:0] sync_argumentNotifierAXI_13_BRESP;
	input sync_argumentNotifierAXI_14_ARREADY;
	output wire sync_argumentNotifierAXI_14_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_14_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_14_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_14_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_14_ARBURST;
	output wire sync_argumentNotifierAXI_14_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_14_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_14_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_14_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_14_ARREGION;
	output wire sync_argumentNotifierAXI_14_RREADY;
	input sync_argumentNotifierAXI_14_RVALID;
	input [31:0] sync_argumentNotifierAXI_14_RDATA;
	input [1:0] sync_argumentNotifierAXI_14_RRESP;
	input sync_argumentNotifierAXI_14_RLAST;
	input sync_argumentNotifierAXI_14_AWREADY;
	output wire sync_argumentNotifierAXI_14_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_14_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_14_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_14_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_14_AWBURST;
	output wire sync_argumentNotifierAXI_14_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_14_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_14_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_14_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_14_AWREGION;
	input sync_argumentNotifierAXI_14_WREADY;
	output wire sync_argumentNotifierAXI_14_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_14_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_14_WSTRB;
	output wire sync_argumentNotifierAXI_14_WLAST;
	output wire sync_argumentNotifierAXI_14_BREADY;
	input sync_argumentNotifierAXI_14_BVALID;
	input [1:0] sync_argumentNotifierAXI_14_BRESP;
	input sync_argumentNotifierAXI_15_ARREADY;
	output wire sync_argumentNotifierAXI_15_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_15_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_15_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_15_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_15_ARBURST;
	output wire sync_argumentNotifierAXI_15_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_15_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_15_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_15_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_15_ARREGION;
	output wire sync_argumentNotifierAXI_15_RREADY;
	input sync_argumentNotifierAXI_15_RVALID;
	input [31:0] sync_argumentNotifierAXI_15_RDATA;
	input [1:0] sync_argumentNotifierAXI_15_RRESP;
	input sync_argumentNotifierAXI_15_RLAST;
	input sync_argumentNotifierAXI_15_AWREADY;
	output wire sync_argumentNotifierAXI_15_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_15_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_15_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_15_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_15_AWBURST;
	output wire sync_argumentNotifierAXI_15_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_15_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_15_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_15_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_15_AWREGION;
	input sync_argumentNotifierAXI_15_WREADY;
	output wire sync_argumentNotifierAXI_15_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_15_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_15_WSTRB;
	output wire sync_argumentNotifierAXI_15_WLAST;
	output wire sync_argumentNotifierAXI_15_BREADY;
	input sync_argumentNotifierAXI_15_BVALID;
	input [1:0] sync_argumentNotifierAXI_15_BRESP;
	input sync_argumentNotifierAXI_16_ARREADY;
	output wire sync_argumentNotifierAXI_16_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_16_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_16_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_16_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_16_ARBURST;
	output wire sync_argumentNotifierAXI_16_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_16_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_16_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_16_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_16_ARREGION;
	output wire sync_argumentNotifierAXI_16_RREADY;
	input sync_argumentNotifierAXI_16_RVALID;
	input [31:0] sync_argumentNotifierAXI_16_RDATA;
	input [1:0] sync_argumentNotifierAXI_16_RRESP;
	input sync_argumentNotifierAXI_16_RLAST;
	input sync_argumentNotifierAXI_16_AWREADY;
	output wire sync_argumentNotifierAXI_16_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_16_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_16_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_16_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_16_AWBURST;
	output wire sync_argumentNotifierAXI_16_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_16_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_16_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_16_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_16_AWREGION;
	input sync_argumentNotifierAXI_16_WREADY;
	output wire sync_argumentNotifierAXI_16_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_16_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_16_WSTRB;
	output wire sync_argumentNotifierAXI_16_WLAST;
	output wire sync_argumentNotifierAXI_16_BREADY;
	input sync_argumentNotifierAXI_16_BVALID;
	input [1:0] sync_argumentNotifierAXI_16_BRESP;
	input sync_argumentNotifierAXI_17_ARREADY;
	output wire sync_argumentNotifierAXI_17_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_17_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_17_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_17_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_17_ARBURST;
	output wire sync_argumentNotifierAXI_17_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_17_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_17_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_17_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_17_ARREGION;
	output wire sync_argumentNotifierAXI_17_RREADY;
	input sync_argumentNotifierAXI_17_RVALID;
	input [31:0] sync_argumentNotifierAXI_17_RDATA;
	input [1:0] sync_argumentNotifierAXI_17_RRESP;
	input sync_argumentNotifierAXI_17_RLAST;
	input sync_argumentNotifierAXI_17_AWREADY;
	output wire sync_argumentNotifierAXI_17_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_17_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_17_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_17_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_17_AWBURST;
	output wire sync_argumentNotifierAXI_17_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_17_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_17_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_17_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_17_AWREGION;
	input sync_argumentNotifierAXI_17_WREADY;
	output wire sync_argumentNotifierAXI_17_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_17_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_17_WSTRB;
	output wire sync_argumentNotifierAXI_17_WLAST;
	output wire sync_argumentNotifierAXI_17_BREADY;
	input sync_argumentNotifierAXI_17_BVALID;
	input [1:0] sync_argumentNotifierAXI_17_BRESP;
	input sync_argumentNotifierAXI_18_ARREADY;
	output wire sync_argumentNotifierAXI_18_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_18_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_18_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_18_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_18_ARBURST;
	output wire sync_argumentNotifierAXI_18_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_18_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_18_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_18_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_18_ARREGION;
	output wire sync_argumentNotifierAXI_18_RREADY;
	input sync_argumentNotifierAXI_18_RVALID;
	input [31:0] sync_argumentNotifierAXI_18_RDATA;
	input [1:0] sync_argumentNotifierAXI_18_RRESP;
	input sync_argumentNotifierAXI_18_RLAST;
	input sync_argumentNotifierAXI_18_AWREADY;
	output wire sync_argumentNotifierAXI_18_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_18_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_18_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_18_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_18_AWBURST;
	output wire sync_argumentNotifierAXI_18_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_18_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_18_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_18_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_18_AWREGION;
	input sync_argumentNotifierAXI_18_WREADY;
	output wire sync_argumentNotifierAXI_18_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_18_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_18_WSTRB;
	output wire sync_argumentNotifierAXI_18_WLAST;
	output wire sync_argumentNotifierAXI_18_BREADY;
	input sync_argumentNotifierAXI_18_BVALID;
	input [1:0] sync_argumentNotifierAXI_18_BRESP;
	input sync_argumentNotifierAXI_19_ARREADY;
	output wire sync_argumentNotifierAXI_19_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_19_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_19_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_19_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_19_ARBURST;
	output wire sync_argumentNotifierAXI_19_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_19_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_19_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_19_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_19_ARREGION;
	output wire sync_argumentNotifierAXI_19_RREADY;
	input sync_argumentNotifierAXI_19_RVALID;
	input [31:0] sync_argumentNotifierAXI_19_RDATA;
	input [1:0] sync_argumentNotifierAXI_19_RRESP;
	input sync_argumentNotifierAXI_19_RLAST;
	input sync_argumentNotifierAXI_19_AWREADY;
	output wire sync_argumentNotifierAXI_19_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_19_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_19_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_19_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_19_AWBURST;
	output wire sync_argumentNotifierAXI_19_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_19_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_19_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_19_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_19_AWREGION;
	input sync_argumentNotifierAXI_19_WREADY;
	output wire sync_argumentNotifierAXI_19_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_19_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_19_WSTRB;
	output wire sync_argumentNotifierAXI_19_WLAST;
	output wire sync_argumentNotifierAXI_19_BREADY;
	input sync_argumentNotifierAXI_19_BVALID;
	input [1:0] sync_argumentNotifierAXI_19_BRESP;
	input sync_argumentNotifierAXI_20_ARREADY;
	output wire sync_argumentNotifierAXI_20_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_20_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_20_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_20_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_20_ARBURST;
	output wire sync_argumentNotifierAXI_20_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_20_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_20_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_20_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_20_ARREGION;
	output wire sync_argumentNotifierAXI_20_RREADY;
	input sync_argumentNotifierAXI_20_RVALID;
	input [31:0] sync_argumentNotifierAXI_20_RDATA;
	input [1:0] sync_argumentNotifierAXI_20_RRESP;
	input sync_argumentNotifierAXI_20_RLAST;
	input sync_argumentNotifierAXI_20_AWREADY;
	output wire sync_argumentNotifierAXI_20_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_20_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_20_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_20_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_20_AWBURST;
	output wire sync_argumentNotifierAXI_20_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_20_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_20_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_20_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_20_AWREGION;
	input sync_argumentNotifierAXI_20_WREADY;
	output wire sync_argumentNotifierAXI_20_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_20_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_20_WSTRB;
	output wire sync_argumentNotifierAXI_20_WLAST;
	output wire sync_argumentNotifierAXI_20_BREADY;
	input sync_argumentNotifierAXI_20_BVALID;
	input [1:0] sync_argumentNotifierAXI_20_BRESP;
	input sync_argumentNotifierAXI_21_ARREADY;
	output wire sync_argumentNotifierAXI_21_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_21_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_21_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_21_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_21_ARBURST;
	output wire sync_argumentNotifierAXI_21_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_21_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_21_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_21_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_21_ARREGION;
	output wire sync_argumentNotifierAXI_21_RREADY;
	input sync_argumentNotifierAXI_21_RVALID;
	input [31:0] sync_argumentNotifierAXI_21_RDATA;
	input [1:0] sync_argumentNotifierAXI_21_RRESP;
	input sync_argumentNotifierAXI_21_RLAST;
	input sync_argumentNotifierAXI_21_AWREADY;
	output wire sync_argumentNotifierAXI_21_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_21_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_21_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_21_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_21_AWBURST;
	output wire sync_argumentNotifierAXI_21_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_21_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_21_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_21_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_21_AWREGION;
	input sync_argumentNotifierAXI_21_WREADY;
	output wire sync_argumentNotifierAXI_21_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_21_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_21_WSTRB;
	output wire sync_argumentNotifierAXI_21_WLAST;
	output wire sync_argumentNotifierAXI_21_BREADY;
	input sync_argumentNotifierAXI_21_BVALID;
	input [1:0] sync_argumentNotifierAXI_21_BRESP;
	input sync_argumentNotifierAXI_22_ARREADY;
	output wire sync_argumentNotifierAXI_22_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_22_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_22_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_22_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_22_ARBURST;
	output wire sync_argumentNotifierAXI_22_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_22_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_22_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_22_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_22_ARREGION;
	output wire sync_argumentNotifierAXI_22_RREADY;
	input sync_argumentNotifierAXI_22_RVALID;
	input [31:0] sync_argumentNotifierAXI_22_RDATA;
	input [1:0] sync_argumentNotifierAXI_22_RRESP;
	input sync_argumentNotifierAXI_22_RLAST;
	input sync_argumentNotifierAXI_22_AWREADY;
	output wire sync_argumentNotifierAXI_22_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_22_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_22_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_22_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_22_AWBURST;
	output wire sync_argumentNotifierAXI_22_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_22_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_22_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_22_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_22_AWREGION;
	input sync_argumentNotifierAXI_22_WREADY;
	output wire sync_argumentNotifierAXI_22_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_22_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_22_WSTRB;
	output wire sync_argumentNotifierAXI_22_WLAST;
	output wire sync_argumentNotifierAXI_22_BREADY;
	input sync_argumentNotifierAXI_22_BVALID;
	input [1:0] sync_argumentNotifierAXI_22_BRESP;
	input sync_argumentNotifierAXI_23_ARREADY;
	output wire sync_argumentNotifierAXI_23_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_23_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_23_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_23_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_23_ARBURST;
	output wire sync_argumentNotifierAXI_23_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_23_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_23_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_23_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_23_ARREGION;
	output wire sync_argumentNotifierAXI_23_RREADY;
	input sync_argumentNotifierAXI_23_RVALID;
	input [31:0] sync_argumentNotifierAXI_23_RDATA;
	input [1:0] sync_argumentNotifierAXI_23_RRESP;
	input sync_argumentNotifierAXI_23_RLAST;
	input sync_argumentNotifierAXI_23_AWREADY;
	output wire sync_argumentNotifierAXI_23_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_23_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_23_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_23_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_23_AWBURST;
	output wire sync_argumentNotifierAXI_23_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_23_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_23_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_23_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_23_AWREGION;
	input sync_argumentNotifierAXI_23_WREADY;
	output wire sync_argumentNotifierAXI_23_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_23_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_23_WSTRB;
	output wire sync_argumentNotifierAXI_23_WLAST;
	output wire sync_argumentNotifierAXI_23_BREADY;
	input sync_argumentNotifierAXI_23_BVALID;
	input [1:0] sync_argumentNotifierAXI_23_BRESP;
	input sync_argumentNotifierAXI_24_ARREADY;
	output wire sync_argumentNotifierAXI_24_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_24_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_24_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_24_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_24_ARBURST;
	output wire sync_argumentNotifierAXI_24_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_24_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_24_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_24_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_24_ARREGION;
	output wire sync_argumentNotifierAXI_24_RREADY;
	input sync_argumentNotifierAXI_24_RVALID;
	input [31:0] sync_argumentNotifierAXI_24_RDATA;
	input [1:0] sync_argumentNotifierAXI_24_RRESP;
	input sync_argumentNotifierAXI_24_RLAST;
	input sync_argumentNotifierAXI_24_AWREADY;
	output wire sync_argumentNotifierAXI_24_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_24_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_24_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_24_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_24_AWBURST;
	output wire sync_argumentNotifierAXI_24_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_24_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_24_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_24_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_24_AWREGION;
	input sync_argumentNotifierAXI_24_WREADY;
	output wire sync_argumentNotifierAXI_24_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_24_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_24_WSTRB;
	output wire sync_argumentNotifierAXI_24_WLAST;
	output wire sync_argumentNotifierAXI_24_BREADY;
	input sync_argumentNotifierAXI_24_BVALID;
	input [1:0] sync_argumentNotifierAXI_24_BRESP;
	input sync_argumentNotifierAXI_25_ARREADY;
	output wire sync_argumentNotifierAXI_25_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_25_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_25_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_25_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_25_ARBURST;
	output wire sync_argumentNotifierAXI_25_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_25_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_25_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_25_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_25_ARREGION;
	output wire sync_argumentNotifierAXI_25_RREADY;
	input sync_argumentNotifierAXI_25_RVALID;
	input [31:0] sync_argumentNotifierAXI_25_RDATA;
	input [1:0] sync_argumentNotifierAXI_25_RRESP;
	input sync_argumentNotifierAXI_25_RLAST;
	input sync_argumentNotifierAXI_25_AWREADY;
	output wire sync_argumentNotifierAXI_25_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_25_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_25_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_25_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_25_AWBURST;
	output wire sync_argumentNotifierAXI_25_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_25_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_25_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_25_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_25_AWREGION;
	input sync_argumentNotifierAXI_25_WREADY;
	output wire sync_argumentNotifierAXI_25_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_25_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_25_WSTRB;
	output wire sync_argumentNotifierAXI_25_WLAST;
	output wire sync_argumentNotifierAXI_25_BREADY;
	input sync_argumentNotifierAXI_25_BVALID;
	input [1:0] sync_argumentNotifierAXI_25_BRESP;
	input sync_argumentNotifierAXI_26_ARREADY;
	output wire sync_argumentNotifierAXI_26_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_26_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_26_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_26_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_26_ARBURST;
	output wire sync_argumentNotifierAXI_26_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_26_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_26_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_26_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_26_ARREGION;
	output wire sync_argumentNotifierAXI_26_RREADY;
	input sync_argumentNotifierAXI_26_RVALID;
	input [31:0] sync_argumentNotifierAXI_26_RDATA;
	input [1:0] sync_argumentNotifierAXI_26_RRESP;
	input sync_argumentNotifierAXI_26_RLAST;
	input sync_argumentNotifierAXI_26_AWREADY;
	output wire sync_argumentNotifierAXI_26_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_26_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_26_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_26_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_26_AWBURST;
	output wire sync_argumentNotifierAXI_26_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_26_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_26_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_26_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_26_AWREGION;
	input sync_argumentNotifierAXI_26_WREADY;
	output wire sync_argumentNotifierAXI_26_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_26_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_26_WSTRB;
	output wire sync_argumentNotifierAXI_26_WLAST;
	output wire sync_argumentNotifierAXI_26_BREADY;
	input sync_argumentNotifierAXI_26_BVALID;
	input [1:0] sync_argumentNotifierAXI_26_BRESP;
	input sync_argumentNotifierAXI_27_ARREADY;
	output wire sync_argumentNotifierAXI_27_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_27_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_27_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_27_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_27_ARBURST;
	output wire sync_argumentNotifierAXI_27_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_27_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_27_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_27_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_27_ARREGION;
	output wire sync_argumentNotifierAXI_27_RREADY;
	input sync_argumentNotifierAXI_27_RVALID;
	input [31:0] sync_argumentNotifierAXI_27_RDATA;
	input [1:0] sync_argumentNotifierAXI_27_RRESP;
	input sync_argumentNotifierAXI_27_RLAST;
	input sync_argumentNotifierAXI_27_AWREADY;
	output wire sync_argumentNotifierAXI_27_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_27_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_27_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_27_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_27_AWBURST;
	output wire sync_argumentNotifierAXI_27_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_27_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_27_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_27_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_27_AWREGION;
	input sync_argumentNotifierAXI_27_WREADY;
	output wire sync_argumentNotifierAXI_27_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_27_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_27_WSTRB;
	output wire sync_argumentNotifierAXI_27_WLAST;
	output wire sync_argumentNotifierAXI_27_BREADY;
	input sync_argumentNotifierAXI_27_BVALID;
	input [1:0] sync_argumentNotifierAXI_27_BRESP;
	input sync_argumentNotifierAXI_28_ARREADY;
	output wire sync_argumentNotifierAXI_28_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_28_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_28_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_28_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_28_ARBURST;
	output wire sync_argumentNotifierAXI_28_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_28_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_28_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_28_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_28_ARREGION;
	output wire sync_argumentNotifierAXI_28_RREADY;
	input sync_argumentNotifierAXI_28_RVALID;
	input [31:0] sync_argumentNotifierAXI_28_RDATA;
	input [1:0] sync_argumentNotifierAXI_28_RRESP;
	input sync_argumentNotifierAXI_28_RLAST;
	input sync_argumentNotifierAXI_28_AWREADY;
	output wire sync_argumentNotifierAXI_28_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_28_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_28_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_28_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_28_AWBURST;
	output wire sync_argumentNotifierAXI_28_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_28_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_28_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_28_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_28_AWREGION;
	input sync_argumentNotifierAXI_28_WREADY;
	output wire sync_argumentNotifierAXI_28_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_28_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_28_WSTRB;
	output wire sync_argumentNotifierAXI_28_WLAST;
	output wire sync_argumentNotifierAXI_28_BREADY;
	input sync_argumentNotifierAXI_28_BVALID;
	input [1:0] sync_argumentNotifierAXI_28_BRESP;
	input sync_argumentNotifierAXI_29_ARREADY;
	output wire sync_argumentNotifierAXI_29_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_29_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_29_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_29_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_29_ARBURST;
	output wire sync_argumentNotifierAXI_29_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_29_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_29_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_29_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_29_ARREGION;
	output wire sync_argumentNotifierAXI_29_RREADY;
	input sync_argumentNotifierAXI_29_RVALID;
	input [31:0] sync_argumentNotifierAXI_29_RDATA;
	input [1:0] sync_argumentNotifierAXI_29_RRESP;
	input sync_argumentNotifierAXI_29_RLAST;
	input sync_argumentNotifierAXI_29_AWREADY;
	output wire sync_argumentNotifierAXI_29_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_29_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_29_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_29_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_29_AWBURST;
	output wire sync_argumentNotifierAXI_29_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_29_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_29_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_29_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_29_AWREGION;
	input sync_argumentNotifierAXI_29_WREADY;
	output wire sync_argumentNotifierAXI_29_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_29_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_29_WSTRB;
	output wire sync_argumentNotifierAXI_29_WLAST;
	output wire sync_argumentNotifierAXI_29_BREADY;
	input sync_argumentNotifierAXI_29_BVALID;
	input [1:0] sync_argumentNotifierAXI_29_BRESP;
	input sync_argumentNotifierAXI_30_ARREADY;
	output wire sync_argumentNotifierAXI_30_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_30_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_30_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_30_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_30_ARBURST;
	output wire sync_argumentNotifierAXI_30_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_30_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_30_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_30_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_30_ARREGION;
	output wire sync_argumentNotifierAXI_30_RREADY;
	input sync_argumentNotifierAXI_30_RVALID;
	input [31:0] sync_argumentNotifierAXI_30_RDATA;
	input [1:0] sync_argumentNotifierAXI_30_RRESP;
	input sync_argumentNotifierAXI_30_RLAST;
	input sync_argumentNotifierAXI_30_AWREADY;
	output wire sync_argumentNotifierAXI_30_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_30_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_30_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_30_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_30_AWBURST;
	output wire sync_argumentNotifierAXI_30_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_30_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_30_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_30_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_30_AWREGION;
	input sync_argumentNotifierAXI_30_WREADY;
	output wire sync_argumentNotifierAXI_30_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_30_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_30_WSTRB;
	output wire sync_argumentNotifierAXI_30_WLAST;
	output wire sync_argumentNotifierAXI_30_BREADY;
	input sync_argumentNotifierAXI_30_BVALID;
	input [1:0] sync_argumentNotifierAXI_30_BRESP;
	input sync_argumentNotifierAXI_31_ARREADY;
	output wire sync_argumentNotifierAXI_31_ARVALID;
	output wire [63:0] sync_argumentNotifierAXI_31_ARADDR;
	output wire [7:0] sync_argumentNotifierAXI_31_ARLEN;
	output wire [2:0] sync_argumentNotifierAXI_31_ARSIZE;
	output wire [1:0] sync_argumentNotifierAXI_31_ARBURST;
	output wire sync_argumentNotifierAXI_31_ARLOCK;
	output wire [3:0] sync_argumentNotifierAXI_31_ARCACHE;
	output wire [2:0] sync_argumentNotifierAXI_31_ARPROT;
	output wire [3:0] sync_argumentNotifierAXI_31_ARQOS;
	output wire [3:0] sync_argumentNotifierAXI_31_ARREGION;
	output wire sync_argumentNotifierAXI_31_RREADY;
	input sync_argumentNotifierAXI_31_RVALID;
	input [31:0] sync_argumentNotifierAXI_31_RDATA;
	input [1:0] sync_argumentNotifierAXI_31_RRESP;
	input sync_argumentNotifierAXI_31_RLAST;
	input sync_argumentNotifierAXI_31_AWREADY;
	output wire sync_argumentNotifierAXI_31_AWVALID;
	output wire [63:0] sync_argumentNotifierAXI_31_AWADDR;
	output wire [7:0] sync_argumentNotifierAXI_31_AWLEN;
	output wire [2:0] sync_argumentNotifierAXI_31_AWSIZE;
	output wire [1:0] sync_argumentNotifierAXI_31_AWBURST;
	output wire sync_argumentNotifierAXI_31_AWLOCK;
	output wire [3:0] sync_argumentNotifierAXI_31_AWCACHE;
	output wire [2:0] sync_argumentNotifierAXI_31_AWPROT;
	output wire [3:0] sync_argumentNotifierAXI_31_AWQOS;
	output wire [3:0] sync_argumentNotifierAXI_31_AWREGION;
	input sync_argumentNotifierAXI_31_WREADY;
	output wire sync_argumentNotifierAXI_31_WVALID;
	output wire [31:0] sync_argumentNotifierAXI_31_WDATA;
	output wire [3:0] sync_argumentNotifierAXI_31_WSTRB;
	output wire sync_argumentNotifierAXI_31_WLAST;
	output wire sync_argumentNotifierAXI_31_BREADY;
	input sync_argumentNotifierAXI_31_BVALID;
	input [1:0] sync_argumentNotifierAXI_31_BRESP;
	wire _ArgumentNotifier_io_export_argIn_0_TREADY;
	wire _ArgumentNotifier_io_export_argIn_1_TREADY;
	wire _ArgumentNotifier_io_export_argIn_2_TREADY;
	wire _ArgumentNotifier_io_export_argIn_3_TREADY;
	wire _ArgumentNotifier_io_export_argIn_4_TREADY;
	wire _ArgumentNotifier_io_export_argIn_5_TREADY;
	wire _ArgumentNotifier_io_export_argIn_6_TREADY;
	wire _ArgumentNotifier_io_export_argIn_7_TREADY;
	wire _ArgumentNotifier_io_export_argIn_8_TREADY;
	wire _ArgumentNotifier_io_export_argIn_9_TREADY;
	wire _ArgumentNotifier_io_export_argIn_10_TREADY;
	wire _ArgumentNotifier_io_export_argIn_11_TREADY;
	wire _ArgumentNotifier_io_export_argIn_12_TREADY;
	wire _ArgumentNotifier_io_export_argIn_13_TREADY;
	wire _ArgumentNotifier_io_export_argIn_14_TREADY;
	wire _ArgumentNotifier_io_export_argIn_15_TREADY;
	wire _ArgumentNotifier_io_export_argIn_16_TREADY;
	wire _ArgumentNotifier_io_export_argIn_17_TREADY;
	wire _ArgumentNotifier_io_export_argIn_18_TREADY;
	wire _ArgumentNotifier_io_export_argIn_19_TREADY;
	wire _ArgumentNotifier_io_export_argIn_20_TREADY;
	wire _ArgumentNotifier_io_export_argIn_21_TREADY;
	wire _ArgumentNotifier_io_export_argIn_22_TREADY;
	wire _ArgumentNotifier_io_export_argIn_23_TREADY;
	wire _ArgumentNotifier_io_export_argIn_24_TREADY;
	wire _ArgumentNotifier_io_export_argIn_25_TREADY;
	wire _ArgumentNotifier_io_export_argIn_26_TREADY;
	wire _ArgumentNotifier_io_export_argIn_27_TREADY;
	wire _ArgumentNotifier_io_export_argIn_28_TREADY;
	wire _ArgumentNotifier_io_export_argIn_29_TREADY;
	wire _ArgumentNotifier_io_export_argIn_30_TREADY;
	wire _ArgumentNotifier_io_export_argIn_31_TREADY;
	wire _ArgumentNotifier_io_export_argIn_32_TREADY;
	wire _ArgumentNotifier_io_export_argIn_33_TREADY;
	wire _ArgumentNotifier_io_export_argIn_34_TREADY;
	wire _ArgumentNotifier_io_export_argIn_35_TREADY;
	wire _ArgumentNotifier_io_export_argIn_36_TREADY;
	wire _ArgumentNotifier_io_export_argIn_37_TREADY;
	wire _ArgumentNotifier_io_export_argIn_38_TREADY;
	wire _ArgumentNotifier_io_export_argIn_39_TREADY;
	wire _ArgumentNotifier_io_export_argIn_40_TREADY;
	wire _ArgumentNotifier_io_export_argIn_41_TREADY;
	wire _ArgumentNotifier_io_export_argIn_42_TREADY;
	wire _ArgumentNotifier_io_export_argIn_43_TREADY;
	wire _ArgumentNotifier_io_export_argIn_44_TREADY;
	wire _ArgumentNotifier_io_export_argIn_45_TREADY;
	wire _ArgumentNotifier_io_export_argIn_46_TREADY;
	wire _ArgumentNotifier_io_export_argIn_47_TREADY;
	wire _ArgumentNotifier_io_export_argIn_48_TREADY;
	wire _ArgumentNotifier_io_export_argIn_49_TREADY;
	wire _ArgumentNotifier_io_export_argIn_50_TREADY;
	wire _ArgumentNotifier_io_export_argIn_51_TREADY;
	wire _ArgumentNotifier_io_export_argIn_52_TREADY;
	wire _ArgumentNotifier_io_export_argIn_53_TREADY;
	wire _ArgumentNotifier_io_export_argIn_54_TREADY;
	wire _ArgumentNotifier_io_export_argIn_55_TREADY;
	wire _ArgumentNotifier_io_export_argIn_56_TREADY;
	wire _ArgumentNotifier_io_export_argIn_57_TREADY;
	wire _ArgumentNotifier_io_export_argIn_58_TREADY;
	wire _ArgumentNotifier_io_export_argIn_59_TREADY;
	wire _ArgumentNotifier_io_export_argIn_60_TREADY;
	wire _ArgumentNotifier_io_export_argIn_61_TREADY;
	wire _ArgumentNotifier_io_export_argIn_62_TREADY;
	wire _ArgumentNotifier_io_export_argIn_63_TREADY;
	wire _ArgumentNotifier_io_export_argIn_64_TREADY;
	wire _ArgumentNotifier_io_export_argIn_65_TREADY;
	wire _ArgumentNotifier_io_export_argIn_66_TREADY;
	wire _ArgumentNotifier_io_export_argIn_67_TREADY;
	wire _ArgumentNotifier_io_export_argIn_68_TREADY;
	wire _ArgumentNotifier_io_export_argIn_69_TREADY;
	wire _ArgumentNotifier_io_export_argIn_70_TREADY;
	wire _ArgumentNotifier_io_export_argIn_71_TREADY;
	wire _ArgumentNotifier_io_export_argIn_72_TREADY;
	wire _ArgumentNotifier_io_export_argIn_73_TREADY;
	wire _ArgumentNotifier_io_export_argIn_74_TREADY;
	wire _ArgumentNotifier_io_export_argIn_75_TREADY;
	wire _ArgumentNotifier_io_export_argIn_76_TREADY;
	wire _ArgumentNotifier_io_export_argIn_77_TREADY;
	wire _ArgumentNotifier_io_export_argIn_78_TREADY;
	wire _ArgumentNotifier_io_export_argIn_79_TREADY;
	wire _ArgumentNotifier_connStealNtw_0_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_0_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_0_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_1_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_1_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_1_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_2_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_2_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_2_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_3_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_3_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_3_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_4_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_4_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_4_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_5_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_5_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_5_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_6_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_6_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_6_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_7_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_7_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_7_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_8_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_8_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_8_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_9_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_9_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_9_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_10_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_10_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_10_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_11_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_11_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_11_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_12_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_12_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_12_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_13_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_13_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_13_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_14_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_14_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_14_data_qOutTask_bits;
	wire _ArgumentNotifier_connStealNtw_15_ctrl_serveStealReq_valid;
	wire _ArgumentNotifier_connStealNtw_15_data_qOutTask_valid;
	wire [127:0] _ArgumentNotifier_connStealNtw_15_data_qOutTask_bits;
	wire _Allocator_io_export_closureOut_0_TVALID;
	wire _Allocator_io_export_closureOut_1_TVALID;
	wire _Allocator_io_export_closureOut_2_TVALID;
	wire _Allocator_io_export_closureOut_3_TVALID;
	wire _Allocator_io_export_closureOut_4_TVALID;
	wire _Allocator_io_export_closureOut_5_TVALID;
	wire _Allocator_io_export_closureOut_6_TVALID;
	wire _Allocator_io_export_closureOut_7_TVALID;
	wire _Allocator_io_export_closureOut_8_TVALID;
	wire _Allocator_io_export_closureOut_9_TVALID;
	wire _Allocator_io_export_closureOut_10_TVALID;
	wire _Allocator_io_export_closureOut_11_TVALID;
	wire _Allocator_io_export_closureOut_12_TVALID;
	wire _Allocator_io_export_closureOut_13_TVALID;
	wire _Allocator_io_export_closureOut_14_TVALID;
	wire _Allocator_io_export_closureOut_15_TVALID;
	wire _Allocator_io_export_closureOut_16_TVALID;
	wire _Allocator_io_export_closureOut_17_TVALID;
	wire _Allocator_io_export_closureOut_18_TVALID;
	wire _Allocator_io_export_closureOut_19_TVALID;
	wire _Allocator_io_export_closureOut_20_TVALID;
	wire _Allocator_io_export_closureOut_21_TVALID;
	wire _Allocator_io_export_closureOut_22_TVALID;
	wire _Allocator_io_export_closureOut_23_TVALID;
	wire _Allocator_io_export_closureOut_24_TVALID;
	wire _Allocator_io_export_closureOut_25_TVALID;
	wire _Allocator_io_export_closureOut_26_TVALID;
	wire _Allocator_io_export_closureOut_27_TVALID;
	wire _Allocator_io_export_closureOut_28_TVALID;
	wire _Allocator_io_export_closureOut_29_TVALID;
	wire _Allocator_io_export_closureOut_30_TVALID;
	wire _Allocator_io_export_closureOut_31_TVALID;
	wire _Allocator_io_export_closureOut_32_TVALID;
	wire _Allocator_io_export_closureOut_33_TVALID;
	wire _Allocator_io_export_closureOut_34_TVALID;
	wire _Allocator_io_export_closureOut_35_TVALID;
	wire _Allocator_io_export_closureOut_36_TVALID;
	wire _Allocator_io_export_closureOut_37_TVALID;
	wire _Allocator_io_export_closureOut_38_TVALID;
	wire _Allocator_io_export_closureOut_39_TVALID;
	wire _Allocator_io_export_closureOut_40_TVALID;
	wire _Allocator_io_export_closureOut_41_TVALID;
	wire _Allocator_io_export_closureOut_42_TVALID;
	wire _Allocator_io_export_closureOut_43_TVALID;
	wire _Allocator_io_export_closureOut_44_TVALID;
	wire _Allocator_io_export_closureOut_45_TVALID;
	wire _Allocator_io_export_closureOut_46_TVALID;
	wire _Allocator_io_export_closureOut_47_TVALID;
	wire _Allocator_io_export_closureOut_48_TVALID;
	wire _Allocator_io_export_closureOut_49_TVALID;
	wire _Allocator_io_export_closureOut_50_TVALID;
	wire _Allocator_io_export_closureOut_51_TVALID;
	wire _Allocator_io_export_closureOut_52_TVALID;
	wire _Allocator_io_export_closureOut_53_TVALID;
	wire _Allocator_io_export_closureOut_54_TVALID;
	wire _Allocator_io_export_closureOut_55_TVALID;
	wire _Allocator_io_export_closureOut_56_TVALID;
	wire _Allocator_io_export_closureOut_57_TVALID;
	wire _Allocator_io_export_closureOut_58_TVALID;
	wire _Allocator_io_export_closureOut_59_TVALID;
	wire _Allocator_io_export_closureOut_60_TVALID;
	wire _Allocator_io_export_closureOut_61_TVALID;
	wire _Allocator_io_export_closureOut_62_TVALID;
	wire _Allocator_io_export_closureOut_63_TVALID;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_0_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_0_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_0_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_0_b_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_1_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_1_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_1_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_1_b_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_2_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_2_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_2_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_2_b_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_ar_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_r_valid;
	wire [63:0] _Allocator_io_internal_axi_mgmt_vcas_3_r_bits_data;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_3_r_bits_resp;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_aw_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_w_ready;
	wire _Allocator_io_internal_axi_mgmt_vcas_3_b_valid;
	wire [1:0] _Allocator_io_internal_axi_mgmt_vcas_3_b_bits_resp;
	wire _Scheduler_1_io_export_taskOut_0_TVALID;
	wire _Scheduler_1_io_export_taskOut_1_TVALID;
	wire _Scheduler_1_io_export_taskOut_2_TVALID;
	wire _Scheduler_1_io_export_taskOut_3_TVALID;
	wire _Scheduler_1_io_export_taskOut_4_TVALID;
	wire _Scheduler_1_io_export_taskOut_5_TVALID;
	wire _Scheduler_1_io_export_taskOut_6_TVALID;
	wire _Scheduler_1_io_export_taskOut_7_TVALID;
	wire _Scheduler_1_io_export_taskOut_8_TVALID;
	wire _Scheduler_1_io_export_taskOut_9_TVALID;
	wire _Scheduler_1_io_export_taskOut_10_TVALID;
	wire _Scheduler_1_io_export_taskOut_11_TVALID;
	wire _Scheduler_1_io_export_taskOut_12_TVALID;
	wire _Scheduler_1_io_export_taskOut_13_TVALID;
	wire _Scheduler_1_io_export_taskOut_14_TVALID;
	wire _Scheduler_1_io_export_taskOut_15_TVALID;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_ar_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_r_valid;
	wire [63:0] _Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_data;
	wire [1:0] _Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_resp;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_aw_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_w_ready;
	wire _Scheduler_1_io_internal_axi_mgmt_vss_0_b_valid;
	wire [1:0] _Scheduler_1_io_internal_axi_mgmt_vss_0_b_bits_resp;
	wire _Scheduler_1_connArgumentNotifier_0_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_0_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_1_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_1_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_2_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_2_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_3_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_3_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_4_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_4_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_5_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_5_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_6_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_6_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_7_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_7_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_8_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_8_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_9_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_9_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_10_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_10_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_11_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_11_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_12_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_12_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_13_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_13_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_14_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_14_data_qOutTask_ready;
	wire _Scheduler_1_connArgumentNotifier_15_ctrl_serveStealReq_ready;
	wire _Scheduler_1_connArgumentNotifier_15_data_qOutTask_ready;
	wire _peArray_15_1_argOut_TVALID;
	wire [63:0] _peArray_15_1_argOut_TDATA;
	wire _peArray_15_1_taskIn_TREADY;
	wire _peArray_14_1_argOut_TVALID;
	wire [63:0] _peArray_14_1_argOut_TDATA;
	wire _peArray_14_1_taskIn_TREADY;
	wire _peArray_13_1_argOut_TVALID;
	wire [63:0] _peArray_13_1_argOut_TDATA;
	wire _peArray_13_1_taskIn_TREADY;
	wire _peArray_12_1_argOut_TVALID;
	wire [63:0] _peArray_12_1_argOut_TDATA;
	wire _peArray_12_1_taskIn_TREADY;
	wire _peArray_11_1_argOut_TVALID;
	wire [63:0] _peArray_11_1_argOut_TDATA;
	wire _peArray_11_1_taskIn_TREADY;
	wire _peArray_10_1_argOut_TVALID;
	wire [63:0] _peArray_10_1_argOut_TDATA;
	wire _peArray_10_1_taskIn_TREADY;
	wire _peArray_9_1_argOut_TVALID;
	wire [63:0] _peArray_9_1_argOut_TDATA;
	wire _peArray_9_1_taskIn_TREADY;
	wire _peArray_8_1_argOut_TVALID;
	wire [63:0] _peArray_8_1_argOut_TDATA;
	wire _peArray_8_1_taskIn_TREADY;
	wire _peArray_7_1_argOut_TVALID;
	wire [63:0] _peArray_7_1_argOut_TDATA;
	wire _peArray_7_1_taskIn_TREADY;
	wire _peArray_6_1_argOut_TVALID;
	wire [63:0] _peArray_6_1_argOut_TDATA;
	wire _peArray_6_1_taskIn_TREADY;
	wire _peArray_5_1_argOut_TVALID;
	wire [63:0] _peArray_5_1_argOut_TDATA;
	wire _peArray_5_1_taskIn_TREADY;
	wire _peArray_4_1_argOut_TVALID;
	wire [63:0] _peArray_4_1_argOut_TDATA;
	wire _peArray_4_1_taskIn_TREADY;
	wire _peArray_3_1_argOut_TVALID;
	wire [63:0] _peArray_3_1_argOut_TDATA;
	wire _peArray_3_1_taskIn_TREADY;
	wire _peArray_2_1_argOut_TVALID;
	wire [63:0] _peArray_2_1_argOut_TDATA;
	wire _peArray_2_1_taskIn_TREADY;
	wire _peArray_1_1_argOut_TVALID;
	wire [63:0] _peArray_1_1_argOut_TDATA;
	wire _peArray_1_1_taskIn_TREADY;
	wire _peArray_0_1_argOut_TVALID;
	wire [63:0] _peArray_0_1_argOut_TDATA;
	wire _peArray_0_1_taskIn_TREADY;
	wire _Scheduler_io_export_taskOut_0_TVALID;
	wire _Scheduler_io_export_taskOut_1_TVALID;
	wire _Scheduler_io_export_taskOut_2_TVALID;
	wire _Scheduler_io_export_taskOut_3_TVALID;
	wire _Scheduler_io_export_taskOut_4_TVALID;
	wire _Scheduler_io_export_taskOut_5_TVALID;
	wire _Scheduler_io_export_taskOut_6_TVALID;
	wire _Scheduler_io_export_taskOut_7_TVALID;
	wire _Scheduler_io_export_taskOut_8_TVALID;
	wire _Scheduler_io_export_taskOut_9_TVALID;
	wire _Scheduler_io_export_taskOut_10_TVALID;
	wire _Scheduler_io_export_taskOut_11_TVALID;
	wire _Scheduler_io_export_taskOut_12_TVALID;
	wire _Scheduler_io_export_taskOut_13_TVALID;
	wire _Scheduler_io_export_taskOut_14_TVALID;
	wire _Scheduler_io_export_taskOut_15_TVALID;
	wire _Scheduler_io_export_taskOut_16_TVALID;
	wire _Scheduler_io_export_taskOut_17_TVALID;
	wire _Scheduler_io_export_taskOut_18_TVALID;
	wire _Scheduler_io_export_taskOut_19_TVALID;
	wire _Scheduler_io_export_taskOut_20_TVALID;
	wire _Scheduler_io_export_taskOut_21_TVALID;
	wire _Scheduler_io_export_taskOut_22_TVALID;
	wire _Scheduler_io_export_taskOut_23_TVALID;
	wire _Scheduler_io_export_taskOut_24_TVALID;
	wire _Scheduler_io_export_taskOut_25_TVALID;
	wire _Scheduler_io_export_taskOut_26_TVALID;
	wire _Scheduler_io_export_taskOut_27_TVALID;
	wire _Scheduler_io_export_taskOut_28_TVALID;
	wire _Scheduler_io_export_taskOut_29_TVALID;
	wire _Scheduler_io_export_taskOut_30_TVALID;
	wire _Scheduler_io_export_taskOut_31_TVALID;
	wire _Scheduler_io_export_taskOut_32_TVALID;
	wire _Scheduler_io_export_taskOut_33_TVALID;
	wire _Scheduler_io_export_taskOut_34_TVALID;
	wire _Scheduler_io_export_taskOut_35_TVALID;
	wire _Scheduler_io_export_taskOut_36_TVALID;
	wire _Scheduler_io_export_taskOut_37_TVALID;
	wire _Scheduler_io_export_taskOut_38_TVALID;
	wire _Scheduler_io_export_taskOut_39_TVALID;
	wire _Scheduler_io_export_taskOut_40_TVALID;
	wire _Scheduler_io_export_taskOut_41_TVALID;
	wire _Scheduler_io_export_taskOut_42_TVALID;
	wire _Scheduler_io_export_taskOut_43_TVALID;
	wire _Scheduler_io_export_taskOut_44_TVALID;
	wire _Scheduler_io_export_taskOut_45_TVALID;
	wire _Scheduler_io_export_taskOut_46_TVALID;
	wire _Scheduler_io_export_taskOut_47_TVALID;
	wire _Scheduler_io_export_taskOut_48_TVALID;
	wire _Scheduler_io_export_taskOut_49_TVALID;
	wire _Scheduler_io_export_taskOut_50_TVALID;
	wire _Scheduler_io_export_taskOut_51_TVALID;
	wire _Scheduler_io_export_taskOut_52_TVALID;
	wire _Scheduler_io_export_taskOut_53_TVALID;
	wire _Scheduler_io_export_taskOut_54_TVALID;
	wire _Scheduler_io_export_taskOut_55_TVALID;
	wire _Scheduler_io_export_taskOut_56_TVALID;
	wire _Scheduler_io_export_taskOut_57_TVALID;
	wire _Scheduler_io_export_taskOut_58_TVALID;
	wire _Scheduler_io_export_taskOut_59_TVALID;
	wire _Scheduler_io_export_taskOut_60_TVALID;
	wire _Scheduler_io_export_taskOut_61_TVALID;
	wire _Scheduler_io_export_taskOut_62_TVALID;
	wire _Scheduler_io_export_taskOut_63_TVALID;
	wire _Scheduler_io_export_taskIn_0_TREADY;
	wire _Scheduler_io_export_taskIn_1_TREADY;
	wire _Scheduler_io_export_taskIn_2_TREADY;
	wire _Scheduler_io_export_taskIn_3_TREADY;
	wire _Scheduler_io_export_taskIn_4_TREADY;
	wire _Scheduler_io_export_taskIn_5_TREADY;
	wire _Scheduler_io_export_taskIn_6_TREADY;
	wire _Scheduler_io_export_taskIn_7_TREADY;
	wire _Scheduler_io_export_taskIn_8_TREADY;
	wire _Scheduler_io_export_taskIn_9_TREADY;
	wire _Scheduler_io_export_taskIn_10_TREADY;
	wire _Scheduler_io_export_taskIn_11_TREADY;
	wire _Scheduler_io_export_taskIn_12_TREADY;
	wire _Scheduler_io_export_taskIn_13_TREADY;
	wire _Scheduler_io_export_taskIn_14_TREADY;
	wire _Scheduler_io_export_taskIn_15_TREADY;
	wire _Scheduler_io_export_taskIn_16_TREADY;
	wire _Scheduler_io_export_taskIn_17_TREADY;
	wire _Scheduler_io_export_taskIn_18_TREADY;
	wire _Scheduler_io_export_taskIn_19_TREADY;
	wire _Scheduler_io_export_taskIn_20_TREADY;
	wire _Scheduler_io_export_taskIn_21_TREADY;
	wire _Scheduler_io_export_taskIn_22_TREADY;
	wire _Scheduler_io_export_taskIn_23_TREADY;
	wire _Scheduler_io_export_taskIn_24_TREADY;
	wire _Scheduler_io_export_taskIn_25_TREADY;
	wire _Scheduler_io_export_taskIn_26_TREADY;
	wire _Scheduler_io_export_taskIn_27_TREADY;
	wire _Scheduler_io_export_taskIn_28_TREADY;
	wire _Scheduler_io_export_taskIn_29_TREADY;
	wire _Scheduler_io_export_taskIn_30_TREADY;
	wire _Scheduler_io_export_taskIn_31_TREADY;
	wire _Scheduler_io_export_taskIn_32_TREADY;
	wire _Scheduler_io_export_taskIn_33_TREADY;
	wire _Scheduler_io_export_taskIn_34_TREADY;
	wire _Scheduler_io_export_taskIn_35_TREADY;
	wire _Scheduler_io_export_taskIn_36_TREADY;
	wire _Scheduler_io_export_taskIn_37_TREADY;
	wire _Scheduler_io_export_taskIn_38_TREADY;
	wire _Scheduler_io_export_taskIn_39_TREADY;
	wire _Scheduler_io_export_taskIn_40_TREADY;
	wire _Scheduler_io_export_taskIn_41_TREADY;
	wire _Scheduler_io_export_taskIn_42_TREADY;
	wire _Scheduler_io_export_taskIn_43_TREADY;
	wire _Scheduler_io_export_taskIn_44_TREADY;
	wire _Scheduler_io_export_taskIn_45_TREADY;
	wire _Scheduler_io_export_taskIn_46_TREADY;
	wire _Scheduler_io_export_taskIn_47_TREADY;
	wire _Scheduler_io_export_taskIn_48_TREADY;
	wire _Scheduler_io_export_taskIn_49_TREADY;
	wire _Scheduler_io_export_taskIn_50_TREADY;
	wire _Scheduler_io_export_taskIn_51_TREADY;
	wire _Scheduler_io_export_taskIn_52_TREADY;
	wire _Scheduler_io_export_taskIn_53_TREADY;
	wire _Scheduler_io_export_taskIn_54_TREADY;
	wire _Scheduler_io_export_taskIn_55_TREADY;
	wire _Scheduler_io_export_taskIn_56_TREADY;
	wire _Scheduler_io_export_taskIn_57_TREADY;
	wire _Scheduler_io_export_taskIn_58_TREADY;
	wire _Scheduler_io_export_taskIn_59_TREADY;
	wire _Scheduler_io_export_taskIn_60_TREADY;
	wire _Scheduler_io_export_taskIn_61_TREADY;
	wire _Scheduler_io_export_taskIn_62_TREADY;
	wire _Scheduler_io_export_taskIn_63_TREADY;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_ar_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_r_valid;
	wire [63:0] _Scheduler_io_internal_axi_mgmt_vss_0_r_bits_data;
	wire [1:0] _Scheduler_io_internal_axi_mgmt_vss_0_r_bits_resp;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_aw_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_w_ready;
	wire _Scheduler_io_internal_axi_mgmt_vss_0_b_valid;
	wire [1:0] _Scheduler_io_internal_axi_mgmt_vss_0_b_bits_resp;
	wire _peArray_63_closureIn_TREADY;
	wire _peArray_63_argOut_TVALID;
	wire [63:0] _peArray_63_argOut_TDATA;
	wire _peArray_63_taskOut_TVALID;
	wire [255:0] _peArray_63_taskOut_TDATA;
	wire _peArray_63_taskIn_TREADY;
	wire _peArray_62_closureIn_TREADY;
	wire _peArray_62_argOut_TVALID;
	wire [63:0] _peArray_62_argOut_TDATA;
	wire _peArray_62_taskOut_TVALID;
	wire [255:0] _peArray_62_taskOut_TDATA;
	wire _peArray_62_taskIn_TREADY;
	wire _peArray_61_closureIn_TREADY;
	wire _peArray_61_argOut_TVALID;
	wire [63:0] _peArray_61_argOut_TDATA;
	wire _peArray_61_taskOut_TVALID;
	wire [255:0] _peArray_61_taskOut_TDATA;
	wire _peArray_61_taskIn_TREADY;
	wire _peArray_60_closureIn_TREADY;
	wire _peArray_60_argOut_TVALID;
	wire [63:0] _peArray_60_argOut_TDATA;
	wire _peArray_60_taskOut_TVALID;
	wire [255:0] _peArray_60_taskOut_TDATA;
	wire _peArray_60_taskIn_TREADY;
	wire _peArray_59_closureIn_TREADY;
	wire _peArray_59_argOut_TVALID;
	wire [63:0] _peArray_59_argOut_TDATA;
	wire _peArray_59_taskOut_TVALID;
	wire [255:0] _peArray_59_taskOut_TDATA;
	wire _peArray_59_taskIn_TREADY;
	wire _peArray_58_closureIn_TREADY;
	wire _peArray_58_argOut_TVALID;
	wire [63:0] _peArray_58_argOut_TDATA;
	wire _peArray_58_taskOut_TVALID;
	wire [255:0] _peArray_58_taskOut_TDATA;
	wire _peArray_58_taskIn_TREADY;
	wire _peArray_57_closureIn_TREADY;
	wire _peArray_57_argOut_TVALID;
	wire [63:0] _peArray_57_argOut_TDATA;
	wire _peArray_57_taskOut_TVALID;
	wire [255:0] _peArray_57_taskOut_TDATA;
	wire _peArray_57_taskIn_TREADY;
	wire _peArray_56_closureIn_TREADY;
	wire _peArray_56_argOut_TVALID;
	wire [63:0] _peArray_56_argOut_TDATA;
	wire _peArray_56_taskOut_TVALID;
	wire [255:0] _peArray_56_taskOut_TDATA;
	wire _peArray_56_taskIn_TREADY;
	wire _peArray_55_closureIn_TREADY;
	wire _peArray_55_argOut_TVALID;
	wire [63:0] _peArray_55_argOut_TDATA;
	wire _peArray_55_taskOut_TVALID;
	wire [255:0] _peArray_55_taskOut_TDATA;
	wire _peArray_55_taskIn_TREADY;
	wire _peArray_54_closureIn_TREADY;
	wire _peArray_54_argOut_TVALID;
	wire [63:0] _peArray_54_argOut_TDATA;
	wire _peArray_54_taskOut_TVALID;
	wire [255:0] _peArray_54_taskOut_TDATA;
	wire _peArray_54_taskIn_TREADY;
	wire _peArray_53_closureIn_TREADY;
	wire _peArray_53_argOut_TVALID;
	wire [63:0] _peArray_53_argOut_TDATA;
	wire _peArray_53_taskOut_TVALID;
	wire [255:0] _peArray_53_taskOut_TDATA;
	wire _peArray_53_taskIn_TREADY;
	wire _peArray_52_closureIn_TREADY;
	wire _peArray_52_argOut_TVALID;
	wire [63:0] _peArray_52_argOut_TDATA;
	wire _peArray_52_taskOut_TVALID;
	wire [255:0] _peArray_52_taskOut_TDATA;
	wire _peArray_52_taskIn_TREADY;
	wire _peArray_51_closureIn_TREADY;
	wire _peArray_51_argOut_TVALID;
	wire [63:0] _peArray_51_argOut_TDATA;
	wire _peArray_51_taskOut_TVALID;
	wire [255:0] _peArray_51_taskOut_TDATA;
	wire _peArray_51_taskIn_TREADY;
	wire _peArray_50_closureIn_TREADY;
	wire _peArray_50_argOut_TVALID;
	wire [63:0] _peArray_50_argOut_TDATA;
	wire _peArray_50_taskOut_TVALID;
	wire [255:0] _peArray_50_taskOut_TDATA;
	wire _peArray_50_taskIn_TREADY;
	wire _peArray_49_closureIn_TREADY;
	wire _peArray_49_argOut_TVALID;
	wire [63:0] _peArray_49_argOut_TDATA;
	wire _peArray_49_taskOut_TVALID;
	wire [255:0] _peArray_49_taskOut_TDATA;
	wire _peArray_49_taskIn_TREADY;
	wire _peArray_48_closureIn_TREADY;
	wire _peArray_48_argOut_TVALID;
	wire [63:0] _peArray_48_argOut_TDATA;
	wire _peArray_48_taskOut_TVALID;
	wire [255:0] _peArray_48_taskOut_TDATA;
	wire _peArray_48_taskIn_TREADY;
	wire _peArray_47_closureIn_TREADY;
	wire _peArray_47_argOut_TVALID;
	wire [63:0] _peArray_47_argOut_TDATA;
	wire _peArray_47_taskOut_TVALID;
	wire [255:0] _peArray_47_taskOut_TDATA;
	wire _peArray_47_taskIn_TREADY;
	wire _peArray_46_closureIn_TREADY;
	wire _peArray_46_argOut_TVALID;
	wire [63:0] _peArray_46_argOut_TDATA;
	wire _peArray_46_taskOut_TVALID;
	wire [255:0] _peArray_46_taskOut_TDATA;
	wire _peArray_46_taskIn_TREADY;
	wire _peArray_45_closureIn_TREADY;
	wire _peArray_45_argOut_TVALID;
	wire [63:0] _peArray_45_argOut_TDATA;
	wire _peArray_45_taskOut_TVALID;
	wire [255:0] _peArray_45_taskOut_TDATA;
	wire _peArray_45_taskIn_TREADY;
	wire _peArray_44_closureIn_TREADY;
	wire _peArray_44_argOut_TVALID;
	wire [63:0] _peArray_44_argOut_TDATA;
	wire _peArray_44_taskOut_TVALID;
	wire [255:0] _peArray_44_taskOut_TDATA;
	wire _peArray_44_taskIn_TREADY;
	wire _peArray_43_closureIn_TREADY;
	wire _peArray_43_argOut_TVALID;
	wire [63:0] _peArray_43_argOut_TDATA;
	wire _peArray_43_taskOut_TVALID;
	wire [255:0] _peArray_43_taskOut_TDATA;
	wire _peArray_43_taskIn_TREADY;
	wire _peArray_42_closureIn_TREADY;
	wire _peArray_42_argOut_TVALID;
	wire [63:0] _peArray_42_argOut_TDATA;
	wire _peArray_42_taskOut_TVALID;
	wire [255:0] _peArray_42_taskOut_TDATA;
	wire _peArray_42_taskIn_TREADY;
	wire _peArray_41_closureIn_TREADY;
	wire _peArray_41_argOut_TVALID;
	wire [63:0] _peArray_41_argOut_TDATA;
	wire _peArray_41_taskOut_TVALID;
	wire [255:0] _peArray_41_taskOut_TDATA;
	wire _peArray_41_taskIn_TREADY;
	wire _peArray_40_closureIn_TREADY;
	wire _peArray_40_argOut_TVALID;
	wire [63:0] _peArray_40_argOut_TDATA;
	wire _peArray_40_taskOut_TVALID;
	wire [255:0] _peArray_40_taskOut_TDATA;
	wire _peArray_40_taskIn_TREADY;
	wire _peArray_39_closureIn_TREADY;
	wire _peArray_39_argOut_TVALID;
	wire [63:0] _peArray_39_argOut_TDATA;
	wire _peArray_39_taskOut_TVALID;
	wire [255:0] _peArray_39_taskOut_TDATA;
	wire _peArray_39_taskIn_TREADY;
	wire _peArray_38_closureIn_TREADY;
	wire _peArray_38_argOut_TVALID;
	wire [63:0] _peArray_38_argOut_TDATA;
	wire _peArray_38_taskOut_TVALID;
	wire [255:0] _peArray_38_taskOut_TDATA;
	wire _peArray_38_taskIn_TREADY;
	wire _peArray_37_closureIn_TREADY;
	wire _peArray_37_argOut_TVALID;
	wire [63:0] _peArray_37_argOut_TDATA;
	wire _peArray_37_taskOut_TVALID;
	wire [255:0] _peArray_37_taskOut_TDATA;
	wire _peArray_37_taskIn_TREADY;
	wire _peArray_36_closureIn_TREADY;
	wire _peArray_36_argOut_TVALID;
	wire [63:0] _peArray_36_argOut_TDATA;
	wire _peArray_36_taskOut_TVALID;
	wire [255:0] _peArray_36_taskOut_TDATA;
	wire _peArray_36_taskIn_TREADY;
	wire _peArray_35_closureIn_TREADY;
	wire _peArray_35_argOut_TVALID;
	wire [63:0] _peArray_35_argOut_TDATA;
	wire _peArray_35_taskOut_TVALID;
	wire [255:0] _peArray_35_taskOut_TDATA;
	wire _peArray_35_taskIn_TREADY;
	wire _peArray_34_closureIn_TREADY;
	wire _peArray_34_argOut_TVALID;
	wire [63:0] _peArray_34_argOut_TDATA;
	wire _peArray_34_taskOut_TVALID;
	wire [255:0] _peArray_34_taskOut_TDATA;
	wire _peArray_34_taskIn_TREADY;
	wire _peArray_33_closureIn_TREADY;
	wire _peArray_33_argOut_TVALID;
	wire [63:0] _peArray_33_argOut_TDATA;
	wire _peArray_33_taskOut_TVALID;
	wire [255:0] _peArray_33_taskOut_TDATA;
	wire _peArray_33_taskIn_TREADY;
	wire _peArray_32_closureIn_TREADY;
	wire _peArray_32_argOut_TVALID;
	wire [63:0] _peArray_32_argOut_TDATA;
	wire _peArray_32_taskOut_TVALID;
	wire [255:0] _peArray_32_taskOut_TDATA;
	wire _peArray_32_taskIn_TREADY;
	wire _peArray_31_closureIn_TREADY;
	wire _peArray_31_argOut_TVALID;
	wire [63:0] _peArray_31_argOut_TDATA;
	wire _peArray_31_taskOut_TVALID;
	wire [255:0] _peArray_31_taskOut_TDATA;
	wire _peArray_31_taskIn_TREADY;
	wire _peArray_30_closureIn_TREADY;
	wire _peArray_30_argOut_TVALID;
	wire [63:0] _peArray_30_argOut_TDATA;
	wire _peArray_30_taskOut_TVALID;
	wire [255:0] _peArray_30_taskOut_TDATA;
	wire _peArray_30_taskIn_TREADY;
	wire _peArray_29_closureIn_TREADY;
	wire _peArray_29_argOut_TVALID;
	wire [63:0] _peArray_29_argOut_TDATA;
	wire _peArray_29_taskOut_TVALID;
	wire [255:0] _peArray_29_taskOut_TDATA;
	wire _peArray_29_taskIn_TREADY;
	wire _peArray_28_closureIn_TREADY;
	wire _peArray_28_argOut_TVALID;
	wire [63:0] _peArray_28_argOut_TDATA;
	wire _peArray_28_taskOut_TVALID;
	wire [255:0] _peArray_28_taskOut_TDATA;
	wire _peArray_28_taskIn_TREADY;
	wire _peArray_27_closureIn_TREADY;
	wire _peArray_27_argOut_TVALID;
	wire [63:0] _peArray_27_argOut_TDATA;
	wire _peArray_27_taskOut_TVALID;
	wire [255:0] _peArray_27_taskOut_TDATA;
	wire _peArray_27_taskIn_TREADY;
	wire _peArray_26_closureIn_TREADY;
	wire _peArray_26_argOut_TVALID;
	wire [63:0] _peArray_26_argOut_TDATA;
	wire _peArray_26_taskOut_TVALID;
	wire [255:0] _peArray_26_taskOut_TDATA;
	wire _peArray_26_taskIn_TREADY;
	wire _peArray_25_closureIn_TREADY;
	wire _peArray_25_argOut_TVALID;
	wire [63:0] _peArray_25_argOut_TDATA;
	wire _peArray_25_taskOut_TVALID;
	wire [255:0] _peArray_25_taskOut_TDATA;
	wire _peArray_25_taskIn_TREADY;
	wire _peArray_24_closureIn_TREADY;
	wire _peArray_24_argOut_TVALID;
	wire [63:0] _peArray_24_argOut_TDATA;
	wire _peArray_24_taskOut_TVALID;
	wire [255:0] _peArray_24_taskOut_TDATA;
	wire _peArray_24_taskIn_TREADY;
	wire _peArray_23_closureIn_TREADY;
	wire _peArray_23_argOut_TVALID;
	wire [63:0] _peArray_23_argOut_TDATA;
	wire _peArray_23_taskOut_TVALID;
	wire [255:0] _peArray_23_taskOut_TDATA;
	wire _peArray_23_taskIn_TREADY;
	wire _peArray_22_closureIn_TREADY;
	wire _peArray_22_argOut_TVALID;
	wire [63:0] _peArray_22_argOut_TDATA;
	wire _peArray_22_taskOut_TVALID;
	wire [255:0] _peArray_22_taskOut_TDATA;
	wire _peArray_22_taskIn_TREADY;
	wire _peArray_21_closureIn_TREADY;
	wire _peArray_21_argOut_TVALID;
	wire [63:0] _peArray_21_argOut_TDATA;
	wire _peArray_21_taskOut_TVALID;
	wire [255:0] _peArray_21_taskOut_TDATA;
	wire _peArray_21_taskIn_TREADY;
	wire _peArray_20_closureIn_TREADY;
	wire _peArray_20_argOut_TVALID;
	wire [63:0] _peArray_20_argOut_TDATA;
	wire _peArray_20_taskOut_TVALID;
	wire [255:0] _peArray_20_taskOut_TDATA;
	wire _peArray_20_taskIn_TREADY;
	wire _peArray_19_closureIn_TREADY;
	wire _peArray_19_argOut_TVALID;
	wire [63:0] _peArray_19_argOut_TDATA;
	wire _peArray_19_taskOut_TVALID;
	wire [255:0] _peArray_19_taskOut_TDATA;
	wire _peArray_19_taskIn_TREADY;
	wire _peArray_18_closureIn_TREADY;
	wire _peArray_18_argOut_TVALID;
	wire [63:0] _peArray_18_argOut_TDATA;
	wire _peArray_18_taskOut_TVALID;
	wire [255:0] _peArray_18_taskOut_TDATA;
	wire _peArray_18_taskIn_TREADY;
	wire _peArray_17_closureIn_TREADY;
	wire _peArray_17_argOut_TVALID;
	wire [63:0] _peArray_17_argOut_TDATA;
	wire _peArray_17_taskOut_TVALID;
	wire [255:0] _peArray_17_taskOut_TDATA;
	wire _peArray_17_taskIn_TREADY;
	wire _peArray_16_closureIn_TREADY;
	wire _peArray_16_argOut_TVALID;
	wire [63:0] _peArray_16_argOut_TDATA;
	wire _peArray_16_taskOut_TVALID;
	wire [255:0] _peArray_16_taskOut_TDATA;
	wire _peArray_16_taskIn_TREADY;
	wire _peArray_15_closureIn_TREADY;
	wire _peArray_15_argOut_TVALID;
	wire [63:0] _peArray_15_argOut_TDATA;
	wire _peArray_15_taskOut_TVALID;
	wire [255:0] _peArray_15_taskOut_TDATA;
	wire _peArray_15_taskIn_TREADY;
	wire _peArray_14_closureIn_TREADY;
	wire _peArray_14_argOut_TVALID;
	wire [63:0] _peArray_14_argOut_TDATA;
	wire _peArray_14_taskOut_TVALID;
	wire [255:0] _peArray_14_taskOut_TDATA;
	wire _peArray_14_taskIn_TREADY;
	wire _peArray_13_closureIn_TREADY;
	wire _peArray_13_argOut_TVALID;
	wire [63:0] _peArray_13_argOut_TDATA;
	wire _peArray_13_taskOut_TVALID;
	wire [255:0] _peArray_13_taskOut_TDATA;
	wire _peArray_13_taskIn_TREADY;
	wire _peArray_12_closureIn_TREADY;
	wire _peArray_12_argOut_TVALID;
	wire [63:0] _peArray_12_argOut_TDATA;
	wire _peArray_12_taskOut_TVALID;
	wire [255:0] _peArray_12_taskOut_TDATA;
	wire _peArray_12_taskIn_TREADY;
	wire _peArray_11_closureIn_TREADY;
	wire _peArray_11_argOut_TVALID;
	wire [63:0] _peArray_11_argOut_TDATA;
	wire _peArray_11_taskOut_TVALID;
	wire [255:0] _peArray_11_taskOut_TDATA;
	wire _peArray_11_taskIn_TREADY;
	wire _peArray_10_closureIn_TREADY;
	wire _peArray_10_argOut_TVALID;
	wire [63:0] _peArray_10_argOut_TDATA;
	wire _peArray_10_taskOut_TVALID;
	wire [255:0] _peArray_10_taskOut_TDATA;
	wire _peArray_10_taskIn_TREADY;
	wire _peArray_9_closureIn_TREADY;
	wire _peArray_9_argOut_TVALID;
	wire [63:0] _peArray_9_argOut_TDATA;
	wire _peArray_9_taskOut_TVALID;
	wire [255:0] _peArray_9_taskOut_TDATA;
	wire _peArray_9_taskIn_TREADY;
	wire _peArray_8_closureIn_TREADY;
	wire _peArray_8_argOut_TVALID;
	wire [63:0] _peArray_8_argOut_TDATA;
	wire _peArray_8_taskOut_TVALID;
	wire [255:0] _peArray_8_taskOut_TDATA;
	wire _peArray_8_taskIn_TREADY;
	wire _peArray_7_closureIn_TREADY;
	wire _peArray_7_argOut_TVALID;
	wire [63:0] _peArray_7_argOut_TDATA;
	wire _peArray_7_taskOut_TVALID;
	wire [255:0] _peArray_7_taskOut_TDATA;
	wire _peArray_7_taskIn_TREADY;
	wire _peArray_6_closureIn_TREADY;
	wire _peArray_6_argOut_TVALID;
	wire [63:0] _peArray_6_argOut_TDATA;
	wire _peArray_6_taskOut_TVALID;
	wire [255:0] _peArray_6_taskOut_TDATA;
	wire _peArray_6_taskIn_TREADY;
	wire _peArray_5_closureIn_TREADY;
	wire _peArray_5_argOut_TVALID;
	wire [63:0] _peArray_5_argOut_TDATA;
	wire _peArray_5_taskOut_TVALID;
	wire [255:0] _peArray_5_taskOut_TDATA;
	wire _peArray_5_taskIn_TREADY;
	wire _peArray_4_closureIn_TREADY;
	wire _peArray_4_argOut_TVALID;
	wire [63:0] _peArray_4_argOut_TDATA;
	wire _peArray_4_taskOut_TVALID;
	wire [255:0] _peArray_4_taskOut_TDATA;
	wire _peArray_4_taskIn_TREADY;
	wire _peArray_3_closureIn_TREADY;
	wire _peArray_3_argOut_TVALID;
	wire [63:0] _peArray_3_argOut_TDATA;
	wire _peArray_3_taskOut_TVALID;
	wire [255:0] _peArray_3_taskOut_TDATA;
	wire _peArray_3_taskIn_TREADY;
	wire _peArray_2_closureIn_TREADY;
	wire _peArray_2_argOut_TVALID;
	wire [63:0] _peArray_2_argOut_TDATA;
	wire _peArray_2_taskOut_TVALID;
	wire [255:0] _peArray_2_taskOut_TDATA;
	wire _peArray_2_taskIn_TREADY;
	wire _peArray_1_closureIn_TREADY;
	wire _peArray_1_argOut_TVALID;
	wire [63:0] _peArray_1_argOut_TDATA;
	wire _peArray_1_taskOut_TVALID;
	wire [255:0] _peArray_1_taskOut_TDATA;
	wire _peArray_1_taskIn_TREADY;
	wire _peArray_0_closureIn_TREADY;
	wire _peArray_0_argOut_TVALID;
	wire [63:0] _peArray_0_argOut_TDATA;
	wire _peArray_0_taskOut_TVALID;
	wire [255:0] _peArray_0_taskOut_TDATA;
	wire _peArray_0_taskIn_TREADY;
	wire _demux_m_axil_0_ar_valid;
	wire [11:0] _demux_m_axil_0_ar_bits_addr;
	wire [2:0] _demux_m_axil_0_ar_bits_prot;
	wire _demux_m_axil_0_r_ready;
	wire _demux_m_axil_0_aw_valid;
	wire [11:0] _demux_m_axil_0_aw_bits_addr;
	wire [2:0] _demux_m_axil_0_aw_bits_prot;
	wire _demux_m_axil_0_w_valid;
	wire [63:0] _demux_m_axil_0_w_bits_data;
	wire [7:0] _demux_m_axil_0_w_bits_strb;
	wire _demux_m_axil_0_b_ready;
	wire _demux_m_axil_1_ar_valid;
	wire [11:0] _demux_m_axil_1_ar_bits_addr;
	wire [2:0] _demux_m_axil_1_ar_bits_prot;
	wire _demux_m_axil_1_r_ready;
	wire _demux_m_axil_1_aw_valid;
	wire [11:0] _demux_m_axil_1_aw_bits_addr;
	wire [2:0] _demux_m_axil_1_aw_bits_prot;
	wire _demux_m_axil_1_w_valid;
	wire [63:0] _demux_m_axil_1_w_bits_data;
	wire [7:0] _demux_m_axil_1_w_bits_strb;
	wire _demux_m_axil_1_b_ready;
	wire _demux_m_axil_2_ar_valid;
	wire [11:0] _demux_m_axil_2_ar_bits_addr;
	wire [2:0] _demux_m_axil_2_ar_bits_prot;
	wire _demux_m_axil_2_r_ready;
	wire _demux_m_axil_2_aw_valid;
	wire [11:0] _demux_m_axil_2_aw_bits_addr;
	wire [2:0] _demux_m_axil_2_aw_bits_prot;
	wire _demux_m_axil_2_w_valid;
	wire [63:0] _demux_m_axil_2_w_bits_data;
	wire [7:0] _demux_m_axil_2_w_bits_strb;
	wire _demux_m_axil_2_b_ready;
	wire _demux_m_axil_3_ar_valid;
	wire [11:0] _demux_m_axil_3_ar_bits_addr;
	wire [2:0] _demux_m_axil_3_ar_bits_prot;
	wire _demux_m_axil_3_r_ready;
	wire _demux_m_axil_3_aw_valid;
	wire [11:0] _demux_m_axil_3_aw_bits_addr;
	wire [2:0] _demux_m_axil_3_aw_bits_prot;
	wire _demux_m_axil_3_w_valid;
	wire [63:0] _demux_m_axil_3_w_bits_data;
	wire [7:0] _demux_m_axil_3_w_bits_strb;
	wire _demux_m_axil_3_b_ready;
	wire _demux_m_axil_4_ar_valid;
	wire [11:0] _demux_m_axil_4_ar_bits_addr;
	wire [2:0] _demux_m_axil_4_ar_bits_prot;
	wire _demux_m_axil_4_r_ready;
	wire _demux_m_axil_4_aw_valid;
	wire [11:0] _demux_m_axil_4_aw_bits_addr;
	wire [2:0] _demux_m_axil_4_aw_bits_prot;
	wire _demux_m_axil_4_w_valid;
	wire [63:0] _demux_m_axil_4_w_bits_data;
	wire [7:0] _demux_m_axil_4_w_bits_strb;
	wire _demux_m_axil_4_b_ready;
	wire _demux_m_axil_5_ar_valid;
	wire [11:0] _demux_m_axil_5_ar_bits_addr;
	wire [2:0] _demux_m_axil_5_ar_bits_prot;
	wire _demux_m_axil_5_r_ready;
	wire _demux_m_axil_5_aw_valid;
	wire [11:0] _demux_m_axil_5_aw_bits_addr;
	wire [2:0] _demux_m_axil_5_aw_bits_prot;
	wire _demux_m_axil_5_w_valid;
	wire [63:0] _demux_m_axil_5_w_bits_data;
	wire [7:0] _demux_m_axil_5_w_bits_strb;
	wire _demux_m_axil_5_b_ready;
	axi4LiteDemux demux(
		.clock(clock),
		.reset(reset),
		.s_axil_ar_ready(s_axil_mgmt_hardcilk_ARREADY),
		.s_axil_ar_valid(s_axil_mgmt_hardcilk_ARVALID),
		.s_axil_ar_bits_addr(s_axil_mgmt_hardcilk_ARADDR),
		.s_axil_ar_bits_prot(s_axil_mgmt_hardcilk_ARPROT),
		.s_axil_r_ready(s_axil_mgmt_hardcilk_RREADY),
		.s_axil_r_valid(s_axil_mgmt_hardcilk_RVALID),
		.s_axil_r_bits_data(s_axil_mgmt_hardcilk_RDATA),
		.s_axil_r_bits_resp(s_axil_mgmt_hardcilk_RRESP),
		.s_axil_aw_ready(s_axil_mgmt_hardcilk_AWREADY),
		.s_axil_aw_valid(s_axil_mgmt_hardcilk_AWVALID),
		.s_axil_aw_bits_addr(s_axil_mgmt_hardcilk_AWADDR),
		.s_axil_aw_bits_prot(s_axil_mgmt_hardcilk_AWPROT),
		.s_axil_w_ready(s_axil_mgmt_hardcilk_WREADY),
		.s_axil_w_valid(s_axil_mgmt_hardcilk_WVALID),
		.s_axil_w_bits_data(s_axil_mgmt_hardcilk_WDATA),
		.s_axil_w_bits_strb(s_axil_mgmt_hardcilk_WSTRB),
		.s_axil_b_ready(s_axil_mgmt_hardcilk_BREADY),
		.s_axil_b_valid(s_axil_mgmt_hardcilk_BVALID),
		.s_axil_b_bits_resp(s_axil_mgmt_hardcilk_BRESP),
		.m_axil_0_ar_ready(_Scheduler_io_internal_axi_mgmt_vss_0_ar_ready),
		.m_axil_0_ar_valid(_demux_m_axil_0_ar_valid),
		.m_axil_0_ar_bits_addr(_demux_m_axil_0_ar_bits_addr),
		.m_axil_0_ar_bits_prot(_demux_m_axil_0_ar_bits_prot),
		.m_axil_0_r_ready(_demux_m_axil_0_r_ready),
		.m_axil_0_r_valid(_Scheduler_io_internal_axi_mgmt_vss_0_r_valid),
		.m_axil_0_r_bits_data(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_data),
		.m_axil_0_r_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.m_axil_0_aw_ready(_Scheduler_io_internal_axi_mgmt_vss_0_aw_ready),
		.m_axil_0_aw_valid(_demux_m_axil_0_aw_valid),
		.m_axil_0_aw_bits_addr(_demux_m_axil_0_aw_bits_addr),
		.m_axil_0_aw_bits_prot(_demux_m_axil_0_aw_bits_prot),
		.m_axil_0_w_ready(_Scheduler_io_internal_axi_mgmt_vss_0_w_ready),
		.m_axil_0_w_valid(_demux_m_axil_0_w_valid),
		.m_axil_0_w_bits_data(_demux_m_axil_0_w_bits_data),
		.m_axil_0_w_bits_strb(_demux_m_axil_0_w_bits_strb),
		.m_axil_0_b_ready(_demux_m_axil_0_b_ready),
		.m_axil_0_b_valid(_Scheduler_io_internal_axi_mgmt_vss_0_b_valid),
		.m_axil_0_b_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.m_axil_1_ar_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_ar_ready),
		.m_axil_1_ar_valid(_demux_m_axil_1_ar_valid),
		.m_axil_1_ar_bits_addr(_demux_m_axil_1_ar_bits_addr),
		.m_axil_1_ar_bits_prot(_demux_m_axil_1_ar_bits_prot),
		.m_axil_1_r_ready(_demux_m_axil_1_r_ready),
		.m_axil_1_r_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_valid),
		.m_axil_1_r_bits_data(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_data),
		.m_axil_1_r_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.m_axil_1_aw_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_aw_ready),
		.m_axil_1_aw_valid(_demux_m_axil_1_aw_valid),
		.m_axil_1_aw_bits_addr(_demux_m_axil_1_aw_bits_addr),
		.m_axil_1_aw_bits_prot(_demux_m_axil_1_aw_bits_prot),
		.m_axil_1_w_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_w_ready),
		.m_axil_1_w_valid(_demux_m_axil_1_w_valid),
		.m_axil_1_w_bits_data(_demux_m_axil_1_w_bits_data),
		.m_axil_1_w_bits_strb(_demux_m_axil_1_w_bits_strb),
		.m_axil_1_b_ready(_demux_m_axil_1_b_ready),
		.m_axil_1_b_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_valid),
		.m_axil_1_b_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.m_axil_2_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_0_ar_ready),
		.m_axil_2_ar_valid(_demux_m_axil_2_ar_valid),
		.m_axil_2_ar_bits_addr(_demux_m_axil_2_ar_bits_addr),
		.m_axil_2_ar_bits_prot(_demux_m_axil_2_ar_bits_prot),
		.m_axil_2_r_ready(_demux_m_axil_2_r_ready),
		.m_axil_2_r_valid(_Allocator_io_internal_axi_mgmt_vcas_0_r_valid),
		.m_axil_2_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_data),
		.m_axil_2_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_resp),
		.m_axil_2_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_0_aw_ready),
		.m_axil_2_aw_valid(_demux_m_axil_2_aw_valid),
		.m_axil_2_aw_bits_addr(_demux_m_axil_2_aw_bits_addr),
		.m_axil_2_aw_bits_prot(_demux_m_axil_2_aw_bits_prot),
		.m_axil_2_w_ready(_Allocator_io_internal_axi_mgmt_vcas_0_w_ready),
		.m_axil_2_w_valid(_demux_m_axil_2_w_valid),
		.m_axil_2_w_bits_data(_demux_m_axil_2_w_bits_data),
		.m_axil_2_w_bits_strb(_demux_m_axil_2_w_bits_strb),
		.m_axil_2_b_ready(_demux_m_axil_2_b_ready),
		.m_axil_2_b_valid(_Allocator_io_internal_axi_mgmt_vcas_0_b_valid),
		.m_axil_2_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_b_bits_resp),
		.m_axil_3_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_1_ar_ready),
		.m_axil_3_ar_valid(_demux_m_axil_3_ar_valid),
		.m_axil_3_ar_bits_addr(_demux_m_axil_3_ar_bits_addr),
		.m_axil_3_ar_bits_prot(_demux_m_axil_3_ar_bits_prot),
		.m_axil_3_r_ready(_demux_m_axil_3_r_ready),
		.m_axil_3_r_valid(_Allocator_io_internal_axi_mgmt_vcas_1_r_valid),
		.m_axil_3_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_data),
		.m_axil_3_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_resp),
		.m_axil_3_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_1_aw_ready),
		.m_axil_3_aw_valid(_demux_m_axil_3_aw_valid),
		.m_axil_3_aw_bits_addr(_demux_m_axil_3_aw_bits_addr),
		.m_axil_3_aw_bits_prot(_demux_m_axil_3_aw_bits_prot),
		.m_axil_3_w_ready(_Allocator_io_internal_axi_mgmt_vcas_1_w_ready),
		.m_axil_3_w_valid(_demux_m_axil_3_w_valid),
		.m_axil_3_w_bits_data(_demux_m_axil_3_w_bits_data),
		.m_axil_3_w_bits_strb(_demux_m_axil_3_w_bits_strb),
		.m_axil_3_b_ready(_demux_m_axil_3_b_ready),
		.m_axil_3_b_valid(_Allocator_io_internal_axi_mgmt_vcas_1_b_valid),
		.m_axil_3_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_b_bits_resp),
		.m_axil_4_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_2_ar_ready),
		.m_axil_4_ar_valid(_demux_m_axil_4_ar_valid),
		.m_axil_4_ar_bits_addr(_demux_m_axil_4_ar_bits_addr),
		.m_axil_4_ar_bits_prot(_demux_m_axil_4_ar_bits_prot),
		.m_axil_4_r_ready(_demux_m_axil_4_r_ready),
		.m_axil_4_r_valid(_Allocator_io_internal_axi_mgmt_vcas_2_r_valid),
		.m_axil_4_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_data),
		.m_axil_4_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_resp),
		.m_axil_4_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_2_aw_ready),
		.m_axil_4_aw_valid(_demux_m_axil_4_aw_valid),
		.m_axil_4_aw_bits_addr(_demux_m_axil_4_aw_bits_addr),
		.m_axil_4_aw_bits_prot(_demux_m_axil_4_aw_bits_prot),
		.m_axil_4_w_ready(_Allocator_io_internal_axi_mgmt_vcas_2_w_ready),
		.m_axil_4_w_valid(_demux_m_axil_4_w_valid),
		.m_axil_4_w_bits_data(_demux_m_axil_4_w_bits_data),
		.m_axil_4_w_bits_strb(_demux_m_axil_4_w_bits_strb),
		.m_axil_4_b_ready(_demux_m_axil_4_b_ready),
		.m_axil_4_b_valid(_Allocator_io_internal_axi_mgmt_vcas_2_b_valid),
		.m_axil_4_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_b_bits_resp),
		.m_axil_5_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_3_ar_ready),
		.m_axil_5_ar_valid(_demux_m_axil_5_ar_valid),
		.m_axil_5_ar_bits_addr(_demux_m_axil_5_ar_bits_addr),
		.m_axil_5_ar_bits_prot(_demux_m_axil_5_ar_bits_prot),
		.m_axil_5_r_ready(_demux_m_axil_5_r_ready),
		.m_axil_5_r_valid(_Allocator_io_internal_axi_mgmt_vcas_3_r_valid),
		.m_axil_5_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_data),
		.m_axil_5_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_resp),
		.m_axil_5_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_3_aw_ready),
		.m_axil_5_aw_valid(_demux_m_axil_5_aw_valid),
		.m_axil_5_aw_bits_addr(_demux_m_axil_5_aw_bits_addr),
		.m_axil_5_aw_bits_prot(_demux_m_axil_5_aw_bits_prot),
		.m_axil_5_w_ready(_Allocator_io_internal_axi_mgmt_vcas_3_w_ready),
		.m_axil_5_w_valid(_demux_m_axil_5_w_valid),
		.m_axil_5_w_bits_data(_demux_m_axil_5_w_bits_data),
		.m_axil_5_w_bits_strb(_demux_m_axil_5_w_bits_strb),
		.m_axil_5_b_ready(_demux_m_axil_5_b_ready),
		.m_axil_5_b_valid(_Allocator_io_internal_axi_mgmt_vcas_3_b_valid),
		.m_axil_5_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_b_bits_resp)
	);
	qsort peArray_0(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_0_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_0_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_0_TREADY),
		.argOut_TVALID(_peArray_0_argOut_TVALID),
		.argOut_TDATA(_peArray_0_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_0_TREADY),
		.taskOut_TVALID(_peArray_0_taskOut_TVALID),
		.taskOut_TDATA(_peArray_0_taskOut_TDATA),
		.taskIn_TREADY(_peArray_0_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_0_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_0_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_0_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_0_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_0_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_0_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_0_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_0_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_0_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_0_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_0_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_0_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_0_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_0_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_0_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_0_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_0_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_0_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_0_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_0_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_0_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_0_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_0_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_0_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_0_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_0_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_0_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_0_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_0_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_0_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_0_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_0_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_0_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_0_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_0_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_0_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_0_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_0_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_0_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_0_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_0_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_0_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_0_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_0_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_0_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_0_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_0_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_0_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_0_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_0_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_0_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_0_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_0_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_0_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_0_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_0_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_0_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_0_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_0_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_0_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_0_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_0_m_axi_gmem_BUSER)
	);
	qsort peArray_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_1_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_1_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_1_TREADY),
		.argOut_TVALID(_peArray_1_argOut_TVALID),
		.argOut_TDATA(_peArray_1_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_1_TREADY),
		.taskOut_TVALID(_peArray_1_taskOut_TVALID),
		.taskOut_TDATA(_peArray_1_taskOut_TDATA),
		.taskIn_TREADY(_peArray_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_1_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_1_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_1_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_1_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_1_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_1_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_1_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_1_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_1_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_1_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_1_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_1_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_1_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_1_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_1_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_1_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_1_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_1_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_1_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_1_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_1_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_1_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_1_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_1_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_1_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_1_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_1_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_1_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_1_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_1_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_1_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_1_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_1_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_1_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_1_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_1_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_1_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_1_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_1_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_1_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_1_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_1_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_1_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_1_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_1_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_1_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_1_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_1_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_1_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_1_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_1_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_1_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_1_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_1_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_1_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_1_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_1_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_1_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_1_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_1_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_1_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_1_m_axi_gmem_BUSER)
	);
	qsort peArray_2(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_2_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_2_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_2_TREADY),
		.argOut_TVALID(_peArray_2_argOut_TVALID),
		.argOut_TDATA(_peArray_2_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_2_TREADY),
		.taskOut_TVALID(_peArray_2_taskOut_TVALID),
		.taskOut_TDATA(_peArray_2_taskOut_TDATA),
		.taskIn_TREADY(_peArray_2_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_2_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_2_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_2_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_2_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_2_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_2_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_2_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_2_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_2_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_2_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_2_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_2_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_2_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_2_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_2_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_2_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_2_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_2_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_2_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_2_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_2_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_2_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_2_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_2_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_2_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_2_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_2_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_2_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_2_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_2_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_2_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_2_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_2_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_2_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_2_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_2_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_2_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_2_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_2_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_2_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_2_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_2_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_2_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_2_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_2_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_2_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_2_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_2_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_2_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_2_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_2_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_2_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_2_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_2_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_2_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_2_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_2_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_2_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_2_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_2_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_2_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_2_m_axi_gmem_BUSER)
	);
	qsort peArray_3(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_3_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_3_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_3_TREADY),
		.argOut_TVALID(_peArray_3_argOut_TVALID),
		.argOut_TDATA(_peArray_3_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_3_TREADY),
		.taskOut_TVALID(_peArray_3_taskOut_TVALID),
		.taskOut_TDATA(_peArray_3_taskOut_TDATA),
		.taskIn_TREADY(_peArray_3_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_3_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_3_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_3_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_3_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_3_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_3_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_3_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_3_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_3_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_3_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_3_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_3_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_3_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_3_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_3_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_3_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_3_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_3_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_3_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_3_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_3_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_3_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_3_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_3_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_3_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_3_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_3_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_3_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_3_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_3_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_3_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_3_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_3_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_3_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_3_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_3_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_3_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_3_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_3_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_3_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_3_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_3_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_3_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_3_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_3_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_3_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_3_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_3_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_3_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_3_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_3_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_3_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_3_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_3_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_3_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_3_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_3_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_3_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_3_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_3_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_3_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_3_m_axi_gmem_BUSER)
	);
	qsort peArray_4(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_4_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_4_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_4_TREADY),
		.argOut_TVALID(_peArray_4_argOut_TVALID),
		.argOut_TDATA(_peArray_4_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_4_TREADY),
		.taskOut_TVALID(_peArray_4_taskOut_TVALID),
		.taskOut_TDATA(_peArray_4_taskOut_TDATA),
		.taskIn_TREADY(_peArray_4_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_4_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_4_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_4_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_4_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_4_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_4_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_4_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_4_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_4_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_4_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_4_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_4_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_4_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_4_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_4_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_4_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_4_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_4_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_4_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_4_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_4_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_4_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_4_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_4_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_4_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_4_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_4_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_4_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_4_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_4_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_4_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_4_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_4_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_4_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_4_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_4_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_4_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_4_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_4_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_4_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_4_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_4_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_4_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_4_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_4_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_4_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_4_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_4_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_4_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_4_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_4_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_4_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_4_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_4_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_4_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_4_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_4_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_4_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_4_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_4_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_4_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_4_m_axi_gmem_BUSER)
	);
	qsort peArray_5(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_5_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_5_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_5_TREADY),
		.argOut_TVALID(_peArray_5_argOut_TVALID),
		.argOut_TDATA(_peArray_5_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_5_TREADY),
		.taskOut_TVALID(_peArray_5_taskOut_TVALID),
		.taskOut_TDATA(_peArray_5_taskOut_TDATA),
		.taskIn_TREADY(_peArray_5_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_5_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_5_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_5_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_5_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_5_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_5_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_5_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_5_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_5_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_5_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_5_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_5_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_5_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_5_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_5_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_5_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_5_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_5_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_5_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_5_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_5_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_5_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_5_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_5_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_5_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_5_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_5_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_5_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_5_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_5_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_5_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_5_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_5_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_5_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_5_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_5_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_5_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_5_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_5_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_5_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_5_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_5_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_5_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_5_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_5_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_5_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_5_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_5_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_5_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_5_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_5_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_5_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_5_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_5_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_5_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_5_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_5_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_5_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_5_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_5_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_5_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_5_m_axi_gmem_BUSER)
	);
	qsort peArray_6(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_6_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_6_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_6_TREADY),
		.argOut_TVALID(_peArray_6_argOut_TVALID),
		.argOut_TDATA(_peArray_6_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_6_TREADY),
		.taskOut_TVALID(_peArray_6_taskOut_TVALID),
		.taskOut_TDATA(_peArray_6_taskOut_TDATA),
		.taskIn_TREADY(_peArray_6_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_6_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_6_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_6_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_6_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_6_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_6_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_6_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_6_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_6_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_6_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_6_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_6_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_6_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_6_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_6_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_6_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_6_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_6_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_6_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_6_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_6_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_6_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_6_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_6_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_6_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_6_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_6_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_6_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_6_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_6_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_6_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_6_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_6_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_6_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_6_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_6_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_6_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_6_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_6_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_6_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_6_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_6_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_6_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_6_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_6_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_6_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_6_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_6_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_6_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_6_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_6_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_6_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_6_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_6_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_6_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_6_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_6_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_6_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_6_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_6_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_6_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_6_m_axi_gmem_BUSER)
	);
	qsort peArray_7(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_7_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_7_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_7_TREADY),
		.argOut_TVALID(_peArray_7_argOut_TVALID),
		.argOut_TDATA(_peArray_7_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_7_TREADY),
		.taskOut_TVALID(_peArray_7_taskOut_TVALID),
		.taskOut_TDATA(_peArray_7_taskOut_TDATA),
		.taskIn_TREADY(_peArray_7_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_7_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_7_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_7_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_7_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_7_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_7_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_7_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_7_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_7_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_7_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_7_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_7_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_7_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_7_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_7_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_7_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_7_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_7_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_7_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_7_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_7_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_7_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_7_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_7_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_7_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_7_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_7_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_7_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_7_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_7_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_7_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_7_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_7_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_7_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_7_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_7_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_7_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_7_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_7_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_7_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_7_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_7_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_7_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_7_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_7_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_7_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_7_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_7_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_7_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_7_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_7_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_7_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_7_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_7_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_7_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_7_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_7_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_7_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_7_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_7_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_7_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_7_m_axi_gmem_BUSER)
	);
	qsort peArray_8(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_8_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_8_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_8_TREADY),
		.argOut_TVALID(_peArray_8_argOut_TVALID),
		.argOut_TDATA(_peArray_8_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_8_TREADY),
		.taskOut_TVALID(_peArray_8_taskOut_TVALID),
		.taskOut_TDATA(_peArray_8_taskOut_TDATA),
		.taskIn_TREADY(_peArray_8_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_8_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_8_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_8_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_8_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_8_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_8_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_8_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_8_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_8_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_8_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_8_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_8_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_8_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_8_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_8_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_8_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_8_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_8_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_8_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_8_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_8_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_8_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_8_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_8_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_8_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_8_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_8_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_8_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_8_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_8_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_8_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_8_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_8_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_8_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_8_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_8_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_8_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_8_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_8_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_8_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_8_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_8_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_8_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_8_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_8_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_8_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_8_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_8_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_8_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_8_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_8_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_8_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_8_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_8_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_8_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_8_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_8_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_8_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_8_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_8_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_8_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_8_m_axi_gmem_BUSER)
	);
	qsort peArray_9(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_9_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_9_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_9_TREADY),
		.argOut_TVALID(_peArray_9_argOut_TVALID),
		.argOut_TDATA(_peArray_9_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_9_TREADY),
		.taskOut_TVALID(_peArray_9_taskOut_TVALID),
		.taskOut_TDATA(_peArray_9_taskOut_TDATA),
		.taskIn_TREADY(_peArray_9_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_9_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_9_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_9_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_9_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_9_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_9_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_9_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_9_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_9_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_9_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_9_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_9_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_9_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_9_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_9_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_9_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_9_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_9_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_9_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_9_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_9_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_9_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_9_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_9_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_9_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_9_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_9_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_9_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_9_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_9_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_9_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_9_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_9_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_9_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_9_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_9_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_9_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_9_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_9_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_9_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_9_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_9_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_9_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_9_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_9_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_9_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_9_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_9_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_9_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_9_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_9_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_9_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_9_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_9_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_9_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_9_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_9_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_9_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_9_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_9_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_9_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_9_m_axi_gmem_BUSER)
	);
	qsort peArray_10(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_10_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_10_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_10_TREADY),
		.argOut_TVALID(_peArray_10_argOut_TVALID),
		.argOut_TDATA(_peArray_10_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_10_TREADY),
		.taskOut_TVALID(_peArray_10_taskOut_TVALID),
		.taskOut_TDATA(_peArray_10_taskOut_TDATA),
		.taskIn_TREADY(_peArray_10_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_10_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_10_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_10_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_10_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_10_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_10_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_10_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_10_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_10_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_10_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_10_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_10_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_10_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_10_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_10_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_10_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_10_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_10_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_10_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_10_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_10_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_10_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_10_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_10_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_10_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_10_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_10_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_10_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_10_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_10_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_10_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_10_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_10_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_10_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_10_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_10_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_10_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_10_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_10_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_10_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_10_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_10_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_10_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_10_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_10_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_10_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_10_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_10_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_10_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_10_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_10_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_10_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_10_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_10_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_10_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_10_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_10_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_10_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_10_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_10_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_10_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_10_m_axi_gmem_BUSER)
	);
	qsort peArray_11(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_11_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_11_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_11_TREADY),
		.argOut_TVALID(_peArray_11_argOut_TVALID),
		.argOut_TDATA(_peArray_11_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_11_TREADY),
		.taskOut_TVALID(_peArray_11_taskOut_TVALID),
		.taskOut_TDATA(_peArray_11_taskOut_TDATA),
		.taskIn_TREADY(_peArray_11_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_11_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_11_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_11_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_11_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_11_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_11_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_11_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_11_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_11_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_11_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_11_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_11_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_11_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_11_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_11_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_11_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_11_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_11_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_11_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_11_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_11_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_11_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_11_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_11_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_11_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_11_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_11_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_11_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_11_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_11_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_11_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_11_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_11_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_11_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_11_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_11_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_11_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_11_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_11_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_11_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_11_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_11_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_11_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_11_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_11_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_11_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_11_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_11_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_11_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_11_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_11_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_11_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_11_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_11_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_11_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_11_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_11_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_11_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_11_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_11_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_11_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_11_m_axi_gmem_BUSER)
	);
	qsort peArray_12(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_12_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_12_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_12_TREADY),
		.argOut_TVALID(_peArray_12_argOut_TVALID),
		.argOut_TDATA(_peArray_12_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_12_TREADY),
		.taskOut_TVALID(_peArray_12_taskOut_TVALID),
		.taskOut_TDATA(_peArray_12_taskOut_TDATA),
		.taskIn_TREADY(_peArray_12_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_12_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_12_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_12_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_12_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_12_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_12_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_12_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_12_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_12_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_12_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_12_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_12_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_12_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_12_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_12_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_12_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_12_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_12_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_12_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_12_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_12_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_12_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_12_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_12_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_12_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_12_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_12_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_12_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_12_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_12_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_12_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_12_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_12_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_12_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_12_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_12_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_12_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_12_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_12_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_12_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_12_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_12_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_12_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_12_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_12_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_12_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_12_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_12_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_12_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_12_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_12_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_12_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_12_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_12_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_12_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_12_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_12_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_12_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_12_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_12_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_12_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_12_m_axi_gmem_BUSER)
	);
	qsort peArray_13(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_13_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_13_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_13_TREADY),
		.argOut_TVALID(_peArray_13_argOut_TVALID),
		.argOut_TDATA(_peArray_13_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_13_TREADY),
		.taskOut_TVALID(_peArray_13_taskOut_TVALID),
		.taskOut_TDATA(_peArray_13_taskOut_TDATA),
		.taskIn_TREADY(_peArray_13_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_13_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_13_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_13_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_13_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_13_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_13_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_13_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_13_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_13_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_13_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_13_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_13_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_13_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_13_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_13_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_13_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_13_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_13_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_13_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_13_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_13_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_13_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_13_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_13_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_13_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_13_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_13_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_13_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_13_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_13_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_13_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_13_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_13_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_13_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_13_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_13_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_13_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_13_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_13_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_13_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_13_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_13_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_13_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_13_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_13_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_13_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_13_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_13_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_13_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_13_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_13_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_13_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_13_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_13_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_13_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_13_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_13_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_13_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_13_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_13_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_13_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_13_m_axi_gmem_BUSER)
	);
	qsort peArray_14(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_14_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_14_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_14_TREADY),
		.argOut_TVALID(_peArray_14_argOut_TVALID),
		.argOut_TDATA(_peArray_14_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_14_TREADY),
		.taskOut_TVALID(_peArray_14_taskOut_TVALID),
		.taskOut_TDATA(_peArray_14_taskOut_TDATA),
		.taskIn_TREADY(_peArray_14_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_14_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_14_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_14_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_14_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_14_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_14_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_14_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_14_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_14_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_14_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_14_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_14_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_14_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_14_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_14_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_14_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_14_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_14_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_14_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_14_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_14_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_14_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_14_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_14_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_14_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_14_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_14_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_14_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_14_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_14_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_14_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_14_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_14_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_14_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_14_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_14_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_14_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_14_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_14_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_14_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_14_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_14_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_14_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_14_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_14_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_14_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_14_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_14_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_14_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_14_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_14_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_14_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_14_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_14_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_14_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_14_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_14_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_14_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_14_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_14_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_14_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_14_m_axi_gmem_BUSER)
	);
	qsort peArray_15(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_15_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_15_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_15_TREADY),
		.argOut_TVALID(_peArray_15_argOut_TVALID),
		.argOut_TDATA(_peArray_15_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_15_TREADY),
		.taskOut_TVALID(_peArray_15_taskOut_TVALID),
		.taskOut_TDATA(_peArray_15_taskOut_TDATA),
		.taskIn_TREADY(_peArray_15_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_15_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_15_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_15_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_15_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_15_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_15_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_15_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_15_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_15_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_15_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_15_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_15_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_15_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_15_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_15_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_15_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_15_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_15_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_15_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_15_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_15_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_15_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_15_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_15_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_15_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_15_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_15_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_15_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_15_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_15_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_15_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_15_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_15_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_15_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_15_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_15_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_15_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_15_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_15_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_15_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_15_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_15_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_15_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_15_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_15_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_15_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_15_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_15_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_15_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_15_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_15_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_15_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_15_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_15_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_15_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_15_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_15_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_15_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_15_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_15_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_15_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_15_m_axi_gmem_BUSER)
	);
	qsort peArray_16(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_16_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_16_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_16_TREADY),
		.argOut_TVALID(_peArray_16_argOut_TVALID),
		.argOut_TDATA(_peArray_16_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_16_TREADY),
		.taskOut_TVALID(_peArray_16_taskOut_TVALID),
		.taskOut_TDATA(_peArray_16_taskOut_TDATA),
		.taskIn_TREADY(_peArray_16_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_16_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_16_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_16_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_16_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_16_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_16_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_16_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_16_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_16_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_16_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_16_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_16_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_16_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_16_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_16_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_16_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_16_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_16_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_16_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_16_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_16_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_16_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_16_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_16_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_16_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_16_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_16_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_16_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_16_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_16_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_16_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_16_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_16_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_16_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_16_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_16_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_16_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_16_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_16_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_16_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_16_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_16_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_16_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_16_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_16_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_16_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_16_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_16_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_16_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_16_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_16_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_16_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_16_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_16_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_16_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_16_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_16_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_16_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_16_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_16_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_16_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_16_m_axi_gmem_BUSER)
	);
	qsort peArray_17(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_17_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_17_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_17_TREADY),
		.argOut_TVALID(_peArray_17_argOut_TVALID),
		.argOut_TDATA(_peArray_17_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_17_TREADY),
		.taskOut_TVALID(_peArray_17_taskOut_TVALID),
		.taskOut_TDATA(_peArray_17_taskOut_TDATA),
		.taskIn_TREADY(_peArray_17_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_17_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_17_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_17_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_17_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_17_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_17_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_17_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_17_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_17_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_17_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_17_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_17_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_17_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_17_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_17_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_17_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_17_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_17_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_17_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_17_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_17_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_17_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_17_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_17_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_17_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_17_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_17_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_17_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_17_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_17_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_17_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_17_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_17_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_17_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_17_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_17_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_17_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_17_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_17_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_17_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_17_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_17_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_17_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_17_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_17_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_17_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_17_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_17_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_17_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_17_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_17_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_17_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_17_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_17_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_17_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_17_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_17_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_17_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_17_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_17_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_17_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_17_m_axi_gmem_BUSER)
	);
	qsort peArray_18(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_18_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_18_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_18_TREADY),
		.argOut_TVALID(_peArray_18_argOut_TVALID),
		.argOut_TDATA(_peArray_18_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_18_TREADY),
		.taskOut_TVALID(_peArray_18_taskOut_TVALID),
		.taskOut_TDATA(_peArray_18_taskOut_TDATA),
		.taskIn_TREADY(_peArray_18_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_18_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_18_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_18_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_18_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_18_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_18_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_18_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_18_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_18_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_18_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_18_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_18_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_18_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_18_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_18_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_18_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_18_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_18_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_18_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_18_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_18_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_18_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_18_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_18_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_18_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_18_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_18_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_18_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_18_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_18_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_18_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_18_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_18_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_18_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_18_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_18_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_18_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_18_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_18_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_18_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_18_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_18_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_18_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_18_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_18_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_18_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_18_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_18_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_18_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_18_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_18_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_18_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_18_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_18_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_18_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_18_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_18_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_18_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_18_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_18_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_18_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_18_m_axi_gmem_BUSER)
	);
	qsort peArray_19(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_19_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_19_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_19_TREADY),
		.argOut_TVALID(_peArray_19_argOut_TVALID),
		.argOut_TDATA(_peArray_19_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_19_TREADY),
		.taskOut_TVALID(_peArray_19_taskOut_TVALID),
		.taskOut_TDATA(_peArray_19_taskOut_TDATA),
		.taskIn_TREADY(_peArray_19_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_19_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_19_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_19_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_19_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_19_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_19_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_19_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_19_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_19_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_19_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_19_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_19_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_19_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_19_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_19_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_19_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_19_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_19_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_19_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_19_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_19_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_19_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_19_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_19_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_19_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_19_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_19_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_19_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_19_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_19_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_19_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_19_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_19_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_19_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_19_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_19_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_19_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_19_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_19_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_19_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_19_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_19_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_19_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_19_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_19_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_19_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_19_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_19_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_19_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_19_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_19_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_19_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_19_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_19_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_19_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_19_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_19_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_19_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_19_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_19_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_19_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_19_m_axi_gmem_BUSER)
	);
	qsort peArray_20(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_20_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_20_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_20_TREADY),
		.argOut_TVALID(_peArray_20_argOut_TVALID),
		.argOut_TDATA(_peArray_20_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_20_TREADY),
		.taskOut_TVALID(_peArray_20_taskOut_TVALID),
		.taskOut_TDATA(_peArray_20_taskOut_TDATA),
		.taskIn_TREADY(_peArray_20_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_20_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_20_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_20_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_20_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_20_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_20_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_20_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_20_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_20_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_20_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_20_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_20_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_20_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_20_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_20_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_20_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_20_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_20_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_20_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_20_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_20_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_20_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_20_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_20_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_20_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_20_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_20_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_20_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_20_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_20_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_20_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_20_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_20_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_20_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_20_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_20_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_20_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_20_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_20_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_20_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_20_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_20_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_20_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_20_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_20_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_20_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_20_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_20_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_20_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_20_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_20_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_20_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_20_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_20_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_20_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_20_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_20_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_20_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_20_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_20_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_20_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_20_m_axi_gmem_BUSER)
	);
	qsort peArray_21(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_21_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_21_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_21_TREADY),
		.argOut_TVALID(_peArray_21_argOut_TVALID),
		.argOut_TDATA(_peArray_21_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_21_TREADY),
		.taskOut_TVALID(_peArray_21_taskOut_TVALID),
		.taskOut_TDATA(_peArray_21_taskOut_TDATA),
		.taskIn_TREADY(_peArray_21_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_21_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_21_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_21_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_21_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_21_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_21_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_21_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_21_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_21_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_21_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_21_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_21_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_21_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_21_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_21_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_21_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_21_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_21_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_21_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_21_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_21_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_21_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_21_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_21_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_21_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_21_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_21_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_21_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_21_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_21_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_21_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_21_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_21_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_21_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_21_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_21_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_21_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_21_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_21_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_21_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_21_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_21_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_21_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_21_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_21_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_21_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_21_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_21_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_21_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_21_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_21_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_21_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_21_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_21_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_21_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_21_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_21_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_21_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_21_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_21_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_21_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_21_m_axi_gmem_BUSER)
	);
	qsort peArray_22(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_22_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_22_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_22_TREADY),
		.argOut_TVALID(_peArray_22_argOut_TVALID),
		.argOut_TDATA(_peArray_22_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_22_TREADY),
		.taskOut_TVALID(_peArray_22_taskOut_TVALID),
		.taskOut_TDATA(_peArray_22_taskOut_TDATA),
		.taskIn_TREADY(_peArray_22_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_22_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_22_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_22_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_22_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_22_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_22_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_22_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_22_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_22_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_22_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_22_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_22_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_22_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_22_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_22_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_22_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_22_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_22_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_22_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_22_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_22_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_22_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_22_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_22_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_22_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_22_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_22_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_22_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_22_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_22_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_22_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_22_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_22_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_22_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_22_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_22_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_22_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_22_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_22_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_22_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_22_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_22_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_22_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_22_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_22_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_22_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_22_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_22_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_22_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_22_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_22_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_22_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_22_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_22_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_22_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_22_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_22_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_22_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_22_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_22_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_22_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_22_m_axi_gmem_BUSER)
	);
	qsort peArray_23(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_23_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_23_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_23_TREADY),
		.argOut_TVALID(_peArray_23_argOut_TVALID),
		.argOut_TDATA(_peArray_23_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_23_TREADY),
		.taskOut_TVALID(_peArray_23_taskOut_TVALID),
		.taskOut_TDATA(_peArray_23_taskOut_TDATA),
		.taskIn_TREADY(_peArray_23_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_23_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_23_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_23_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_23_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_23_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_23_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_23_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_23_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_23_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_23_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_23_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_23_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_23_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_23_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_23_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_23_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_23_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_23_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_23_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_23_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_23_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_23_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_23_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_23_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_23_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_23_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_23_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_23_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_23_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_23_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_23_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_23_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_23_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_23_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_23_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_23_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_23_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_23_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_23_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_23_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_23_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_23_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_23_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_23_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_23_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_23_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_23_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_23_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_23_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_23_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_23_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_23_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_23_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_23_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_23_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_23_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_23_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_23_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_23_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_23_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_23_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_23_m_axi_gmem_BUSER)
	);
	qsort peArray_24(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_24_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_24_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_24_TREADY),
		.argOut_TVALID(_peArray_24_argOut_TVALID),
		.argOut_TDATA(_peArray_24_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_24_TREADY),
		.taskOut_TVALID(_peArray_24_taskOut_TVALID),
		.taskOut_TDATA(_peArray_24_taskOut_TDATA),
		.taskIn_TREADY(_peArray_24_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_24_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_24_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_24_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_24_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_24_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_24_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_24_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_24_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_24_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_24_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_24_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_24_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_24_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_24_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_24_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_24_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_24_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_24_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_24_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_24_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_24_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_24_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_24_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_24_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_24_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_24_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_24_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_24_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_24_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_24_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_24_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_24_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_24_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_24_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_24_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_24_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_24_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_24_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_24_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_24_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_24_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_24_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_24_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_24_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_24_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_24_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_24_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_24_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_24_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_24_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_24_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_24_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_24_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_24_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_24_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_24_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_24_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_24_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_24_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_24_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_24_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_24_m_axi_gmem_BUSER)
	);
	qsort peArray_25(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_25_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_25_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_25_TREADY),
		.argOut_TVALID(_peArray_25_argOut_TVALID),
		.argOut_TDATA(_peArray_25_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_25_TREADY),
		.taskOut_TVALID(_peArray_25_taskOut_TVALID),
		.taskOut_TDATA(_peArray_25_taskOut_TDATA),
		.taskIn_TREADY(_peArray_25_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_25_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_25_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_25_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_25_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_25_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_25_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_25_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_25_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_25_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_25_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_25_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_25_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_25_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_25_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_25_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_25_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_25_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_25_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_25_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_25_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_25_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_25_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_25_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_25_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_25_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_25_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_25_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_25_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_25_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_25_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_25_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_25_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_25_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_25_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_25_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_25_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_25_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_25_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_25_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_25_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_25_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_25_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_25_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_25_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_25_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_25_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_25_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_25_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_25_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_25_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_25_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_25_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_25_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_25_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_25_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_25_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_25_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_25_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_25_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_25_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_25_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_25_m_axi_gmem_BUSER)
	);
	qsort peArray_26(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_26_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_26_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_26_TREADY),
		.argOut_TVALID(_peArray_26_argOut_TVALID),
		.argOut_TDATA(_peArray_26_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_26_TREADY),
		.taskOut_TVALID(_peArray_26_taskOut_TVALID),
		.taskOut_TDATA(_peArray_26_taskOut_TDATA),
		.taskIn_TREADY(_peArray_26_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_26_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_26_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_26_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_26_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_26_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_26_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_26_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_26_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_26_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_26_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_26_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_26_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_26_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_26_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_26_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_26_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_26_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_26_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_26_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_26_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_26_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_26_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_26_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_26_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_26_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_26_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_26_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_26_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_26_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_26_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_26_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_26_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_26_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_26_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_26_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_26_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_26_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_26_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_26_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_26_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_26_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_26_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_26_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_26_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_26_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_26_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_26_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_26_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_26_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_26_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_26_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_26_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_26_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_26_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_26_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_26_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_26_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_26_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_26_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_26_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_26_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_26_m_axi_gmem_BUSER)
	);
	qsort peArray_27(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_27_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_27_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_27_TREADY),
		.argOut_TVALID(_peArray_27_argOut_TVALID),
		.argOut_TDATA(_peArray_27_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_27_TREADY),
		.taskOut_TVALID(_peArray_27_taskOut_TVALID),
		.taskOut_TDATA(_peArray_27_taskOut_TDATA),
		.taskIn_TREADY(_peArray_27_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_27_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_27_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_27_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_27_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_27_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_27_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_27_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_27_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_27_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_27_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_27_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_27_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_27_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_27_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_27_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_27_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_27_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_27_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_27_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_27_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_27_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_27_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_27_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_27_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_27_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_27_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_27_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_27_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_27_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_27_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_27_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_27_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_27_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_27_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_27_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_27_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_27_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_27_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_27_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_27_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_27_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_27_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_27_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_27_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_27_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_27_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_27_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_27_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_27_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_27_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_27_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_27_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_27_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_27_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_27_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_27_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_27_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_27_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_27_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_27_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_27_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_27_m_axi_gmem_BUSER)
	);
	qsort peArray_28(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_28_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_28_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_28_TREADY),
		.argOut_TVALID(_peArray_28_argOut_TVALID),
		.argOut_TDATA(_peArray_28_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_28_TREADY),
		.taskOut_TVALID(_peArray_28_taskOut_TVALID),
		.taskOut_TDATA(_peArray_28_taskOut_TDATA),
		.taskIn_TREADY(_peArray_28_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_28_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_28_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_28_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_28_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_28_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_28_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_28_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_28_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_28_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_28_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_28_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_28_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_28_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_28_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_28_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_28_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_28_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_28_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_28_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_28_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_28_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_28_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_28_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_28_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_28_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_28_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_28_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_28_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_28_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_28_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_28_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_28_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_28_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_28_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_28_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_28_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_28_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_28_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_28_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_28_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_28_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_28_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_28_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_28_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_28_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_28_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_28_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_28_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_28_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_28_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_28_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_28_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_28_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_28_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_28_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_28_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_28_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_28_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_28_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_28_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_28_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_28_m_axi_gmem_BUSER)
	);
	qsort peArray_29(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_29_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_29_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_29_TREADY),
		.argOut_TVALID(_peArray_29_argOut_TVALID),
		.argOut_TDATA(_peArray_29_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_29_TREADY),
		.taskOut_TVALID(_peArray_29_taskOut_TVALID),
		.taskOut_TDATA(_peArray_29_taskOut_TDATA),
		.taskIn_TREADY(_peArray_29_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_29_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_29_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_29_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_29_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_29_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_29_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_29_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_29_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_29_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_29_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_29_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_29_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_29_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_29_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_29_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_29_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_29_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_29_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_29_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_29_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_29_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_29_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_29_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_29_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_29_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_29_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_29_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_29_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_29_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_29_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_29_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_29_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_29_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_29_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_29_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_29_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_29_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_29_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_29_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_29_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_29_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_29_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_29_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_29_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_29_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_29_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_29_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_29_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_29_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_29_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_29_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_29_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_29_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_29_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_29_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_29_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_29_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_29_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_29_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_29_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_29_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_29_m_axi_gmem_BUSER)
	);
	qsort peArray_30(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_30_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_30_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_30_TREADY),
		.argOut_TVALID(_peArray_30_argOut_TVALID),
		.argOut_TDATA(_peArray_30_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_30_TREADY),
		.taskOut_TVALID(_peArray_30_taskOut_TVALID),
		.taskOut_TDATA(_peArray_30_taskOut_TDATA),
		.taskIn_TREADY(_peArray_30_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_30_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_30_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_30_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_30_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_30_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_30_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_30_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_30_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_30_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_30_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_30_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_30_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_30_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_30_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_30_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_30_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_30_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_30_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_30_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_30_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_30_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_30_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_30_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_30_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_30_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_30_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_30_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_30_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_30_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_30_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_30_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_30_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_30_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_30_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_30_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_30_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_30_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_30_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_30_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_30_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_30_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_30_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_30_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_30_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_30_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_30_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_30_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_30_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_30_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_30_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_30_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_30_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_30_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_30_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_30_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_30_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_30_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_30_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_30_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_30_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_30_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_30_m_axi_gmem_BUSER)
	);
	qsort peArray_31(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_31_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_31_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_31_TREADY),
		.argOut_TVALID(_peArray_31_argOut_TVALID),
		.argOut_TDATA(_peArray_31_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_31_TREADY),
		.taskOut_TVALID(_peArray_31_taskOut_TVALID),
		.taskOut_TDATA(_peArray_31_taskOut_TDATA),
		.taskIn_TREADY(_peArray_31_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_31_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_31_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_31_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_31_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_31_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_31_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_31_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_31_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_31_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_31_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_31_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_31_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_31_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_31_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_31_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_31_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_31_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_31_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_31_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_31_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_31_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_31_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_31_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_31_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_31_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_31_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_31_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_31_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_31_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_31_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_31_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_31_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_31_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_31_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_31_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_31_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_31_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_31_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_31_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_31_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_31_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_31_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_31_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_31_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_31_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_31_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_31_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_31_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_31_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_31_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_31_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_31_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_31_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_31_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_31_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_31_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_31_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_31_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_31_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_31_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_31_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_31_m_axi_gmem_BUSER)
	);
	qsort peArray_32(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_32_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_32_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_32_TREADY),
		.argOut_TVALID(_peArray_32_argOut_TVALID),
		.argOut_TDATA(_peArray_32_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_32_TREADY),
		.taskOut_TVALID(_peArray_32_taskOut_TVALID),
		.taskOut_TDATA(_peArray_32_taskOut_TDATA),
		.taskIn_TREADY(_peArray_32_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_32_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_32_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_32_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_32_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_32_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_32_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_32_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_32_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_32_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_32_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_32_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_32_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_32_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_32_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_32_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_32_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_32_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_32_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_32_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_32_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_32_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_32_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_32_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_32_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_32_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_32_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_32_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_32_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_32_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_32_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_32_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_32_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_32_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_32_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_32_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_32_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_32_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_32_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_32_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_32_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_32_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_32_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_32_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_32_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_32_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_32_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_32_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_32_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_32_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_32_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_32_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_32_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_32_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_32_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_32_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_32_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_32_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_32_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_32_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_32_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_32_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_32_m_axi_gmem_BUSER)
	);
	qsort peArray_33(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_33_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_33_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_33_TREADY),
		.argOut_TVALID(_peArray_33_argOut_TVALID),
		.argOut_TDATA(_peArray_33_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_33_TREADY),
		.taskOut_TVALID(_peArray_33_taskOut_TVALID),
		.taskOut_TDATA(_peArray_33_taskOut_TDATA),
		.taskIn_TREADY(_peArray_33_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_33_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_33_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_33_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_33_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_33_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_33_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_33_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_33_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_33_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_33_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_33_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_33_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_33_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_33_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_33_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_33_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_33_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_33_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_33_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_33_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_33_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_33_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_33_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_33_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_33_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_33_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_33_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_33_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_33_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_33_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_33_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_33_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_33_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_33_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_33_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_33_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_33_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_33_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_33_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_33_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_33_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_33_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_33_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_33_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_33_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_33_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_33_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_33_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_33_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_33_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_33_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_33_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_33_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_33_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_33_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_33_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_33_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_33_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_33_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_33_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_33_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_33_m_axi_gmem_BUSER)
	);
	qsort peArray_34(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_34_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_34_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_34_TREADY),
		.argOut_TVALID(_peArray_34_argOut_TVALID),
		.argOut_TDATA(_peArray_34_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_34_TREADY),
		.taskOut_TVALID(_peArray_34_taskOut_TVALID),
		.taskOut_TDATA(_peArray_34_taskOut_TDATA),
		.taskIn_TREADY(_peArray_34_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_34_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_34_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_34_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_34_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_34_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_34_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_34_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_34_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_34_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_34_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_34_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_34_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_34_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_34_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_34_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_34_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_34_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_34_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_34_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_34_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_34_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_34_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_34_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_34_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_34_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_34_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_34_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_34_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_34_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_34_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_34_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_34_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_34_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_34_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_34_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_34_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_34_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_34_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_34_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_34_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_34_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_34_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_34_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_34_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_34_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_34_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_34_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_34_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_34_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_34_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_34_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_34_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_34_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_34_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_34_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_34_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_34_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_34_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_34_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_34_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_34_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_34_m_axi_gmem_BUSER)
	);
	qsort peArray_35(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_35_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_35_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_35_TREADY),
		.argOut_TVALID(_peArray_35_argOut_TVALID),
		.argOut_TDATA(_peArray_35_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_35_TREADY),
		.taskOut_TVALID(_peArray_35_taskOut_TVALID),
		.taskOut_TDATA(_peArray_35_taskOut_TDATA),
		.taskIn_TREADY(_peArray_35_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_35_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_35_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_35_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_35_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_35_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_35_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_35_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_35_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_35_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_35_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_35_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_35_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_35_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_35_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_35_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_35_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_35_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_35_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_35_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_35_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_35_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_35_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_35_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_35_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_35_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_35_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_35_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_35_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_35_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_35_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_35_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_35_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_35_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_35_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_35_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_35_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_35_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_35_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_35_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_35_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_35_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_35_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_35_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_35_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_35_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_35_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_35_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_35_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_35_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_35_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_35_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_35_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_35_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_35_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_35_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_35_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_35_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_35_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_35_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_35_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_35_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_35_m_axi_gmem_BUSER)
	);
	qsort peArray_36(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_36_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_36_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_36_TREADY),
		.argOut_TVALID(_peArray_36_argOut_TVALID),
		.argOut_TDATA(_peArray_36_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_36_TREADY),
		.taskOut_TVALID(_peArray_36_taskOut_TVALID),
		.taskOut_TDATA(_peArray_36_taskOut_TDATA),
		.taskIn_TREADY(_peArray_36_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_36_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_36_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_36_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_36_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_36_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_36_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_36_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_36_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_36_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_36_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_36_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_36_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_36_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_36_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_36_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_36_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_36_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_36_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_36_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_36_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_36_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_36_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_36_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_36_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_36_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_36_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_36_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_36_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_36_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_36_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_36_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_36_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_36_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_36_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_36_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_36_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_36_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_36_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_36_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_36_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_36_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_36_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_36_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_36_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_36_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_36_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_36_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_36_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_36_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_36_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_36_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_36_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_36_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_36_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_36_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_36_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_36_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_36_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_36_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_36_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_36_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_36_m_axi_gmem_BUSER)
	);
	qsort peArray_37(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_37_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_37_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_37_TREADY),
		.argOut_TVALID(_peArray_37_argOut_TVALID),
		.argOut_TDATA(_peArray_37_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_37_TREADY),
		.taskOut_TVALID(_peArray_37_taskOut_TVALID),
		.taskOut_TDATA(_peArray_37_taskOut_TDATA),
		.taskIn_TREADY(_peArray_37_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_37_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_37_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_37_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_37_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_37_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_37_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_37_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_37_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_37_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_37_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_37_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_37_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_37_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_37_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_37_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_37_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_37_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_37_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_37_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_37_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_37_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_37_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_37_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_37_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_37_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_37_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_37_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_37_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_37_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_37_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_37_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_37_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_37_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_37_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_37_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_37_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_37_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_37_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_37_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_37_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_37_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_37_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_37_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_37_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_37_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_37_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_37_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_37_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_37_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_37_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_37_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_37_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_37_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_37_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_37_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_37_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_37_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_37_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_37_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_37_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_37_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_37_m_axi_gmem_BUSER)
	);
	qsort peArray_38(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_38_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_38_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_38_TREADY),
		.argOut_TVALID(_peArray_38_argOut_TVALID),
		.argOut_TDATA(_peArray_38_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_38_TREADY),
		.taskOut_TVALID(_peArray_38_taskOut_TVALID),
		.taskOut_TDATA(_peArray_38_taskOut_TDATA),
		.taskIn_TREADY(_peArray_38_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_38_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_38_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_38_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_38_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_38_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_38_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_38_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_38_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_38_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_38_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_38_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_38_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_38_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_38_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_38_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_38_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_38_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_38_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_38_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_38_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_38_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_38_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_38_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_38_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_38_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_38_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_38_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_38_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_38_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_38_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_38_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_38_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_38_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_38_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_38_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_38_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_38_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_38_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_38_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_38_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_38_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_38_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_38_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_38_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_38_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_38_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_38_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_38_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_38_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_38_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_38_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_38_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_38_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_38_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_38_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_38_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_38_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_38_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_38_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_38_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_38_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_38_m_axi_gmem_BUSER)
	);
	qsort peArray_39(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_39_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_39_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_39_TREADY),
		.argOut_TVALID(_peArray_39_argOut_TVALID),
		.argOut_TDATA(_peArray_39_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_39_TREADY),
		.taskOut_TVALID(_peArray_39_taskOut_TVALID),
		.taskOut_TDATA(_peArray_39_taskOut_TDATA),
		.taskIn_TREADY(_peArray_39_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_39_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_39_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_39_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_39_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_39_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_39_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_39_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_39_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_39_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_39_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_39_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_39_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_39_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_39_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_39_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_39_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_39_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_39_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_39_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_39_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_39_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_39_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_39_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_39_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_39_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_39_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_39_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_39_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_39_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_39_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_39_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_39_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_39_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_39_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_39_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_39_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_39_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_39_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_39_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_39_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_39_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_39_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_39_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_39_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_39_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_39_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_39_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_39_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_39_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_39_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_39_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_39_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_39_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_39_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_39_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_39_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_39_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_39_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_39_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_39_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_39_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_39_m_axi_gmem_BUSER)
	);
	qsort peArray_40(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_40_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_40_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_40_TREADY),
		.argOut_TVALID(_peArray_40_argOut_TVALID),
		.argOut_TDATA(_peArray_40_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_40_TREADY),
		.taskOut_TVALID(_peArray_40_taskOut_TVALID),
		.taskOut_TDATA(_peArray_40_taskOut_TDATA),
		.taskIn_TREADY(_peArray_40_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_40_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_40_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_40_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_40_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_40_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_40_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_40_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_40_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_40_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_40_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_40_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_40_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_40_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_40_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_40_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_40_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_40_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_40_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_40_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_40_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_40_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_40_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_40_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_40_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_40_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_40_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_40_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_40_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_40_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_40_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_40_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_40_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_40_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_40_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_40_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_40_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_40_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_40_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_40_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_40_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_40_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_40_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_40_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_40_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_40_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_40_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_40_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_40_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_40_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_40_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_40_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_40_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_40_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_40_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_40_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_40_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_40_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_40_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_40_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_40_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_40_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_40_m_axi_gmem_BUSER)
	);
	qsort peArray_41(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_41_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_41_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_41_TREADY),
		.argOut_TVALID(_peArray_41_argOut_TVALID),
		.argOut_TDATA(_peArray_41_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_41_TREADY),
		.taskOut_TVALID(_peArray_41_taskOut_TVALID),
		.taskOut_TDATA(_peArray_41_taskOut_TDATA),
		.taskIn_TREADY(_peArray_41_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_41_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_41_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_41_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_41_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_41_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_41_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_41_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_41_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_41_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_41_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_41_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_41_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_41_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_41_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_41_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_41_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_41_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_41_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_41_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_41_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_41_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_41_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_41_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_41_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_41_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_41_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_41_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_41_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_41_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_41_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_41_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_41_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_41_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_41_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_41_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_41_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_41_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_41_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_41_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_41_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_41_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_41_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_41_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_41_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_41_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_41_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_41_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_41_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_41_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_41_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_41_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_41_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_41_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_41_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_41_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_41_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_41_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_41_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_41_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_41_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_41_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_41_m_axi_gmem_BUSER)
	);
	qsort peArray_42(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_42_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_42_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_42_TREADY),
		.argOut_TVALID(_peArray_42_argOut_TVALID),
		.argOut_TDATA(_peArray_42_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_42_TREADY),
		.taskOut_TVALID(_peArray_42_taskOut_TVALID),
		.taskOut_TDATA(_peArray_42_taskOut_TDATA),
		.taskIn_TREADY(_peArray_42_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_42_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_42_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_42_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_42_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_42_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_42_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_42_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_42_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_42_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_42_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_42_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_42_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_42_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_42_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_42_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_42_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_42_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_42_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_42_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_42_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_42_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_42_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_42_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_42_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_42_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_42_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_42_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_42_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_42_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_42_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_42_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_42_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_42_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_42_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_42_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_42_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_42_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_42_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_42_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_42_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_42_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_42_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_42_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_42_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_42_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_42_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_42_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_42_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_42_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_42_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_42_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_42_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_42_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_42_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_42_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_42_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_42_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_42_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_42_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_42_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_42_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_42_m_axi_gmem_BUSER)
	);
	qsort peArray_43(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_43_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_43_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_43_TREADY),
		.argOut_TVALID(_peArray_43_argOut_TVALID),
		.argOut_TDATA(_peArray_43_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_43_TREADY),
		.taskOut_TVALID(_peArray_43_taskOut_TVALID),
		.taskOut_TDATA(_peArray_43_taskOut_TDATA),
		.taskIn_TREADY(_peArray_43_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_43_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_43_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_43_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_43_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_43_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_43_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_43_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_43_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_43_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_43_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_43_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_43_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_43_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_43_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_43_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_43_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_43_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_43_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_43_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_43_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_43_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_43_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_43_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_43_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_43_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_43_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_43_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_43_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_43_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_43_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_43_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_43_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_43_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_43_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_43_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_43_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_43_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_43_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_43_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_43_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_43_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_43_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_43_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_43_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_43_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_43_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_43_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_43_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_43_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_43_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_43_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_43_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_43_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_43_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_43_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_43_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_43_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_43_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_43_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_43_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_43_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_43_m_axi_gmem_BUSER)
	);
	qsort peArray_44(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_44_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_44_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_44_TREADY),
		.argOut_TVALID(_peArray_44_argOut_TVALID),
		.argOut_TDATA(_peArray_44_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_44_TREADY),
		.taskOut_TVALID(_peArray_44_taskOut_TVALID),
		.taskOut_TDATA(_peArray_44_taskOut_TDATA),
		.taskIn_TREADY(_peArray_44_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_44_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_44_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_44_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_44_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_44_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_44_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_44_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_44_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_44_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_44_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_44_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_44_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_44_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_44_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_44_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_44_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_44_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_44_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_44_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_44_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_44_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_44_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_44_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_44_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_44_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_44_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_44_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_44_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_44_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_44_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_44_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_44_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_44_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_44_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_44_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_44_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_44_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_44_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_44_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_44_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_44_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_44_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_44_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_44_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_44_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_44_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_44_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_44_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_44_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_44_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_44_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_44_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_44_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_44_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_44_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_44_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_44_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_44_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_44_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_44_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_44_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_44_m_axi_gmem_BUSER)
	);
	qsort peArray_45(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_45_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_45_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_45_TREADY),
		.argOut_TVALID(_peArray_45_argOut_TVALID),
		.argOut_TDATA(_peArray_45_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_45_TREADY),
		.taskOut_TVALID(_peArray_45_taskOut_TVALID),
		.taskOut_TDATA(_peArray_45_taskOut_TDATA),
		.taskIn_TREADY(_peArray_45_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_45_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_45_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_45_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_45_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_45_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_45_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_45_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_45_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_45_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_45_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_45_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_45_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_45_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_45_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_45_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_45_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_45_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_45_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_45_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_45_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_45_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_45_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_45_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_45_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_45_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_45_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_45_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_45_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_45_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_45_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_45_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_45_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_45_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_45_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_45_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_45_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_45_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_45_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_45_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_45_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_45_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_45_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_45_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_45_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_45_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_45_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_45_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_45_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_45_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_45_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_45_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_45_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_45_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_45_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_45_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_45_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_45_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_45_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_45_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_45_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_45_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_45_m_axi_gmem_BUSER)
	);
	qsort peArray_46(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_46_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_46_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_46_TREADY),
		.argOut_TVALID(_peArray_46_argOut_TVALID),
		.argOut_TDATA(_peArray_46_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_46_TREADY),
		.taskOut_TVALID(_peArray_46_taskOut_TVALID),
		.taskOut_TDATA(_peArray_46_taskOut_TDATA),
		.taskIn_TREADY(_peArray_46_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_46_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_46_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_46_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_46_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_46_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_46_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_46_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_46_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_46_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_46_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_46_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_46_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_46_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_46_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_46_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_46_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_46_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_46_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_46_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_46_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_46_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_46_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_46_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_46_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_46_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_46_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_46_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_46_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_46_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_46_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_46_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_46_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_46_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_46_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_46_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_46_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_46_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_46_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_46_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_46_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_46_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_46_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_46_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_46_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_46_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_46_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_46_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_46_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_46_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_46_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_46_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_46_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_46_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_46_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_46_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_46_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_46_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_46_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_46_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_46_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_46_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_46_m_axi_gmem_BUSER)
	);
	qsort peArray_47(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_47_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_47_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_47_TREADY),
		.argOut_TVALID(_peArray_47_argOut_TVALID),
		.argOut_TDATA(_peArray_47_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_47_TREADY),
		.taskOut_TVALID(_peArray_47_taskOut_TVALID),
		.taskOut_TDATA(_peArray_47_taskOut_TDATA),
		.taskIn_TREADY(_peArray_47_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_47_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_47_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_47_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_47_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_47_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_47_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_47_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_47_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_47_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_47_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_47_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_47_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_47_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_47_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_47_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_47_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_47_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_47_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_47_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_47_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_47_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_47_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_47_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_47_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_47_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_47_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_47_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_47_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_47_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_47_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_47_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_47_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_47_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_47_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_47_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_47_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_47_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_47_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_47_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_47_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_47_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_47_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_47_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_47_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_47_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_47_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_47_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_47_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_47_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_47_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_47_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_47_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_47_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_47_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_47_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_47_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_47_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_47_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_47_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_47_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_47_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_47_m_axi_gmem_BUSER)
	);
	qsort peArray_48(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_48_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_48_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_48_TREADY),
		.argOut_TVALID(_peArray_48_argOut_TVALID),
		.argOut_TDATA(_peArray_48_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_48_TREADY),
		.taskOut_TVALID(_peArray_48_taskOut_TVALID),
		.taskOut_TDATA(_peArray_48_taskOut_TDATA),
		.taskIn_TREADY(_peArray_48_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_48_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_48_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_48_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_48_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_48_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_48_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_48_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_48_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_48_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_48_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_48_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_48_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_48_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_48_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_48_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_48_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_48_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_48_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_48_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_48_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_48_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_48_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_48_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_48_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_48_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_48_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_48_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_48_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_48_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_48_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_48_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_48_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_48_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_48_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_48_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_48_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_48_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_48_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_48_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_48_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_48_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_48_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_48_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_48_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_48_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_48_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_48_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_48_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_48_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_48_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_48_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_48_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_48_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_48_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_48_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_48_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_48_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_48_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_48_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_48_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_48_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_48_m_axi_gmem_BUSER)
	);
	qsort peArray_49(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_49_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_49_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_49_TREADY),
		.argOut_TVALID(_peArray_49_argOut_TVALID),
		.argOut_TDATA(_peArray_49_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_49_TREADY),
		.taskOut_TVALID(_peArray_49_taskOut_TVALID),
		.taskOut_TDATA(_peArray_49_taskOut_TDATA),
		.taskIn_TREADY(_peArray_49_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_49_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_49_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_49_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_49_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_49_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_49_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_49_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_49_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_49_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_49_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_49_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_49_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_49_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_49_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_49_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_49_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_49_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_49_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_49_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_49_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_49_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_49_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_49_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_49_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_49_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_49_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_49_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_49_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_49_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_49_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_49_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_49_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_49_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_49_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_49_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_49_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_49_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_49_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_49_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_49_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_49_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_49_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_49_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_49_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_49_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_49_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_49_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_49_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_49_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_49_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_49_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_49_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_49_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_49_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_49_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_49_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_49_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_49_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_49_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_49_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_49_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_49_m_axi_gmem_BUSER)
	);
	qsort peArray_50(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_50_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_50_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_50_TREADY),
		.argOut_TVALID(_peArray_50_argOut_TVALID),
		.argOut_TDATA(_peArray_50_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_50_TREADY),
		.taskOut_TVALID(_peArray_50_taskOut_TVALID),
		.taskOut_TDATA(_peArray_50_taskOut_TDATA),
		.taskIn_TREADY(_peArray_50_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_50_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_50_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_50_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_50_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_50_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_50_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_50_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_50_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_50_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_50_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_50_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_50_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_50_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_50_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_50_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_50_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_50_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_50_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_50_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_50_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_50_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_50_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_50_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_50_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_50_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_50_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_50_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_50_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_50_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_50_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_50_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_50_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_50_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_50_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_50_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_50_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_50_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_50_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_50_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_50_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_50_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_50_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_50_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_50_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_50_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_50_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_50_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_50_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_50_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_50_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_50_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_50_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_50_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_50_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_50_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_50_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_50_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_50_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_50_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_50_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_50_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_50_m_axi_gmem_BUSER)
	);
	qsort peArray_51(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_51_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_51_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_51_TREADY),
		.argOut_TVALID(_peArray_51_argOut_TVALID),
		.argOut_TDATA(_peArray_51_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_51_TREADY),
		.taskOut_TVALID(_peArray_51_taskOut_TVALID),
		.taskOut_TDATA(_peArray_51_taskOut_TDATA),
		.taskIn_TREADY(_peArray_51_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_51_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_51_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_51_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_51_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_51_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_51_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_51_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_51_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_51_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_51_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_51_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_51_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_51_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_51_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_51_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_51_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_51_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_51_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_51_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_51_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_51_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_51_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_51_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_51_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_51_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_51_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_51_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_51_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_51_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_51_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_51_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_51_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_51_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_51_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_51_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_51_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_51_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_51_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_51_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_51_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_51_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_51_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_51_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_51_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_51_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_51_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_51_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_51_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_51_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_51_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_51_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_51_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_51_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_51_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_51_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_51_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_51_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_51_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_51_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_51_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_51_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_51_m_axi_gmem_BUSER)
	);
	qsort peArray_52(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_52_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_52_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_52_TREADY),
		.argOut_TVALID(_peArray_52_argOut_TVALID),
		.argOut_TDATA(_peArray_52_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_52_TREADY),
		.taskOut_TVALID(_peArray_52_taskOut_TVALID),
		.taskOut_TDATA(_peArray_52_taskOut_TDATA),
		.taskIn_TREADY(_peArray_52_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_52_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_52_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_52_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_52_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_52_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_52_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_52_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_52_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_52_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_52_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_52_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_52_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_52_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_52_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_52_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_52_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_52_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_52_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_52_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_52_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_52_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_52_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_52_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_52_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_52_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_52_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_52_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_52_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_52_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_52_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_52_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_52_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_52_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_52_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_52_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_52_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_52_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_52_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_52_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_52_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_52_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_52_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_52_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_52_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_52_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_52_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_52_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_52_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_52_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_52_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_52_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_52_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_52_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_52_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_52_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_52_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_52_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_52_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_52_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_52_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_52_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_52_m_axi_gmem_BUSER)
	);
	qsort peArray_53(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_53_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_53_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_53_TREADY),
		.argOut_TVALID(_peArray_53_argOut_TVALID),
		.argOut_TDATA(_peArray_53_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_53_TREADY),
		.taskOut_TVALID(_peArray_53_taskOut_TVALID),
		.taskOut_TDATA(_peArray_53_taskOut_TDATA),
		.taskIn_TREADY(_peArray_53_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_53_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_53_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_53_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_53_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_53_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_53_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_53_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_53_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_53_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_53_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_53_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_53_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_53_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_53_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_53_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_53_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_53_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_53_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_53_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_53_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_53_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_53_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_53_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_53_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_53_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_53_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_53_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_53_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_53_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_53_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_53_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_53_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_53_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_53_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_53_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_53_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_53_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_53_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_53_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_53_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_53_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_53_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_53_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_53_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_53_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_53_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_53_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_53_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_53_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_53_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_53_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_53_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_53_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_53_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_53_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_53_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_53_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_53_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_53_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_53_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_53_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_53_m_axi_gmem_BUSER)
	);
	qsort peArray_54(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_54_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_54_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_54_TREADY),
		.argOut_TVALID(_peArray_54_argOut_TVALID),
		.argOut_TDATA(_peArray_54_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_54_TREADY),
		.taskOut_TVALID(_peArray_54_taskOut_TVALID),
		.taskOut_TDATA(_peArray_54_taskOut_TDATA),
		.taskIn_TREADY(_peArray_54_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_54_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_54_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_54_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_54_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_54_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_54_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_54_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_54_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_54_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_54_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_54_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_54_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_54_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_54_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_54_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_54_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_54_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_54_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_54_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_54_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_54_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_54_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_54_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_54_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_54_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_54_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_54_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_54_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_54_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_54_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_54_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_54_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_54_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_54_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_54_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_54_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_54_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_54_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_54_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_54_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_54_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_54_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_54_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_54_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_54_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_54_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_54_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_54_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_54_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_54_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_54_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_54_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_54_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_54_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_54_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_54_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_54_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_54_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_54_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_54_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_54_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_54_m_axi_gmem_BUSER)
	);
	qsort peArray_55(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_55_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_55_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_55_TREADY),
		.argOut_TVALID(_peArray_55_argOut_TVALID),
		.argOut_TDATA(_peArray_55_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_55_TREADY),
		.taskOut_TVALID(_peArray_55_taskOut_TVALID),
		.taskOut_TDATA(_peArray_55_taskOut_TDATA),
		.taskIn_TREADY(_peArray_55_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_55_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_55_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_55_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_55_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_55_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_55_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_55_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_55_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_55_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_55_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_55_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_55_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_55_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_55_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_55_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_55_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_55_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_55_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_55_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_55_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_55_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_55_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_55_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_55_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_55_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_55_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_55_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_55_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_55_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_55_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_55_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_55_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_55_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_55_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_55_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_55_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_55_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_55_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_55_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_55_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_55_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_55_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_55_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_55_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_55_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_55_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_55_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_55_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_55_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_55_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_55_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_55_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_55_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_55_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_55_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_55_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_55_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_55_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_55_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_55_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_55_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_55_m_axi_gmem_BUSER)
	);
	qsort peArray_56(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_56_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_56_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_56_TREADY),
		.argOut_TVALID(_peArray_56_argOut_TVALID),
		.argOut_TDATA(_peArray_56_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_56_TREADY),
		.taskOut_TVALID(_peArray_56_taskOut_TVALID),
		.taskOut_TDATA(_peArray_56_taskOut_TDATA),
		.taskIn_TREADY(_peArray_56_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_56_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_56_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_56_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_56_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_56_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_56_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_56_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_56_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_56_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_56_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_56_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_56_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_56_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_56_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_56_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_56_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_56_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_56_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_56_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_56_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_56_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_56_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_56_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_56_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_56_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_56_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_56_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_56_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_56_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_56_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_56_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_56_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_56_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_56_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_56_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_56_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_56_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_56_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_56_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_56_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_56_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_56_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_56_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_56_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_56_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_56_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_56_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_56_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_56_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_56_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_56_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_56_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_56_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_56_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_56_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_56_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_56_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_56_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_56_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_56_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_56_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_56_m_axi_gmem_BUSER)
	);
	qsort peArray_57(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_57_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_57_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_57_TREADY),
		.argOut_TVALID(_peArray_57_argOut_TVALID),
		.argOut_TDATA(_peArray_57_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_57_TREADY),
		.taskOut_TVALID(_peArray_57_taskOut_TVALID),
		.taskOut_TDATA(_peArray_57_taskOut_TDATA),
		.taskIn_TREADY(_peArray_57_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_57_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_57_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_57_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_57_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_57_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_57_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_57_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_57_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_57_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_57_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_57_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_57_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_57_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_57_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_57_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_57_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_57_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_57_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_57_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_57_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_57_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_57_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_57_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_57_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_57_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_57_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_57_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_57_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_57_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_57_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_57_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_57_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_57_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_57_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_57_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_57_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_57_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_57_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_57_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_57_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_57_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_57_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_57_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_57_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_57_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_57_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_57_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_57_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_57_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_57_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_57_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_57_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_57_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_57_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_57_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_57_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_57_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_57_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_57_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_57_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_57_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_57_m_axi_gmem_BUSER)
	);
	qsort peArray_58(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_58_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_58_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_58_TREADY),
		.argOut_TVALID(_peArray_58_argOut_TVALID),
		.argOut_TDATA(_peArray_58_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_58_TREADY),
		.taskOut_TVALID(_peArray_58_taskOut_TVALID),
		.taskOut_TDATA(_peArray_58_taskOut_TDATA),
		.taskIn_TREADY(_peArray_58_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_58_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_58_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_58_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_58_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_58_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_58_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_58_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_58_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_58_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_58_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_58_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_58_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_58_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_58_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_58_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_58_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_58_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_58_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_58_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_58_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_58_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_58_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_58_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_58_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_58_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_58_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_58_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_58_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_58_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_58_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_58_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_58_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_58_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_58_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_58_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_58_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_58_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_58_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_58_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_58_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_58_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_58_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_58_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_58_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_58_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_58_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_58_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_58_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_58_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_58_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_58_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_58_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_58_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_58_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_58_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_58_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_58_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_58_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_58_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_58_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_58_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_58_m_axi_gmem_BUSER)
	);
	qsort peArray_59(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_59_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_59_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_59_TREADY),
		.argOut_TVALID(_peArray_59_argOut_TVALID),
		.argOut_TDATA(_peArray_59_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_59_TREADY),
		.taskOut_TVALID(_peArray_59_taskOut_TVALID),
		.taskOut_TDATA(_peArray_59_taskOut_TDATA),
		.taskIn_TREADY(_peArray_59_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_59_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_59_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_59_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_59_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_59_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_59_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_59_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_59_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_59_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_59_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_59_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_59_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_59_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_59_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_59_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_59_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_59_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_59_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_59_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_59_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_59_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_59_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_59_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_59_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_59_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_59_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_59_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_59_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_59_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_59_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_59_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_59_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_59_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_59_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_59_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_59_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_59_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_59_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_59_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_59_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_59_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_59_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_59_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_59_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_59_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_59_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_59_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_59_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_59_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_59_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_59_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_59_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_59_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_59_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_59_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_59_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_59_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_59_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_59_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_59_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_59_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_59_m_axi_gmem_BUSER)
	);
	qsort peArray_60(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_60_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_60_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_60_TREADY),
		.argOut_TVALID(_peArray_60_argOut_TVALID),
		.argOut_TDATA(_peArray_60_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_60_TREADY),
		.taskOut_TVALID(_peArray_60_taskOut_TVALID),
		.taskOut_TDATA(_peArray_60_taskOut_TDATA),
		.taskIn_TREADY(_peArray_60_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_60_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_60_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_60_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_60_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_60_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_60_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_60_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_60_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_60_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_60_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_60_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_60_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_60_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_60_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_60_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_60_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_60_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_60_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_60_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_60_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_60_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_60_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_60_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_60_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_60_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_60_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_60_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_60_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_60_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_60_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_60_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_60_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_60_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_60_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_60_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_60_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_60_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_60_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_60_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_60_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_60_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_60_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_60_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_60_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_60_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_60_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_60_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_60_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_60_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_60_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_60_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_60_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_60_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_60_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_60_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_60_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_60_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_60_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_60_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_60_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_60_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_60_m_axi_gmem_BUSER)
	);
	qsort peArray_61(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_61_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_61_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_61_TREADY),
		.argOut_TVALID(_peArray_61_argOut_TVALID),
		.argOut_TDATA(_peArray_61_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_61_TREADY),
		.taskOut_TVALID(_peArray_61_taskOut_TVALID),
		.taskOut_TDATA(_peArray_61_taskOut_TDATA),
		.taskIn_TREADY(_peArray_61_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_61_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_61_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_61_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_61_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_61_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_61_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_61_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_61_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_61_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_61_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_61_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_61_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_61_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_61_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_61_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_61_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_61_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_61_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_61_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_61_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_61_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_61_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_61_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_61_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_61_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_61_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_61_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_61_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_61_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_61_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_61_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_61_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_61_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_61_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_61_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_61_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_61_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_61_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_61_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_61_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_61_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_61_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_61_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_61_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_61_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_61_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_61_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_61_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_61_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_61_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_61_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_61_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_61_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_61_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_61_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_61_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_61_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_61_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_61_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_61_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_61_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_61_m_axi_gmem_BUSER)
	);
	qsort peArray_62(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_62_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_62_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_62_TREADY),
		.argOut_TVALID(_peArray_62_argOut_TVALID),
		.argOut_TDATA(_peArray_62_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_62_TREADY),
		.taskOut_TVALID(_peArray_62_taskOut_TVALID),
		.taskOut_TDATA(_peArray_62_taskOut_TDATA),
		.taskIn_TREADY(_peArray_62_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_62_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_62_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_62_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_62_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_62_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_62_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_62_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_62_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_62_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_62_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_62_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_62_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_62_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_62_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_62_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_62_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_62_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_62_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_62_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_62_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_62_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_62_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_62_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_62_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_62_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_62_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_62_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_62_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_62_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_62_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_62_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_62_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_62_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_62_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_62_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_62_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_62_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_62_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_62_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_62_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_62_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_62_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_62_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_62_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_62_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_62_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_62_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_62_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_62_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_62_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_62_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_62_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_62_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_62_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_62_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_62_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_62_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_62_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_62_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_62_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_62_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_62_m_axi_gmem_BUSER)
	);
	qsort peArray_63(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.ap_ready(),
		.ap_idle(),
		.ap_done(),
		.ap_start(1'h1),
		.closureIn_TREADY(_peArray_63_closureIn_TREADY),
		.closureIn_TVALID(_Allocator_io_export_closureOut_63_TVALID),
		.closureIn_TDATA(64'h0000000000000000),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_63_TREADY),
		.argOut_TVALID(_peArray_63_argOut_TVALID),
		.argOut_TDATA(_peArray_63_argOut_TDATA),
		.taskOut_TREADY(_Scheduler_io_export_taskIn_63_TREADY),
		.taskOut_TVALID(_peArray_63_taskOut_TVALID),
		.taskOut_TDATA(_peArray_63_taskOut_TDATA),
		.taskIn_TREADY(_peArray_63_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_io_export_taskOut_63_TVALID),
		.taskIn_TDATA(256'h0000000000000000000000000000000000000000000000000000000000000000),
		.s_axi_control_ARREADY(qsort_63_s_axi_control_ARREADY),
		.s_axi_control_ARVALID(qsort_63_s_axi_control_ARVALID),
		.s_axi_control_ARADDR(qsort_63_s_axi_control_ARADDR),
		.s_axi_control_RREADY(qsort_63_s_axi_control_RREADY),
		.s_axi_control_RVALID(qsort_63_s_axi_control_RVALID),
		.s_axi_control_RDATA(qsort_63_s_axi_control_RDATA),
		.s_axi_control_RRESP(qsort_63_s_axi_control_RRESP),
		.s_axi_control_AWREADY(qsort_63_s_axi_control_AWREADY),
		.s_axi_control_AWVALID(qsort_63_s_axi_control_AWVALID),
		.s_axi_control_AWADDR(qsort_63_s_axi_control_AWADDR),
		.s_axi_control_WREADY(qsort_63_s_axi_control_WREADY),
		.s_axi_control_WVALID(qsort_63_s_axi_control_WVALID),
		.s_axi_control_WDATA(qsort_63_s_axi_control_WDATA),
		.s_axi_control_WSTRB(qsort_63_s_axi_control_WSTRB),
		.s_axi_control_BREADY(qsort_63_s_axi_control_BREADY),
		.s_axi_control_BVALID(qsort_63_s_axi_control_BVALID),
		.s_axi_control_BRESP(qsort_63_s_axi_control_BRESP),
		.m_axi_gmem_ARREADY(qsort_63_m_axi_gmem_ARREADY),
		.m_axi_gmem_ARVALID(qsort_63_m_axi_gmem_ARVALID),
		.m_axi_gmem_ARID(qsort_63_m_axi_gmem_ARID),
		.m_axi_gmem_ARADDR(qsort_63_m_axi_gmem_ARADDR),
		.m_axi_gmem_ARLEN(qsort_63_m_axi_gmem_ARLEN),
		.m_axi_gmem_ARSIZE(qsort_63_m_axi_gmem_ARSIZE),
		.m_axi_gmem_ARBURST(qsort_63_m_axi_gmem_ARBURST),
		.m_axi_gmem_ARLOCK(qsort_63_m_axi_gmem_ARLOCK),
		.m_axi_gmem_ARCACHE(qsort_63_m_axi_gmem_ARCACHE),
		.m_axi_gmem_ARPROT(qsort_63_m_axi_gmem_ARPROT),
		.m_axi_gmem_ARQOS(qsort_63_m_axi_gmem_ARQOS),
		.m_axi_gmem_ARREGION(qsort_63_m_axi_gmem_ARREGION),
		.m_axi_gmem_ARUSER(qsort_63_m_axi_gmem_ARUSER),
		.m_axi_gmem_RREADY(qsort_63_m_axi_gmem_RREADY),
		.m_axi_gmem_RVALID(qsort_63_m_axi_gmem_RVALID),
		.m_axi_gmem_RID(qsort_63_m_axi_gmem_RID),
		.m_axi_gmem_RDATA(qsort_63_m_axi_gmem_RDATA),
		.m_axi_gmem_RRESP(qsort_63_m_axi_gmem_RRESP),
		.m_axi_gmem_RLAST(qsort_63_m_axi_gmem_RLAST),
		.m_axi_gmem_RUSER(qsort_63_m_axi_gmem_RUSER),
		.m_axi_gmem_AWREADY(qsort_63_m_axi_gmem_AWREADY),
		.m_axi_gmem_AWVALID(qsort_63_m_axi_gmem_AWVALID),
		.m_axi_gmem_AWID(qsort_63_m_axi_gmem_AWID),
		.m_axi_gmem_AWADDR(qsort_63_m_axi_gmem_AWADDR),
		.m_axi_gmem_AWLEN(qsort_63_m_axi_gmem_AWLEN),
		.m_axi_gmem_AWSIZE(qsort_63_m_axi_gmem_AWSIZE),
		.m_axi_gmem_AWBURST(qsort_63_m_axi_gmem_AWBURST),
		.m_axi_gmem_AWLOCK(qsort_63_m_axi_gmem_AWLOCK),
		.m_axi_gmem_AWCACHE(qsort_63_m_axi_gmem_AWCACHE),
		.m_axi_gmem_AWPROT(qsort_63_m_axi_gmem_AWPROT),
		.m_axi_gmem_AWQOS(qsort_63_m_axi_gmem_AWQOS),
		.m_axi_gmem_AWREGION(qsort_63_m_axi_gmem_AWREGION),
		.m_axi_gmem_AWUSER(qsort_63_m_axi_gmem_AWUSER),
		.m_axi_gmem_WREADY(qsort_63_m_axi_gmem_WREADY),
		.m_axi_gmem_WVALID(qsort_63_m_axi_gmem_WVALID),
		.m_axi_gmem_WDATA(qsort_63_m_axi_gmem_WDATA),
		.m_axi_gmem_WSTRB(qsort_63_m_axi_gmem_WSTRB),
		.m_axi_gmem_WLAST(qsort_63_m_axi_gmem_WLAST),
		.m_axi_gmem_WUSER(qsort_63_m_axi_gmem_WUSER),
		.m_axi_gmem_BREADY(qsort_63_m_axi_gmem_BREADY),
		.m_axi_gmem_BVALID(qsort_63_m_axi_gmem_BVALID),
		.m_axi_gmem_BID(qsort_63_m_axi_gmem_BID),
		.m_axi_gmem_BRESP(qsort_63_m_axi_gmem_BRESP),
		.m_axi_gmem_BUSER(qsort_63_m_axi_gmem_BUSER)
	);
	Scheduler Scheduler(
		.clock(clock),
		.reset(reset),
		.io_export_taskOut_0_TREADY(_peArray_0_taskIn_TREADY),
		.io_export_taskOut_0_TVALID(_Scheduler_io_export_taskOut_0_TVALID),
		.io_export_taskOut_1_TREADY(_peArray_1_taskIn_TREADY),
		.io_export_taskOut_1_TVALID(_Scheduler_io_export_taskOut_1_TVALID),
		.io_export_taskOut_2_TREADY(_peArray_2_taskIn_TREADY),
		.io_export_taskOut_2_TVALID(_Scheduler_io_export_taskOut_2_TVALID),
		.io_export_taskOut_3_TREADY(_peArray_3_taskIn_TREADY),
		.io_export_taskOut_3_TVALID(_Scheduler_io_export_taskOut_3_TVALID),
		.io_export_taskOut_4_TREADY(_peArray_4_taskIn_TREADY),
		.io_export_taskOut_4_TVALID(_Scheduler_io_export_taskOut_4_TVALID),
		.io_export_taskOut_5_TREADY(_peArray_5_taskIn_TREADY),
		.io_export_taskOut_5_TVALID(_Scheduler_io_export_taskOut_5_TVALID),
		.io_export_taskOut_6_TREADY(_peArray_6_taskIn_TREADY),
		.io_export_taskOut_6_TVALID(_Scheduler_io_export_taskOut_6_TVALID),
		.io_export_taskOut_7_TREADY(_peArray_7_taskIn_TREADY),
		.io_export_taskOut_7_TVALID(_Scheduler_io_export_taskOut_7_TVALID),
		.io_export_taskOut_8_TREADY(_peArray_8_taskIn_TREADY),
		.io_export_taskOut_8_TVALID(_Scheduler_io_export_taskOut_8_TVALID),
		.io_export_taskOut_9_TREADY(_peArray_9_taskIn_TREADY),
		.io_export_taskOut_9_TVALID(_Scheduler_io_export_taskOut_9_TVALID),
		.io_export_taskOut_10_TREADY(_peArray_10_taskIn_TREADY),
		.io_export_taskOut_10_TVALID(_Scheduler_io_export_taskOut_10_TVALID),
		.io_export_taskOut_11_TREADY(_peArray_11_taskIn_TREADY),
		.io_export_taskOut_11_TVALID(_Scheduler_io_export_taskOut_11_TVALID),
		.io_export_taskOut_12_TREADY(_peArray_12_taskIn_TREADY),
		.io_export_taskOut_12_TVALID(_Scheduler_io_export_taskOut_12_TVALID),
		.io_export_taskOut_13_TREADY(_peArray_13_taskIn_TREADY),
		.io_export_taskOut_13_TVALID(_Scheduler_io_export_taskOut_13_TVALID),
		.io_export_taskOut_14_TREADY(_peArray_14_taskIn_TREADY),
		.io_export_taskOut_14_TVALID(_Scheduler_io_export_taskOut_14_TVALID),
		.io_export_taskOut_15_TREADY(_peArray_15_taskIn_TREADY),
		.io_export_taskOut_15_TVALID(_Scheduler_io_export_taskOut_15_TVALID),
		.io_export_taskOut_16_TREADY(_peArray_16_taskIn_TREADY),
		.io_export_taskOut_16_TVALID(_Scheduler_io_export_taskOut_16_TVALID),
		.io_export_taskOut_17_TREADY(_peArray_17_taskIn_TREADY),
		.io_export_taskOut_17_TVALID(_Scheduler_io_export_taskOut_17_TVALID),
		.io_export_taskOut_18_TREADY(_peArray_18_taskIn_TREADY),
		.io_export_taskOut_18_TVALID(_Scheduler_io_export_taskOut_18_TVALID),
		.io_export_taskOut_19_TREADY(_peArray_19_taskIn_TREADY),
		.io_export_taskOut_19_TVALID(_Scheduler_io_export_taskOut_19_TVALID),
		.io_export_taskOut_20_TREADY(_peArray_20_taskIn_TREADY),
		.io_export_taskOut_20_TVALID(_Scheduler_io_export_taskOut_20_TVALID),
		.io_export_taskOut_21_TREADY(_peArray_21_taskIn_TREADY),
		.io_export_taskOut_21_TVALID(_Scheduler_io_export_taskOut_21_TVALID),
		.io_export_taskOut_22_TREADY(_peArray_22_taskIn_TREADY),
		.io_export_taskOut_22_TVALID(_Scheduler_io_export_taskOut_22_TVALID),
		.io_export_taskOut_23_TREADY(_peArray_23_taskIn_TREADY),
		.io_export_taskOut_23_TVALID(_Scheduler_io_export_taskOut_23_TVALID),
		.io_export_taskOut_24_TREADY(_peArray_24_taskIn_TREADY),
		.io_export_taskOut_24_TVALID(_Scheduler_io_export_taskOut_24_TVALID),
		.io_export_taskOut_25_TREADY(_peArray_25_taskIn_TREADY),
		.io_export_taskOut_25_TVALID(_Scheduler_io_export_taskOut_25_TVALID),
		.io_export_taskOut_26_TREADY(_peArray_26_taskIn_TREADY),
		.io_export_taskOut_26_TVALID(_Scheduler_io_export_taskOut_26_TVALID),
		.io_export_taskOut_27_TREADY(_peArray_27_taskIn_TREADY),
		.io_export_taskOut_27_TVALID(_Scheduler_io_export_taskOut_27_TVALID),
		.io_export_taskOut_28_TREADY(_peArray_28_taskIn_TREADY),
		.io_export_taskOut_28_TVALID(_Scheduler_io_export_taskOut_28_TVALID),
		.io_export_taskOut_29_TREADY(_peArray_29_taskIn_TREADY),
		.io_export_taskOut_29_TVALID(_Scheduler_io_export_taskOut_29_TVALID),
		.io_export_taskOut_30_TREADY(_peArray_30_taskIn_TREADY),
		.io_export_taskOut_30_TVALID(_Scheduler_io_export_taskOut_30_TVALID),
		.io_export_taskOut_31_TREADY(_peArray_31_taskIn_TREADY),
		.io_export_taskOut_31_TVALID(_Scheduler_io_export_taskOut_31_TVALID),
		.io_export_taskOut_32_TREADY(_peArray_32_taskIn_TREADY),
		.io_export_taskOut_32_TVALID(_Scheduler_io_export_taskOut_32_TVALID),
		.io_export_taskOut_33_TREADY(_peArray_33_taskIn_TREADY),
		.io_export_taskOut_33_TVALID(_Scheduler_io_export_taskOut_33_TVALID),
		.io_export_taskOut_34_TREADY(_peArray_34_taskIn_TREADY),
		.io_export_taskOut_34_TVALID(_Scheduler_io_export_taskOut_34_TVALID),
		.io_export_taskOut_35_TREADY(_peArray_35_taskIn_TREADY),
		.io_export_taskOut_35_TVALID(_Scheduler_io_export_taskOut_35_TVALID),
		.io_export_taskOut_36_TREADY(_peArray_36_taskIn_TREADY),
		.io_export_taskOut_36_TVALID(_Scheduler_io_export_taskOut_36_TVALID),
		.io_export_taskOut_37_TREADY(_peArray_37_taskIn_TREADY),
		.io_export_taskOut_37_TVALID(_Scheduler_io_export_taskOut_37_TVALID),
		.io_export_taskOut_38_TREADY(_peArray_38_taskIn_TREADY),
		.io_export_taskOut_38_TVALID(_Scheduler_io_export_taskOut_38_TVALID),
		.io_export_taskOut_39_TREADY(_peArray_39_taskIn_TREADY),
		.io_export_taskOut_39_TVALID(_Scheduler_io_export_taskOut_39_TVALID),
		.io_export_taskOut_40_TREADY(_peArray_40_taskIn_TREADY),
		.io_export_taskOut_40_TVALID(_Scheduler_io_export_taskOut_40_TVALID),
		.io_export_taskOut_41_TREADY(_peArray_41_taskIn_TREADY),
		.io_export_taskOut_41_TVALID(_Scheduler_io_export_taskOut_41_TVALID),
		.io_export_taskOut_42_TREADY(_peArray_42_taskIn_TREADY),
		.io_export_taskOut_42_TVALID(_Scheduler_io_export_taskOut_42_TVALID),
		.io_export_taskOut_43_TREADY(_peArray_43_taskIn_TREADY),
		.io_export_taskOut_43_TVALID(_Scheduler_io_export_taskOut_43_TVALID),
		.io_export_taskOut_44_TREADY(_peArray_44_taskIn_TREADY),
		.io_export_taskOut_44_TVALID(_Scheduler_io_export_taskOut_44_TVALID),
		.io_export_taskOut_45_TREADY(_peArray_45_taskIn_TREADY),
		.io_export_taskOut_45_TVALID(_Scheduler_io_export_taskOut_45_TVALID),
		.io_export_taskOut_46_TREADY(_peArray_46_taskIn_TREADY),
		.io_export_taskOut_46_TVALID(_Scheduler_io_export_taskOut_46_TVALID),
		.io_export_taskOut_47_TREADY(_peArray_47_taskIn_TREADY),
		.io_export_taskOut_47_TVALID(_Scheduler_io_export_taskOut_47_TVALID),
		.io_export_taskOut_48_TREADY(_peArray_48_taskIn_TREADY),
		.io_export_taskOut_48_TVALID(_Scheduler_io_export_taskOut_48_TVALID),
		.io_export_taskOut_49_TREADY(_peArray_49_taskIn_TREADY),
		.io_export_taskOut_49_TVALID(_Scheduler_io_export_taskOut_49_TVALID),
		.io_export_taskOut_50_TREADY(_peArray_50_taskIn_TREADY),
		.io_export_taskOut_50_TVALID(_Scheduler_io_export_taskOut_50_TVALID),
		.io_export_taskOut_51_TREADY(_peArray_51_taskIn_TREADY),
		.io_export_taskOut_51_TVALID(_Scheduler_io_export_taskOut_51_TVALID),
		.io_export_taskOut_52_TREADY(_peArray_52_taskIn_TREADY),
		.io_export_taskOut_52_TVALID(_Scheduler_io_export_taskOut_52_TVALID),
		.io_export_taskOut_53_TREADY(_peArray_53_taskIn_TREADY),
		.io_export_taskOut_53_TVALID(_Scheduler_io_export_taskOut_53_TVALID),
		.io_export_taskOut_54_TREADY(_peArray_54_taskIn_TREADY),
		.io_export_taskOut_54_TVALID(_Scheduler_io_export_taskOut_54_TVALID),
		.io_export_taskOut_55_TREADY(_peArray_55_taskIn_TREADY),
		.io_export_taskOut_55_TVALID(_Scheduler_io_export_taskOut_55_TVALID),
		.io_export_taskOut_56_TREADY(_peArray_56_taskIn_TREADY),
		.io_export_taskOut_56_TVALID(_Scheduler_io_export_taskOut_56_TVALID),
		.io_export_taskOut_57_TREADY(_peArray_57_taskIn_TREADY),
		.io_export_taskOut_57_TVALID(_Scheduler_io_export_taskOut_57_TVALID),
		.io_export_taskOut_58_TREADY(_peArray_58_taskIn_TREADY),
		.io_export_taskOut_58_TVALID(_Scheduler_io_export_taskOut_58_TVALID),
		.io_export_taskOut_59_TREADY(_peArray_59_taskIn_TREADY),
		.io_export_taskOut_59_TVALID(_Scheduler_io_export_taskOut_59_TVALID),
		.io_export_taskOut_60_TREADY(_peArray_60_taskIn_TREADY),
		.io_export_taskOut_60_TVALID(_Scheduler_io_export_taskOut_60_TVALID),
		.io_export_taskOut_61_TREADY(_peArray_61_taskIn_TREADY),
		.io_export_taskOut_61_TVALID(_Scheduler_io_export_taskOut_61_TVALID),
		.io_export_taskOut_62_TREADY(_peArray_62_taskIn_TREADY),
		.io_export_taskOut_62_TVALID(_Scheduler_io_export_taskOut_62_TVALID),
		.io_export_taskOut_63_TREADY(_peArray_63_taskIn_TREADY),
		.io_export_taskOut_63_TVALID(_Scheduler_io_export_taskOut_63_TVALID),
		.io_export_taskIn_0_TREADY(_Scheduler_io_export_taskIn_0_TREADY),
		.io_export_taskIn_0_TVALID(_peArray_0_taskOut_TVALID),
		.io_export_taskIn_0_TDATA(_peArray_0_taskOut_TDATA[31:0]),
		.io_export_taskIn_1_TREADY(_Scheduler_io_export_taskIn_1_TREADY),
		.io_export_taskIn_1_TVALID(_peArray_1_taskOut_TVALID),
		.io_export_taskIn_1_TDATA(_peArray_1_taskOut_TDATA[31:0]),
		.io_export_taskIn_2_TREADY(_Scheduler_io_export_taskIn_2_TREADY),
		.io_export_taskIn_2_TVALID(_peArray_2_taskOut_TVALID),
		.io_export_taskIn_2_TDATA(_peArray_2_taskOut_TDATA[31:0]),
		.io_export_taskIn_3_TREADY(_Scheduler_io_export_taskIn_3_TREADY),
		.io_export_taskIn_3_TVALID(_peArray_3_taskOut_TVALID),
		.io_export_taskIn_3_TDATA(_peArray_3_taskOut_TDATA[31:0]),
		.io_export_taskIn_4_TREADY(_Scheduler_io_export_taskIn_4_TREADY),
		.io_export_taskIn_4_TVALID(_peArray_4_taskOut_TVALID),
		.io_export_taskIn_4_TDATA(_peArray_4_taskOut_TDATA[31:0]),
		.io_export_taskIn_5_TREADY(_Scheduler_io_export_taskIn_5_TREADY),
		.io_export_taskIn_5_TVALID(_peArray_5_taskOut_TVALID),
		.io_export_taskIn_5_TDATA(_peArray_5_taskOut_TDATA[31:0]),
		.io_export_taskIn_6_TREADY(_Scheduler_io_export_taskIn_6_TREADY),
		.io_export_taskIn_6_TVALID(_peArray_6_taskOut_TVALID),
		.io_export_taskIn_6_TDATA(_peArray_6_taskOut_TDATA[31:0]),
		.io_export_taskIn_7_TREADY(_Scheduler_io_export_taskIn_7_TREADY),
		.io_export_taskIn_7_TVALID(_peArray_7_taskOut_TVALID),
		.io_export_taskIn_7_TDATA(_peArray_7_taskOut_TDATA[31:0]),
		.io_export_taskIn_8_TREADY(_Scheduler_io_export_taskIn_8_TREADY),
		.io_export_taskIn_8_TVALID(_peArray_8_taskOut_TVALID),
		.io_export_taskIn_8_TDATA(_peArray_8_taskOut_TDATA[31:0]),
		.io_export_taskIn_9_TREADY(_Scheduler_io_export_taskIn_9_TREADY),
		.io_export_taskIn_9_TVALID(_peArray_9_taskOut_TVALID),
		.io_export_taskIn_9_TDATA(_peArray_9_taskOut_TDATA[31:0]),
		.io_export_taskIn_10_TREADY(_Scheduler_io_export_taskIn_10_TREADY),
		.io_export_taskIn_10_TVALID(_peArray_10_taskOut_TVALID),
		.io_export_taskIn_10_TDATA(_peArray_10_taskOut_TDATA[31:0]),
		.io_export_taskIn_11_TREADY(_Scheduler_io_export_taskIn_11_TREADY),
		.io_export_taskIn_11_TVALID(_peArray_11_taskOut_TVALID),
		.io_export_taskIn_11_TDATA(_peArray_11_taskOut_TDATA[31:0]),
		.io_export_taskIn_12_TREADY(_Scheduler_io_export_taskIn_12_TREADY),
		.io_export_taskIn_12_TVALID(_peArray_12_taskOut_TVALID),
		.io_export_taskIn_12_TDATA(_peArray_12_taskOut_TDATA[31:0]),
		.io_export_taskIn_13_TREADY(_Scheduler_io_export_taskIn_13_TREADY),
		.io_export_taskIn_13_TVALID(_peArray_13_taskOut_TVALID),
		.io_export_taskIn_13_TDATA(_peArray_13_taskOut_TDATA[31:0]),
		.io_export_taskIn_14_TREADY(_Scheduler_io_export_taskIn_14_TREADY),
		.io_export_taskIn_14_TVALID(_peArray_14_taskOut_TVALID),
		.io_export_taskIn_14_TDATA(_peArray_14_taskOut_TDATA[31:0]),
		.io_export_taskIn_15_TREADY(_Scheduler_io_export_taskIn_15_TREADY),
		.io_export_taskIn_15_TVALID(_peArray_15_taskOut_TVALID),
		.io_export_taskIn_15_TDATA(_peArray_15_taskOut_TDATA[31:0]),
		.io_export_taskIn_16_TREADY(_Scheduler_io_export_taskIn_16_TREADY),
		.io_export_taskIn_16_TVALID(_peArray_16_taskOut_TVALID),
		.io_export_taskIn_16_TDATA(_peArray_16_taskOut_TDATA[31:0]),
		.io_export_taskIn_17_TREADY(_Scheduler_io_export_taskIn_17_TREADY),
		.io_export_taskIn_17_TVALID(_peArray_17_taskOut_TVALID),
		.io_export_taskIn_17_TDATA(_peArray_17_taskOut_TDATA[31:0]),
		.io_export_taskIn_18_TREADY(_Scheduler_io_export_taskIn_18_TREADY),
		.io_export_taskIn_18_TVALID(_peArray_18_taskOut_TVALID),
		.io_export_taskIn_18_TDATA(_peArray_18_taskOut_TDATA[31:0]),
		.io_export_taskIn_19_TREADY(_Scheduler_io_export_taskIn_19_TREADY),
		.io_export_taskIn_19_TVALID(_peArray_19_taskOut_TVALID),
		.io_export_taskIn_19_TDATA(_peArray_19_taskOut_TDATA[31:0]),
		.io_export_taskIn_20_TREADY(_Scheduler_io_export_taskIn_20_TREADY),
		.io_export_taskIn_20_TVALID(_peArray_20_taskOut_TVALID),
		.io_export_taskIn_20_TDATA(_peArray_20_taskOut_TDATA[31:0]),
		.io_export_taskIn_21_TREADY(_Scheduler_io_export_taskIn_21_TREADY),
		.io_export_taskIn_21_TVALID(_peArray_21_taskOut_TVALID),
		.io_export_taskIn_21_TDATA(_peArray_21_taskOut_TDATA[31:0]),
		.io_export_taskIn_22_TREADY(_Scheduler_io_export_taskIn_22_TREADY),
		.io_export_taskIn_22_TVALID(_peArray_22_taskOut_TVALID),
		.io_export_taskIn_22_TDATA(_peArray_22_taskOut_TDATA[31:0]),
		.io_export_taskIn_23_TREADY(_Scheduler_io_export_taskIn_23_TREADY),
		.io_export_taskIn_23_TVALID(_peArray_23_taskOut_TVALID),
		.io_export_taskIn_23_TDATA(_peArray_23_taskOut_TDATA[31:0]),
		.io_export_taskIn_24_TREADY(_Scheduler_io_export_taskIn_24_TREADY),
		.io_export_taskIn_24_TVALID(_peArray_24_taskOut_TVALID),
		.io_export_taskIn_24_TDATA(_peArray_24_taskOut_TDATA[31:0]),
		.io_export_taskIn_25_TREADY(_Scheduler_io_export_taskIn_25_TREADY),
		.io_export_taskIn_25_TVALID(_peArray_25_taskOut_TVALID),
		.io_export_taskIn_25_TDATA(_peArray_25_taskOut_TDATA[31:0]),
		.io_export_taskIn_26_TREADY(_Scheduler_io_export_taskIn_26_TREADY),
		.io_export_taskIn_26_TVALID(_peArray_26_taskOut_TVALID),
		.io_export_taskIn_26_TDATA(_peArray_26_taskOut_TDATA[31:0]),
		.io_export_taskIn_27_TREADY(_Scheduler_io_export_taskIn_27_TREADY),
		.io_export_taskIn_27_TVALID(_peArray_27_taskOut_TVALID),
		.io_export_taskIn_27_TDATA(_peArray_27_taskOut_TDATA[31:0]),
		.io_export_taskIn_28_TREADY(_Scheduler_io_export_taskIn_28_TREADY),
		.io_export_taskIn_28_TVALID(_peArray_28_taskOut_TVALID),
		.io_export_taskIn_28_TDATA(_peArray_28_taskOut_TDATA[31:0]),
		.io_export_taskIn_29_TREADY(_Scheduler_io_export_taskIn_29_TREADY),
		.io_export_taskIn_29_TVALID(_peArray_29_taskOut_TVALID),
		.io_export_taskIn_29_TDATA(_peArray_29_taskOut_TDATA[31:0]),
		.io_export_taskIn_30_TREADY(_Scheduler_io_export_taskIn_30_TREADY),
		.io_export_taskIn_30_TVALID(_peArray_30_taskOut_TVALID),
		.io_export_taskIn_30_TDATA(_peArray_30_taskOut_TDATA[31:0]),
		.io_export_taskIn_31_TREADY(_Scheduler_io_export_taskIn_31_TREADY),
		.io_export_taskIn_31_TVALID(_peArray_31_taskOut_TVALID),
		.io_export_taskIn_31_TDATA(_peArray_31_taskOut_TDATA[31:0]),
		.io_export_taskIn_32_TREADY(_Scheduler_io_export_taskIn_32_TREADY),
		.io_export_taskIn_32_TVALID(_peArray_32_taskOut_TVALID),
		.io_export_taskIn_32_TDATA(_peArray_32_taskOut_TDATA[31:0]),
		.io_export_taskIn_33_TREADY(_Scheduler_io_export_taskIn_33_TREADY),
		.io_export_taskIn_33_TVALID(_peArray_33_taskOut_TVALID),
		.io_export_taskIn_33_TDATA(_peArray_33_taskOut_TDATA[31:0]),
		.io_export_taskIn_34_TREADY(_Scheduler_io_export_taskIn_34_TREADY),
		.io_export_taskIn_34_TVALID(_peArray_34_taskOut_TVALID),
		.io_export_taskIn_34_TDATA(_peArray_34_taskOut_TDATA[31:0]),
		.io_export_taskIn_35_TREADY(_Scheduler_io_export_taskIn_35_TREADY),
		.io_export_taskIn_35_TVALID(_peArray_35_taskOut_TVALID),
		.io_export_taskIn_35_TDATA(_peArray_35_taskOut_TDATA[31:0]),
		.io_export_taskIn_36_TREADY(_Scheduler_io_export_taskIn_36_TREADY),
		.io_export_taskIn_36_TVALID(_peArray_36_taskOut_TVALID),
		.io_export_taskIn_36_TDATA(_peArray_36_taskOut_TDATA[31:0]),
		.io_export_taskIn_37_TREADY(_Scheduler_io_export_taskIn_37_TREADY),
		.io_export_taskIn_37_TVALID(_peArray_37_taskOut_TVALID),
		.io_export_taskIn_37_TDATA(_peArray_37_taskOut_TDATA[31:0]),
		.io_export_taskIn_38_TREADY(_Scheduler_io_export_taskIn_38_TREADY),
		.io_export_taskIn_38_TVALID(_peArray_38_taskOut_TVALID),
		.io_export_taskIn_38_TDATA(_peArray_38_taskOut_TDATA[31:0]),
		.io_export_taskIn_39_TREADY(_Scheduler_io_export_taskIn_39_TREADY),
		.io_export_taskIn_39_TVALID(_peArray_39_taskOut_TVALID),
		.io_export_taskIn_39_TDATA(_peArray_39_taskOut_TDATA[31:0]),
		.io_export_taskIn_40_TREADY(_Scheduler_io_export_taskIn_40_TREADY),
		.io_export_taskIn_40_TVALID(_peArray_40_taskOut_TVALID),
		.io_export_taskIn_40_TDATA(_peArray_40_taskOut_TDATA[31:0]),
		.io_export_taskIn_41_TREADY(_Scheduler_io_export_taskIn_41_TREADY),
		.io_export_taskIn_41_TVALID(_peArray_41_taskOut_TVALID),
		.io_export_taskIn_41_TDATA(_peArray_41_taskOut_TDATA[31:0]),
		.io_export_taskIn_42_TREADY(_Scheduler_io_export_taskIn_42_TREADY),
		.io_export_taskIn_42_TVALID(_peArray_42_taskOut_TVALID),
		.io_export_taskIn_42_TDATA(_peArray_42_taskOut_TDATA[31:0]),
		.io_export_taskIn_43_TREADY(_Scheduler_io_export_taskIn_43_TREADY),
		.io_export_taskIn_43_TVALID(_peArray_43_taskOut_TVALID),
		.io_export_taskIn_43_TDATA(_peArray_43_taskOut_TDATA[31:0]),
		.io_export_taskIn_44_TREADY(_Scheduler_io_export_taskIn_44_TREADY),
		.io_export_taskIn_44_TVALID(_peArray_44_taskOut_TVALID),
		.io_export_taskIn_44_TDATA(_peArray_44_taskOut_TDATA[31:0]),
		.io_export_taskIn_45_TREADY(_Scheduler_io_export_taskIn_45_TREADY),
		.io_export_taskIn_45_TVALID(_peArray_45_taskOut_TVALID),
		.io_export_taskIn_45_TDATA(_peArray_45_taskOut_TDATA[31:0]),
		.io_export_taskIn_46_TREADY(_Scheduler_io_export_taskIn_46_TREADY),
		.io_export_taskIn_46_TVALID(_peArray_46_taskOut_TVALID),
		.io_export_taskIn_46_TDATA(_peArray_46_taskOut_TDATA[31:0]),
		.io_export_taskIn_47_TREADY(_Scheduler_io_export_taskIn_47_TREADY),
		.io_export_taskIn_47_TVALID(_peArray_47_taskOut_TVALID),
		.io_export_taskIn_47_TDATA(_peArray_47_taskOut_TDATA[31:0]),
		.io_export_taskIn_48_TREADY(_Scheduler_io_export_taskIn_48_TREADY),
		.io_export_taskIn_48_TVALID(_peArray_48_taskOut_TVALID),
		.io_export_taskIn_48_TDATA(_peArray_48_taskOut_TDATA[31:0]),
		.io_export_taskIn_49_TREADY(_Scheduler_io_export_taskIn_49_TREADY),
		.io_export_taskIn_49_TVALID(_peArray_49_taskOut_TVALID),
		.io_export_taskIn_49_TDATA(_peArray_49_taskOut_TDATA[31:0]),
		.io_export_taskIn_50_TREADY(_Scheduler_io_export_taskIn_50_TREADY),
		.io_export_taskIn_50_TVALID(_peArray_50_taskOut_TVALID),
		.io_export_taskIn_50_TDATA(_peArray_50_taskOut_TDATA[31:0]),
		.io_export_taskIn_51_TREADY(_Scheduler_io_export_taskIn_51_TREADY),
		.io_export_taskIn_51_TVALID(_peArray_51_taskOut_TVALID),
		.io_export_taskIn_51_TDATA(_peArray_51_taskOut_TDATA[31:0]),
		.io_export_taskIn_52_TREADY(_Scheduler_io_export_taskIn_52_TREADY),
		.io_export_taskIn_52_TVALID(_peArray_52_taskOut_TVALID),
		.io_export_taskIn_52_TDATA(_peArray_52_taskOut_TDATA[31:0]),
		.io_export_taskIn_53_TREADY(_Scheduler_io_export_taskIn_53_TREADY),
		.io_export_taskIn_53_TVALID(_peArray_53_taskOut_TVALID),
		.io_export_taskIn_53_TDATA(_peArray_53_taskOut_TDATA[31:0]),
		.io_export_taskIn_54_TREADY(_Scheduler_io_export_taskIn_54_TREADY),
		.io_export_taskIn_54_TVALID(_peArray_54_taskOut_TVALID),
		.io_export_taskIn_54_TDATA(_peArray_54_taskOut_TDATA[31:0]),
		.io_export_taskIn_55_TREADY(_Scheduler_io_export_taskIn_55_TREADY),
		.io_export_taskIn_55_TVALID(_peArray_55_taskOut_TVALID),
		.io_export_taskIn_55_TDATA(_peArray_55_taskOut_TDATA[31:0]),
		.io_export_taskIn_56_TREADY(_Scheduler_io_export_taskIn_56_TREADY),
		.io_export_taskIn_56_TVALID(_peArray_56_taskOut_TVALID),
		.io_export_taskIn_56_TDATA(_peArray_56_taskOut_TDATA[31:0]),
		.io_export_taskIn_57_TREADY(_Scheduler_io_export_taskIn_57_TREADY),
		.io_export_taskIn_57_TVALID(_peArray_57_taskOut_TVALID),
		.io_export_taskIn_57_TDATA(_peArray_57_taskOut_TDATA[31:0]),
		.io_export_taskIn_58_TREADY(_Scheduler_io_export_taskIn_58_TREADY),
		.io_export_taskIn_58_TVALID(_peArray_58_taskOut_TVALID),
		.io_export_taskIn_58_TDATA(_peArray_58_taskOut_TDATA[31:0]),
		.io_export_taskIn_59_TREADY(_Scheduler_io_export_taskIn_59_TREADY),
		.io_export_taskIn_59_TVALID(_peArray_59_taskOut_TVALID),
		.io_export_taskIn_59_TDATA(_peArray_59_taskOut_TDATA[31:0]),
		.io_export_taskIn_60_TREADY(_Scheduler_io_export_taskIn_60_TREADY),
		.io_export_taskIn_60_TVALID(_peArray_60_taskOut_TVALID),
		.io_export_taskIn_60_TDATA(_peArray_60_taskOut_TDATA[31:0]),
		.io_export_taskIn_61_TREADY(_Scheduler_io_export_taskIn_61_TREADY),
		.io_export_taskIn_61_TVALID(_peArray_61_taskOut_TVALID),
		.io_export_taskIn_61_TDATA(_peArray_61_taskOut_TDATA[31:0]),
		.io_export_taskIn_62_TREADY(_Scheduler_io_export_taskIn_62_TREADY),
		.io_export_taskIn_62_TVALID(_peArray_62_taskOut_TVALID),
		.io_export_taskIn_62_TDATA(_peArray_62_taskOut_TDATA[31:0]),
		.io_export_taskIn_63_TREADY(_Scheduler_io_export_taskIn_63_TREADY),
		.io_export_taskIn_63_TVALID(_peArray_63_taskOut_TVALID),
		.io_export_taskIn_63_TDATA(_peArray_63_taskOut_TDATA[31:0]),
		.io_internal_vss_axi_full_0_ar_ready(qsort_schedulerAXI_0_ARREADY),
		.io_internal_vss_axi_full_0_ar_valid(qsort_schedulerAXI_0_ARVALID),
		.io_internal_vss_axi_full_0_ar_bits_addr(qsort_schedulerAXI_0_ARADDR),
		.io_internal_vss_axi_full_0_ar_bits_len(qsort_schedulerAXI_0_ARLEN),
		.io_internal_vss_axi_full_0_ar_bits_size(qsort_schedulerAXI_0_ARSIZE),
		.io_internal_vss_axi_full_0_ar_bits_burst(qsort_schedulerAXI_0_ARBURST),
		.io_internal_vss_axi_full_0_ar_bits_lock(qsort_schedulerAXI_0_ARLOCK),
		.io_internal_vss_axi_full_0_ar_bits_cache(qsort_schedulerAXI_0_ARCACHE),
		.io_internal_vss_axi_full_0_ar_bits_prot(qsort_schedulerAXI_0_ARPROT),
		.io_internal_vss_axi_full_0_ar_bits_qos(qsort_schedulerAXI_0_ARQOS),
		.io_internal_vss_axi_full_0_ar_bits_region(qsort_schedulerAXI_0_ARREGION),
		.io_internal_vss_axi_full_0_r_ready(qsort_schedulerAXI_0_RREADY),
		.io_internal_vss_axi_full_0_r_valid(qsort_schedulerAXI_0_RVALID),
		.io_internal_vss_axi_full_0_r_bits_data(qsort_schedulerAXI_0_RDATA),
		.io_internal_vss_axi_full_0_aw_ready(qsort_schedulerAXI_0_AWREADY),
		.io_internal_vss_axi_full_0_aw_valid(qsort_schedulerAXI_0_AWVALID),
		.io_internal_vss_axi_full_0_aw_bits_addr(qsort_schedulerAXI_0_AWADDR),
		.io_internal_vss_axi_full_0_aw_bits_len(qsort_schedulerAXI_0_AWLEN),
		.io_internal_vss_axi_full_0_aw_bits_size(qsort_schedulerAXI_0_AWSIZE),
		.io_internal_vss_axi_full_0_aw_bits_burst(qsort_schedulerAXI_0_AWBURST),
		.io_internal_vss_axi_full_0_aw_bits_lock(qsort_schedulerAXI_0_AWLOCK),
		.io_internal_vss_axi_full_0_aw_bits_cache(qsort_schedulerAXI_0_AWCACHE),
		.io_internal_vss_axi_full_0_aw_bits_prot(qsort_schedulerAXI_0_AWPROT),
		.io_internal_vss_axi_full_0_aw_bits_qos(qsort_schedulerAXI_0_AWQOS),
		.io_internal_vss_axi_full_0_aw_bits_region(qsort_schedulerAXI_0_AWREGION),
		.io_internal_vss_axi_full_0_w_ready(qsort_schedulerAXI_0_WREADY),
		.io_internal_vss_axi_full_0_w_valid(qsort_schedulerAXI_0_WVALID),
		.io_internal_vss_axi_full_0_w_bits_data(qsort_schedulerAXI_0_WDATA),
		.io_internal_vss_axi_full_0_w_bits_last(qsort_schedulerAXI_0_WLAST),
		.io_internal_vss_axi_full_0_b_valid(qsort_schedulerAXI_0_BVALID),
		.io_internal_axi_mgmt_vss_0_ar_ready(_Scheduler_io_internal_axi_mgmt_vss_0_ar_ready),
		.io_internal_axi_mgmt_vss_0_ar_valid(_demux_m_axil_0_ar_valid),
		.io_internal_axi_mgmt_vss_0_ar_bits_addr(_demux_m_axil_0_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_ar_bits_prot(_demux_m_axil_0_ar_bits_prot),
		.io_internal_axi_mgmt_vss_0_r_ready(_demux_m_axil_0_r_ready),
		.io_internal_axi_mgmt_vss_0_r_valid(_Scheduler_io_internal_axi_mgmt_vss_0_r_valid),
		.io_internal_axi_mgmt_vss_0_r_bits_data(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_internal_axi_mgmt_vss_0_r_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_internal_axi_mgmt_vss_0_aw_ready(_Scheduler_io_internal_axi_mgmt_vss_0_aw_ready),
		.io_internal_axi_mgmt_vss_0_aw_valid(_demux_m_axil_0_aw_valid),
		.io_internal_axi_mgmt_vss_0_aw_bits_addr(_demux_m_axil_0_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_aw_bits_prot(_demux_m_axil_0_aw_bits_prot),
		.io_internal_axi_mgmt_vss_0_w_ready(_Scheduler_io_internal_axi_mgmt_vss_0_w_ready),
		.io_internal_axi_mgmt_vss_0_w_valid(_demux_m_axil_0_w_valid),
		.io_internal_axi_mgmt_vss_0_w_bits_data(_demux_m_axil_0_w_bits_data),
		.io_internal_axi_mgmt_vss_0_w_bits_strb(_demux_m_axil_0_w_bits_strb),
		.io_internal_axi_mgmt_vss_0_b_ready(_demux_m_axil_0_b_ready),
		.io_internal_axi_mgmt_vss_0_b_valid(_Scheduler_io_internal_axi_mgmt_vss_0_b_valid),
		.io_internal_axi_mgmt_vss_0_b_bits_resp(_Scheduler_io_internal_axi_mgmt_vss_0_b_bits_resp)
	);
	sync peArray_0_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_64_TREADY),
		.argOut_TVALID(_peArray_0_1_argOut_TVALID),
		.argOut_TDATA(_peArray_0_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_0_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_0_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_1_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_65_TREADY),
		.argOut_TVALID(_peArray_1_1_argOut_TVALID),
		.argOut_TDATA(_peArray_1_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_1_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_1_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_2_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_66_TREADY),
		.argOut_TVALID(_peArray_2_1_argOut_TVALID),
		.argOut_TDATA(_peArray_2_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_2_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_2_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_3_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_67_TREADY),
		.argOut_TVALID(_peArray_3_1_argOut_TVALID),
		.argOut_TDATA(_peArray_3_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_3_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_3_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_4_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_68_TREADY),
		.argOut_TVALID(_peArray_4_1_argOut_TVALID),
		.argOut_TDATA(_peArray_4_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_4_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_4_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_5_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_69_TREADY),
		.argOut_TVALID(_peArray_5_1_argOut_TVALID),
		.argOut_TDATA(_peArray_5_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_5_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_5_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_6_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_70_TREADY),
		.argOut_TVALID(_peArray_6_1_argOut_TVALID),
		.argOut_TDATA(_peArray_6_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_6_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_6_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_7_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_71_TREADY),
		.argOut_TVALID(_peArray_7_1_argOut_TVALID),
		.argOut_TDATA(_peArray_7_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_7_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_7_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_8_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_72_TREADY),
		.argOut_TVALID(_peArray_8_1_argOut_TVALID),
		.argOut_TDATA(_peArray_8_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_8_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_8_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_9_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_73_TREADY),
		.argOut_TVALID(_peArray_9_1_argOut_TVALID),
		.argOut_TDATA(_peArray_9_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_9_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_9_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_10_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_74_TREADY),
		.argOut_TVALID(_peArray_10_1_argOut_TVALID),
		.argOut_TDATA(_peArray_10_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_10_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_10_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_11_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_75_TREADY),
		.argOut_TVALID(_peArray_11_1_argOut_TVALID),
		.argOut_TDATA(_peArray_11_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_11_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_11_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_12_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_76_TREADY),
		.argOut_TVALID(_peArray_12_1_argOut_TVALID),
		.argOut_TDATA(_peArray_12_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_12_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_12_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_13_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_77_TREADY),
		.argOut_TVALID(_peArray_13_1_argOut_TVALID),
		.argOut_TDATA(_peArray_13_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_13_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_13_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_14_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_78_TREADY),
		.argOut_TVALID(_peArray_14_1_argOut_TVALID),
		.argOut_TDATA(_peArray_14_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_14_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_14_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	sync peArray_15_1(
		.ap_rst_n(~reset),
		.ap_clk(clock),
		.argOut_TREADY(_ArgumentNotifier_io_export_argIn_79_TREADY),
		.argOut_TVALID(_peArray_15_1_argOut_TVALID),
		.argOut_TDATA(_peArray_15_1_argOut_TDATA),
		.taskIn_TREADY(_peArray_15_1_taskIn_TREADY),
		.taskIn_TVALID(_Scheduler_1_io_export_taskOut_15_TVALID),
		.taskIn_TDATA(128'h00000000000000000000000000000000)
	);
	Scheduler_1 Scheduler_1(
		.clock(clock),
		.reset(reset),
		.io_export_taskOut_0_TREADY(_peArray_0_1_taskIn_TREADY),
		.io_export_taskOut_0_TVALID(_Scheduler_1_io_export_taskOut_0_TVALID),
		.io_export_taskOut_1_TREADY(_peArray_1_1_taskIn_TREADY),
		.io_export_taskOut_1_TVALID(_Scheduler_1_io_export_taskOut_1_TVALID),
		.io_export_taskOut_2_TREADY(_peArray_2_1_taskIn_TREADY),
		.io_export_taskOut_2_TVALID(_Scheduler_1_io_export_taskOut_2_TVALID),
		.io_export_taskOut_3_TREADY(_peArray_3_1_taskIn_TREADY),
		.io_export_taskOut_3_TVALID(_Scheduler_1_io_export_taskOut_3_TVALID),
		.io_export_taskOut_4_TREADY(_peArray_4_1_taskIn_TREADY),
		.io_export_taskOut_4_TVALID(_Scheduler_1_io_export_taskOut_4_TVALID),
		.io_export_taskOut_5_TREADY(_peArray_5_1_taskIn_TREADY),
		.io_export_taskOut_5_TVALID(_Scheduler_1_io_export_taskOut_5_TVALID),
		.io_export_taskOut_6_TREADY(_peArray_6_1_taskIn_TREADY),
		.io_export_taskOut_6_TVALID(_Scheduler_1_io_export_taskOut_6_TVALID),
		.io_export_taskOut_7_TREADY(_peArray_7_1_taskIn_TREADY),
		.io_export_taskOut_7_TVALID(_Scheduler_1_io_export_taskOut_7_TVALID),
		.io_export_taskOut_8_TREADY(_peArray_8_1_taskIn_TREADY),
		.io_export_taskOut_8_TVALID(_Scheduler_1_io_export_taskOut_8_TVALID),
		.io_export_taskOut_9_TREADY(_peArray_9_1_taskIn_TREADY),
		.io_export_taskOut_9_TVALID(_Scheduler_1_io_export_taskOut_9_TVALID),
		.io_export_taskOut_10_TREADY(_peArray_10_1_taskIn_TREADY),
		.io_export_taskOut_10_TVALID(_Scheduler_1_io_export_taskOut_10_TVALID),
		.io_export_taskOut_11_TREADY(_peArray_11_1_taskIn_TREADY),
		.io_export_taskOut_11_TVALID(_Scheduler_1_io_export_taskOut_11_TVALID),
		.io_export_taskOut_12_TREADY(_peArray_12_1_taskIn_TREADY),
		.io_export_taskOut_12_TVALID(_Scheduler_1_io_export_taskOut_12_TVALID),
		.io_export_taskOut_13_TREADY(_peArray_13_1_taskIn_TREADY),
		.io_export_taskOut_13_TVALID(_Scheduler_1_io_export_taskOut_13_TVALID),
		.io_export_taskOut_14_TREADY(_peArray_14_1_taskIn_TREADY),
		.io_export_taskOut_14_TVALID(_Scheduler_1_io_export_taskOut_14_TVALID),
		.io_export_taskOut_15_TREADY(_peArray_15_1_taskIn_TREADY),
		.io_export_taskOut_15_TVALID(_Scheduler_1_io_export_taskOut_15_TVALID),
		.io_internal_vss_axi_full_0_ar_ready(sync_schedulerAXI_0_ARREADY),
		.io_internal_vss_axi_full_0_ar_valid(sync_schedulerAXI_0_ARVALID),
		.io_internal_vss_axi_full_0_ar_bits_addr(sync_schedulerAXI_0_ARADDR),
		.io_internal_vss_axi_full_0_ar_bits_len(sync_schedulerAXI_0_ARLEN),
		.io_internal_vss_axi_full_0_ar_bits_size(sync_schedulerAXI_0_ARSIZE),
		.io_internal_vss_axi_full_0_ar_bits_burst(sync_schedulerAXI_0_ARBURST),
		.io_internal_vss_axi_full_0_ar_bits_lock(sync_schedulerAXI_0_ARLOCK),
		.io_internal_vss_axi_full_0_ar_bits_cache(sync_schedulerAXI_0_ARCACHE),
		.io_internal_vss_axi_full_0_ar_bits_prot(sync_schedulerAXI_0_ARPROT),
		.io_internal_vss_axi_full_0_ar_bits_qos(sync_schedulerAXI_0_ARQOS),
		.io_internal_vss_axi_full_0_ar_bits_region(sync_schedulerAXI_0_ARREGION),
		.io_internal_vss_axi_full_0_r_ready(sync_schedulerAXI_0_RREADY),
		.io_internal_vss_axi_full_0_r_valid(sync_schedulerAXI_0_RVALID),
		.io_internal_vss_axi_full_0_r_bits_data(sync_schedulerAXI_0_RDATA),
		.io_internal_vss_axi_full_0_aw_ready(sync_schedulerAXI_0_AWREADY),
		.io_internal_vss_axi_full_0_aw_valid(sync_schedulerAXI_0_AWVALID),
		.io_internal_vss_axi_full_0_aw_bits_addr(sync_schedulerAXI_0_AWADDR),
		.io_internal_vss_axi_full_0_aw_bits_len(sync_schedulerAXI_0_AWLEN),
		.io_internal_vss_axi_full_0_aw_bits_size(sync_schedulerAXI_0_AWSIZE),
		.io_internal_vss_axi_full_0_aw_bits_burst(sync_schedulerAXI_0_AWBURST),
		.io_internal_vss_axi_full_0_aw_bits_lock(sync_schedulerAXI_0_AWLOCK),
		.io_internal_vss_axi_full_0_aw_bits_cache(sync_schedulerAXI_0_AWCACHE),
		.io_internal_vss_axi_full_0_aw_bits_prot(sync_schedulerAXI_0_AWPROT),
		.io_internal_vss_axi_full_0_aw_bits_qos(sync_schedulerAXI_0_AWQOS),
		.io_internal_vss_axi_full_0_aw_bits_region(sync_schedulerAXI_0_AWREGION),
		.io_internal_vss_axi_full_0_w_ready(sync_schedulerAXI_0_WREADY),
		.io_internal_vss_axi_full_0_w_valid(sync_schedulerAXI_0_WVALID),
		.io_internal_vss_axi_full_0_w_bits_data(sync_schedulerAXI_0_WDATA),
		.io_internal_vss_axi_full_0_w_bits_last(sync_schedulerAXI_0_WLAST),
		.io_internal_vss_axi_full_0_b_valid(sync_schedulerAXI_0_BVALID),
		.io_internal_axi_mgmt_vss_0_ar_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_ar_ready),
		.io_internal_axi_mgmt_vss_0_ar_valid(_demux_m_axil_1_ar_valid),
		.io_internal_axi_mgmt_vss_0_ar_bits_addr(_demux_m_axil_1_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_ar_bits_prot(_demux_m_axil_1_ar_bits_prot),
		.io_internal_axi_mgmt_vss_0_r_ready(_demux_m_axil_1_r_ready),
		.io_internal_axi_mgmt_vss_0_r_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_valid),
		.io_internal_axi_mgmt_vss_0_r_bits_data(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_data),
		.io_internal_axi_mgmt_vss_0_r_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_r_bits_resp),
		.io_internal_axi_mgmt_vss_0_aw_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_aw_ready),
		.io_internal_axi_mgmt_vss_0_aw_valid(_demux_m_axil_1_aw_valid),
		.io_internal_axi_mgmt_vss_0_aw_bits_addr(_demux_m_axil_1_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vss_0_aw_bits_prot(_demux_m_axil_1_aw_bits_prot),
		.io_internal_axi_mgmt_vss_0_w_ready(_Scheduler_1_io_internal_axi_mgmt_vss_0_w_ready),
		.io_internal_axi_mgmt_vss_0_w_valid(_demux_m_axil_1_w_valid),
		.io_internal_axi_mgmt_vss_0_w_bits_data(_demux_m_axil_1_w_bits_data),
		.io_internal_axi_mgmt_vss_0_w_bits_strb(_demux_m_axil_1_w_bits_strb),
		.io_internal_axi_mgmt_vss_0_b_ready(_demux_m_axil_1_b_ready),
		.io_internal_axi_mgmt_vss_0_b_valid(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_valid),
		.io_internal_axi_mgmt_vss_0_b_bits_resp(_Scheduler_1_io_internal_axi_mgmt_vss_0_b_bits_resp),
		.connArgumentNotifier_0_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_0_ctrl_serveStealReq_valid),
		.connArgumentNotifier_0_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_0_ctrl_serveStealReq_ready),
		.connArgumentNotifier_0_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_0_data_qOutTask_ready),
		.connArgumentNotifier_0_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_0_data_qOutTask_valid),
		.connArgumentNotifier_0_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_0_data_qOutTask_bits),
		.connArgumentNotifier_1_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_1_ctrl_serveStealReq_valid),
		.connArgumentNotifier_1_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_1_ctrl_serveStealReq_ready),
		.connArgumentNotifier_1_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_1_data_qOutTask_ready),
		.connArgumentNotifier_1_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_1_data_qOutTask_valid),
		.connArgumentNotifier_1_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_1_data_qOutTask_bits),
		.connArgumentNotifier_2_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_2_ctrl_serveStealReq_valid),
		.connArgumentNotifier_2_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_2_ctrl_serveStealReq_ready),
		.connArgumentNotifier_2_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_2_data_qOutTask_ready),
		.connArgumentNotifier_2_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_2_data_qOutTask_valid),
		.connArgumentNotifier_2_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_2_data_qOutTask_bits),
		.connArgumentNotifier_3_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_3_ctrl_serveStealReq_valid),
		.connArgumentNotifier_3_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_3_ctrl_serveStealReq_ready),
		.connArgumentNotifier_3_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_3_data_qOutTask_ready),
		.connArgumentNotifier_3_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_3_data_qOutTask_valid),
		.connArgumentNotifier_3_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_3_data_qOutTask_bits),
		.connArgumentNotifier_4_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_4_ctrl_serveStealReq_valid),
		.connArgumentNotifier_4_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_4_ctrl_serveStealReq_ready),
		.connArgumentNotifier_4_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_4_data_qOutTask_ready),
		.connArgumentNotifier_4_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_4_data_qOutTask_valid),
		.connArgumentNotifier_4_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_4_data_qOutTask_bits),
		.connArgumentNotifier_5_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_5_ctrl_serveStealReq_valid),
		.connArgumentNotifier_5_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_5_ctrl_serveStealReq_ready),
		.connArgumentNotifier_5_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_5_data_qOutTask_ready),
		.connArgumentNotifier_5_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_5_data_qOutTask_valid),
		.connArgumentNotifier_5_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_5_data_qOutTask_bits),
		.connArgumentNotifier_6_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_6_ctrl_serveStealReq_valid),
		.connArgumentNotifier_6_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_6_ctrl_serveStealReq_ready),
		.connArgumentNotifier_6_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_6_data_qOutTask_ready),
		.connArgumentNotifier_6_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_6_data_qOutTask_valid),
		.connArgumentNotifier_6_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_6_data_qOutTask_bits),
		.connArgumentNotifier_7_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_7_ctrl_serveStealReq_valid),
		.connArgumentNotifier_7_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_7_ctrl_serveStealReq_ready),
		.connArgumentNotifier_7_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_7_data_qOutTask_ready),
		.connArgumentNotifier_7_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_7_data_qOutTask_valid),
		.connArgumentNotifier_7_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_7_data_qOutTask_bits),
		.connArgumentNotifier_8_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_8_ctrl_serveStealReq_valid),
		.connArgumentNotifier_8_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_8_ctrl_serveStealReq_ready),
		.connArgumentNotifier_8_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_8_data_qOutTask_ready),
		.connArgumentNotifier_8_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_8_data_qOutTask_valid),
		.connArgumentNotifier_8_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_8_data_qOutTask_bits),
		.connArgumentNotifier_9_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_9_ctrl_serveStealReq_valid),
		.connArgumentNotifier_9_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_9_ctrl_serveStealReq_ready),
		.connArgumentNotifier_9_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_9_data_qOutTask_ready),
		.connArgumentNotifier_9_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_9_data_qOutTask_valid),
		.connArgumentNotifier_9_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_9_data_qOutTask_bits),
		.connArgumentNotifier_10_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_10_ctrl_serveStealReq_valid),
		.connArgumentNotifier_10_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_10_ctrl_serveStealReq_ready),
		.connArgumentNotifier_10_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_10_data_qOutTask_ready),
		.connArgumentNotifier_10_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_10_data_qOutTask_valid),
		.connArgumentNotifier_10_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_10_data_qOutTask_bits),
		.connArgumentNotifier_11_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_11_ctrl_serveStealReq_valid),
		.connArgumentNotifier_11_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_11_ctrl_serveStealReq_ready),
		.connArgumentNotifier_11_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_11_data_qOutTask_ready),
		.connArgumentNotifier_11_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_11_data_qOutTask_valid),
		.connArgumentNotifier_11_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_11_data_qOutTask_bits),
		.connArgumentNotifier_12_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_12_ctrl_serveStealReq_valid),
		.connArgumentNotifier_12_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_12_ctrl_serveStealReq_ready),
		.connArgumentNotifier_12_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_12_data_qOutTask_ready),
		.connArgumentNotifier_12_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_12_data_qOutTask_valid),
		.connArgumentNotifier_12_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_12_data_qOutTask_bits),
		.connArgumentNotifier_13_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_13_ctrl_serveStealReq_valid),
		.connArgumentNotifier_13_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_13_ctrl_serveStealReq_ready),
		.connArgumentNotifier_13_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_13_data_qOutTask_ready),
		.connArgumentNotifier_13_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_13_data_qOutTask_valid),
		.connArgumentNotifier_13_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_13_data_qOutTask_bits),
		.connArgumentNotifier_14_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_14_ctrl_serveStealReq_valid),
		.connArgumentNotifier_14_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_14_ctrl_serveStealReq_ready),
		.connArgumentNotifier_14_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_14_data_qOutTask_ready),
		.connArgumentNotifier_14_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_14_data_qOutTask_valid),
		.connArgumentNotifier_14_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_14_data_qOutTask_bits),
		.connArgumentNotifier_15_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_15_ctrl_serveStealReq_valid),
		.connArgumentNotifier_15_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_15_ctrl_serveStealReq_ready),
		.connArgumentNotifier_15_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_15_data_qOutTask_ready),
		.connArgumentNotifier_15_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_15_data_qOutTask_valid),
		.connArgumentNotifier_15_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_15_data_qOutTask_bits)
	);
	Allocator Allocator(
		.clock(clock),
		.reset(reset),
		.io_export_closureOut_0_TREADY(_peArray_0_closureIn_TREADY),
		.io_export_closureOut_0_TVALID(_Allocator_io_export_closureOut_0_TVALID),
		.io_export_closureOut_1_TREADY(_peArray_1_closureIn_TREADY),
		.io_export_closureOut_1_TVALID(_Allocator_io_export_closureOut_1_TVALID),
		.io_export_closureOut_2_TREADY(_peArray_2_closureIn_TREADY),
		.io_export_closureOut_2_TVALID(_Allocator_io_export_closureOut_2_TVALID),
		.io_export_closureOut_3_TREADY(_peArray_3_closureIn_TREADY),
		.io_export_closureOut_3_TVALID(_Allocator_io_export_closureOut_3_TVALID),
		.io_export_closureOut_4_TREADY(_peArray_4_closureIn_TREADY),
		.io_export_closureOut_4_TVALID(_Allocator_io_export_closureOut_4_TVALID),
		.io_export_closureOut_5_TREADY(_peArray_5_closureIn_TREADY),
		.io_export_closureOut_5_TVALID(_Allocator_io_export_closureOut_5_TVALID),
		.io_export_closureOut_6_TREADY(_peArray_6_closureIn_TREADY),
		.io_export_closureOut_6_TVALID(_Allocator_io_export_closureOut_6_TVALID),
		.io_export_closureOut_7_TREADY(_peArray_7_closureIn_TREADY),
		.io_export_closureOut_7_TVALID(_Allocator_io_export_closureOut_7_TVALID),
		.io_export_closureOut_8_TREADY(_peArray_8_closureIn_TREADY),
		.io_export_closureOut_8_TVALID(_Allocator_io_export_closureOut_8_TVALID),
		.io_export_closureOut_9_TREADY(_peArray_9_closureIn_TREADY),
		.io_export_closureOut_9_TVALID(_Allocator_io_export_closureOut_9_TVALID),
		.io_export_closureOut_10_TREADY(_peArray_10_closureIn_TREADY),
		.io_export_closureOut_10_TVALID(_Allocator_io_export_closureOut_10_TVALID),
		.io_export_closureOut_11_TREADY(_peArray_11_closureIn_TREADY),
		.io_export_closureOut_11_TVALID(_Allocator_io_export_closureOut_11_TVALID),
		.io_export_closureOut_12_TREADY(_peArray_12_closureIn_TREADY),
		.io_export_closureOut_12_TVALID(_Allocator_io_export_closureOut_12_TVALID),
		.io_export_closureOut_13_TREADY(_peArray_13_closureIn_TREADY),
		.io_export_closureOut_13_TVALID(_Allocator_io_export_closureOut_13_TVALID),
		.io_export_closureOut_14_TREADY(_peArray_14_closureIn_TREADY),
		.io_export_closureOut_14_TVALID(_Allocator_io_export_closureOut_14_TVALID),
		.io_export_closureOut_15_TREADY(_peArray_15_closureIn_TREADY),
		.io_export_closureOut_15_TVALID(_Allocator_io_export_closureOut_15_TVALID),
		.io_export_closureOut_16_TREADY(_peArray_16_closureIn_TREADY),
		.io_export_closureOut_16_TVALID(_Allocator_io_export_closureOut_16_TVALID),
		.io_export_closureOut_17_TREADY(_peArray_17_closureIn_TREADY),
		.io_export_closureOut_17_TVALID(_Allocator_io_export_closureOut_17_TVALID),
		.io_export_closureOut_18_TREADY(_peArray_18_closureIn_TREADY),
		.io_export_closureOut_18_TVALID(_Allocator_io_export_closureOut_18_TVALID),
		.io_export_closureOut_19_TREADY(_peArray_19_closureIn_TREADY),
		.io_export_closureOut_19_TVALID(_Allocator_io_export_closureOut_19_TVALID),
		.io_export_closureOut_20_TREADY(_peArray_20_closureIn_TREADY),
		.io_export_closureOut_20_TVALID(_Allocator_io_export_closureOut_20_TVALID),
		.io_export_closureOut_21_TREADY(_peArray_21_closureIn_TREADY),
		.io_export_closureOut_21_TVALID(_Allocator_io_export_closureOut_21_TVALID),
		.io_export_closureOut_22_TREADY(_peArray_22_closureIn_TREADY),
		.io_export_closureOut_22_TVALID(_Allocator_io_export_closureOut_22_TVALID),
		.io_export_closureOut_23_TREADY(_peArray_23_closureIn_TREADY),
		.io_export_closureOut_23_TVALID(_Allocator_io_export_closureOut_23_TVALID),
		.io_export_closureOut_24_TREADY(_peArray_24_closureIn_TREADY),
		.io_export_closureOut_24_TVALID(_Allocator_io_export_closureOut_24_TVALID),
		.io_export_closureOut_25_TREADY(_peArray_25_closureIn_TREADY),
		.io_export_closureOut_25_TVALID(_Allocator_io_export_closureOut_25_TVALID),
		.io_export_closureOut_26_TREADY(_peArray_26_closureIn_TREADY),
		.io_export_closureOut_26_TVALID(_Allocator_io_export_closureOut_26_TVALID),
		.io_export_closureOut_27_TREADY(_peArray_27_closureIn_TREADY),
		.io_export_closureOut_27_TVALID(_Allocator_io_export_closureOut_27_TVALID),
		.io_export_closureOut_28_TREADY(_peArray_28_closureIn_TREADY),
		.io_export_closureOut_28_TVALID(_Allocator_io_export_closureOut_28_TVALID),
		.io_export_closureOut_29_TREADY(_peArray_29_closureIn_TREADY),
		.io_export_closureOut_29_TVALID(_Allocator_io_export_closureOut_29_TVALID),
		.io_export_closureOut_30_TREADY(_peArray_30_closureIn_TREADY),
		.io_export_closureOut_30_TVALID(_Allocator_io_export_closureOut_30_TVALID),
		.io_export_closureOut_31_TREADY(_peArray_31_closureIn_TREADY),
		.io_export_closureOut_31_TVALID(_Allocator_io_export_closureOut_31_TVALID),
		.io_export_closureOut_32_TREADY(_peArray_32_closureIn_TREADY),
		.io_export_closureOut_32_TVALID(_Allocator_io_export_closureOut_32_TVALID),
		.io_export_closureOut_33_TREADY(_peArray_33_closureIn_TREADY),
		.io_export_closureOut_33_TVALID(_Allocator_io_export_closureOut_33_TVALID),
		.io_export_closureOut_34_TREADY(_peArray_34_closureIn_TREADY),
		.io_export_closureOut_34_TVALID(_Allocator_io_export_closureOut_34_TVALID),
		.io_export_closureOut_35_TREADY(_peArray_35_closureIn_TREADY),
		.io_export_closureOut_35_TVALID(_Allocator_io_export_closureOut_35_TVALID),
		.io_export_closureOut_36_TREADY(_peArray_36_closureIn_TREADY),
		.io_export_closureOut_36_TVALID(_Allocator_io_export_closureOut_36_TVALID),
		.io_export_closureOut_37_TREADY(_peArray_37_closureIn_TREADY),
		.io_export_closureOut_37_TVALID(_Allocator_io_export_closureOut_37_TVALID),
		.io_export_closureOut_38_TREADY(_peArray_38_closureIn_TREADY),
		.io_export_closureOut_38_TVALID(_Allocator_io_export_closureOut_38_TVALID),
		.io_export_closureOut_39_TREADY(_peArray_39_closureIn_TREADY),
		.io_export_closureOut_39_TVALID(_Allocator_io_export_closureOut_39_TVALID),
		.io_export_closureOut_40_TREADY(_peArray_40_closureIn_TREADY),
		.io_export_closureOut_40_TVALID(_Allocator_io_export_closureOut_40_TVALID),
		.io_export_closureOut_41_TREADY(_peArray_41_closureIn_TREADY),
		.io_export_closureOut_41_TVALID(_Allocator_io_export_closureOut_41_TVALID),
		.io_export_closureOut_42_TREADY(_peArray_42_closureIn_TREADY),
		.io_export_closureOut_42_TVALID(_Allocator_io_export_closureOut_42_TVALID),
		.io_export_closureOut_43_TREADY(_peArray_43_closureIn_TREADY),
		.io_export_closureOut_43_TVALID(_Allocator_io_export_closureOut_43_TVALID),
		.io_export_closureOut_44_TREADY(_peArray_44_closureIn_TREADY),
		.io_export_closureOut_44_TVALID(_Allocator_io_export_closureOut_44_TVALID),
		.io_export_closureOut_45_TREADY(_peArray_45_closureIn_TREADY),
		.io_export_closureOut_45_TVALID(_Allocator_io_export_closureOut_45_TVALID),
		.io_export_closureOut_46_TREADY(_peArray_46_closureIn_TREADY),
		.io_export_closureOut_46_TVALID(_Allocator_io_export_closureOut_46_TVALID),
		.io_export_closureOut_47_TREADY(_peArray_47_closureIn_TREADY),
		.io_export_closureOut_47_TVALID(_Allocator_io_export_closureOut_47_TVALID),
		.io_export_closureOut_48_TREADY(_peArray_48_closureIn_TREADY),
		.io_export_closureOut_48_TVALID(_Allocator_io_export_closureOut_48_TVALID),
		.io_export_closureOut_49_TREADY(_peArray_49_closureIn_TREADY),
		.io_export_closureOut_49_TVALID(_Allocator_io_export_closureOut_49_TVALID),
		.io_export_closureOut_50_TREADY(_peArray_50_closureIn_TREADY),
		.io_export_closureOut_50_TVALID(_Allocator_io_export_closureOut_50_TVALID),
		.io_export_closureOut_51_TREADY(_peArray_51_closureIn_TREADY),
		.io_export_closureOut_51_TVALID(_Allocator_io_export_closureOut_51_TVALID),
		.io_export_closureOut_52_TREADY(_peArray_52_closureIn_TREADY),
		.io_export_closureOut_52_TVALID(_Allocator_io_export_closureOut_52_TVALID),
		.io_export_closureOut_53_TREADY(_peArray_53_closureIn_TREADY),
		.io_export_closureOut_53_TVALID(_Allocator_io_export_closureOut_53_TVALID),
		.io_export_closureOut_54_TREADY(_peArray_54_closureIn_TREADY),
		.io_export_closureOut_54_TVALID(_Allocator_io_export_closureOut_54_TVALID),
		.io_export_closureOut_55_TREADY(_peArray_55_closureIn_TREADY),
		.io_export_closureOut_55_TVALID(_Allocator_io_export_closureOut_55_TVALID),
		.io_export_closureOut_56_TREADY(_peArray_56_closureIn_TREADY),
		.io_export_closureOut_56_TVALID(_Allocator_io_export_closureOut_56_TVALID),
		.io_export_closureOut_57_TREADY(_peArray_57_closureIn_TREADY),
		.io_export_closureOut_57_TVALID(_Allocator_io_export_closureOut_57_TVALID),
		.io_export_closureOut_58_TREADY(_peArray_58_closureIn_TREADY),
		.io_export_closureOut_58_TVALID(_Allocator_io_export_closureOut_58_TVALID),
		.io_export_closureOut_59_TREADY(_peArray_59_closureIn_TREADY),
		.io_export_closureOut_59_TVALID(_Allocator_io_export_closureOut_59_TVALID),
		.io_export_closureOut_60_TREADY(_peArray_60_closureIn_TREADY),
		.io_export_closureOut_60_TVALID(_Allocator_io_export_closureOut_60_TVALID),
		.io_export_closureOut_61_TREADY(_peArray_61_closureIn_TREADY),
		.io_export_closureOut_61_TVALID(_Allocator_io_export_closureOut_61_TVALID),
		.io_export_closureOut_62_TREADY(_peArray_62_closureIn_TREADY),
		.io_export_closureOut_62_TVALID(_Allocator_io_export_closureOut_62_TVALID),
		.io_export_closureOut_63_TREADY(_peArray_63_closureIn_TREADY),
		.io_export_closureOut_63_TVALID(_Allocator_io_export_closureOut_63_TVALID),
		.io_internal_vcas_axi_full_0_ar_ready(sync_closureAllocatorAXI_0_ARREADY),
		.io_internal_vcas_axi_full_0_ar_valid(sync_closureAllocatorAXI_0_ARVALID),
		.io_internal_vcas_axi_full_0_ar_bits_addr(sync_closureAllocatorAXI_0_ARADDR),
		.io_internal_vcas_axi_full_0_r_ready(sync_closureAllocatorAXI_0_RREADY),
		.io_internal_vcas_axi_full_0_r_valid(sync_closureAllocatorAXI_0_RVALID),
		.io_internal_vcas_axi_full_0_r_bits_data(sync_closureAllocatorAXI_0_RDATA),
		.io_internal_vcas_axi_full_1_ar_ready(sync_closureAllocatorAXI_1_ARREADY),
		.io_internal_vcas_axi_full_1_ar_valid(sync_closureAllocatorAXI_1_ARVALID),
		.io_internal_vcas_axi_full_1_ar_bits_addr(sync_closureAllocatorAXI_1_ARADDR),
		.io_internal_vcas_axi_full_1_r_ready(sync_closureAllocatorAXI_1_RREADY),
		.io_internal_vcas_axi_full_1_r_valid(sync_closureAllocatorAXI_1_RVALID),
		.io_internal_vcas_axi_full_1_r_bits_data(sync_closureAllocatorAXI_1_RDATA),
		.io_internal_vcas_axi_full_2_ar_ready(sync_closureAllocatorAXI_2_ARREADY),
		.io_internal_vcas_axi_full_2_ar_valid(sync_closureAllocatorAXI_2_ARVALID),
		.io_internal_vcas_axi_full_2_ar_bits_addr(sync_closureAllocatorAXI_2_ARADDR),
		.io_internal_vcas_axi_full_2_r_ready(sync_closureAllocatorAXI_2_RREADY),
		.io_internal_vcas_axi_full_2_r_valid(sync_closureAllocatorAXI_2_RVALID),
		.io_internal_vcas_axi_full_2_r_bits_data(sync_closureAllocatorAXI_2_RDATA),
		.io_internal_vcas_axi_full_3_ar_ready(sync_closureAllocatorAXI_3_ARREADY),
		.io_internal_vcas_axi_full_3_ar_valid(sync_closureAllocatorAXI_3_ARVALID),
		.io_internal_vcas_axi_full_3_ar_bits_addr(sync_closureAllocatorAXI_3_ARADDR),
		.io_internal_vcas_axi_full_3_r_ready(sync_closureAllocatorAXI_3_RREADY),
		.io_internal_vcas_axi_full_3_r_valid(sync_closureAllocatorAXI_3_RVALID),
		.io_internal_vcas_axi_full_3_r_bits_data(sync_closureAllocatorAXI_3_RDATA),
		.io_internal_axi_mgmt_vcas_0_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_0_ar_ready),
		.io_internal_axi_mgmt_vcas_0_ar_valid(_demux_m_axil_2_ar_valid),
		.io_internal_axi_mgmt_vcas_0_ar_bits_addr(_demux_m_axil_2_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_0_ar_bits_prot(_demux_m_axil_2_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_0_r_ready(_demux_m_axil_2_r_ready),
		.io_internal_axi_mgmt_vcas_0_r_valid(_Allocator_io_internal_axi_mgmt_vcas_0_r_valid),
		.io_internal_axi_mgmt_vcas_0_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_data),
		.io_internal_axi_mgmt_vcas_0_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_r_bits_resp),
		.io_internal_axi_mgmt_vcas_0_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_0_aw_ready),
		.io_internal_axi_mgmt_vcas_0_aw_valid(_demux_m_axil_2_aw_valid),
		.io_internal_axi_mgmt_vcas_0_aw_bits_addr(_demux_m_axil_2_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_0_aw_bits_prot(_demux_m_axil_2_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_0_w_ready(_Allocator_io_internal_axi_mgmt_vcas_0_w_ready),
		.io_internal_axi_mgmt_vcas_0_w_valid(_demux_m_axil_2_w_valid),
		.io_internal_axi_mgmt_vcas_0_w_bits_data(_demux_m_axil_2_w_bits_data),
		.io_internal_axi_mgmt_vcas_0_w_bits_strb(_demux_m_axil_2_w_bits_strb),
		.io_internal_axi_mgmt_vcas_0_b_ready(_demux_m_axil_2_b_ready),
		.io_internal_axi_mgmt_vcas_0_b_valid(_Allocator_io_internal_axi_mgmt_vcas_0_b_valid),
		.io_internal_axi_mgmt_vcas_0_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_0_b_bits_resp),
		.io_internal_axi_mgmt_vcas_1_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_1_ar_ready),
		.io_internal_axi_mgmt_vcas_1_ar_valid(_demux_m_axil_3_ar_valid),
		.io_internal_axi_mgmt_vcas_1_ar_bits_addr(_demux_m_axil_3_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_1_ar_bits_prot(_demux_m_axil_3_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_1_r_ready(_demux_m_axil_3_r_ready),
		.io_internal_axi_mgmt_vcas_1_r_valid(_Allocator_io_internal_axi_mgmt_vcas_1_r_valid),
		.io_internal_axi_mgmt_vcas_1_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_data),
		.io_internal_axi_mgmt_vcas_1_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_r_bits_resp),
		.io_internal_axi_mgmt_vcas_1_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_1_aw_ready),
		.io_internal_axi_mgmt_vcas_1_aw_valid(_demux_m_axil_3_aw_valid),
		.io_internal_axi_mgmt_vcas_1_aw_bits_addr(_demux_m_axil_3_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_1_aw_bits_prot(_demux_m_axil_3_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_1_w_ready(_Allocator_io_internal_axi_mgmt_vcas_1_w_ready),
		.io_internal_axi_mgmt_vcas_1_w_valid(_demux_m_axil_3_w_valid),
		.io_internal_axi_mgmt_vcas_1_w_bits_data(_demux_m_axil_3_w_bits_data),
		.io_internal_axi_mgmt_vcas_1_w_bits_strb(_demux_m_axil_3_w_bits_strb),
		.io_internal_axi_mgmt_vcas_1_b_ready(_demux_m_axil_3_b_ready),
		.io_internal_axi_mgmt_vcas_1_b_valid(_Allocator_io_internal_axi_mgmt_vcas_1_b_valid),
		.io_internal_axi_mgmt_vcas_1_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_1_b_bits_resp),
		.io_internal_axi_mgmt_vcas_2_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_2_ar_ready),
		.io_internal_axi_mgmt_vcas_2_ar_valid(_demux_m_axil_4_ar_valid),
		.io_internal_axi_mgmt_vcas_2_ar_bits_addr(_demux_m_axil_4_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_2_ar_bits_prot(_demux_m_axil_4_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_2_r_ready(_demux_m_axil_4_r_ready),
		.io_internal_axi_mgmt_vcas_2_r_valid(_Allocator_io_internal_axi_mgmt_vcas_2_r_valid),
		.io_internal_axi_mgmt_vcas_2_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_data),
		.io_internal_axi_mgmt_vcas_2_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_r_bits_resp),
		.io_internal_axi_mgmt_vcas_2_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_2_aw_ready),
		.io_internal_axi_mgmt_vcas_2_aw_valid(_demux_m_axil_4_aw_valid),
		.io_internal_axi_mgmt_vcas_2_aw_bits_addr(_demux_m_axil_4_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_2_aw_bits_prot(_demux_m_axil_4_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_2_w_ready(_Allocator_io_internal_axi_mgmt_vcas_2_w_ready),
		.io_internal_axi_mgmt_vcas_2_w_valid(_demux_m_axil_4_w_valid),
		.io_internal_axi_mgmt_vcas_2_w_bits_data(_demux_m_axil_4_w_bits_data),
		.io_internal_axi_mgmt_vcas_2_w_bits_strb(_demux_m_axil_4_w_bits_strb),
		.io_internal_axi_mgmt_vcas_2_b_ready(_demux_m_axil_4_b_ready),
		.io_internal_axi_mgmt_vcas_2_b_valid(_Allocator_io_internal_axi_mgmt_vcas_2_b_valid),
		.io_internal_axi_mgmt_vcas_2_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_2_b_bits_resp),
		.io_internal_axi_mgmt_vcas_3_ar_ready(_Allocator_io_internal_axi_mgmt_vcas_3_ar_ready),
		.io_internal_axi_mgmt_vcas_3_ar_valid(_demux_m_axil_5_ar_valid),
		.io_internal_axi_mgmt_vcas_3_ar_bits_addr(_demux_m_axil_5_ar_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_3_ar_bits_prot(_demux_m_axil_5_ar_bits_prot),
		.io_internal_axi_mgmt_vcas_3_r_ready(_demux_m_axil_5_r_ready),
		.io_internal_axi_mgmt_vcas_3_r_valid(_Allocator_io_internal_axi_mgmt_vcas_3_r_valid),
		.io_internal_axi_mgmt_vcas_3_r_bits_data(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_data),
		.io_internal_axi_mgmt_vcas_3_r_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_r_bits_resp),
		.io_internal_axi_mgmt_vcas_3_aw_ready(_Allocator_io_internal_axi_mgmt_vcas_3_aw_ready),
		.io_internal_axi_mgmt_vcas_3_aw_valid(_demux_m_axil_5_aw_valid),
		.io_internal_axi_mgmt_vcas_3_aw_bits_addr(_demux_m_axil_5_aw_bits_addr[5:0]),
		.io_internal_axi_mgmt_vcas_3_aw_bits_prot(_demux_m_axil_5_aw_bits_prot),
		.io_internal_axi_mgmt_vcas_3_w_ready(_Allocator_io_internal_axi_mgmt_vcas_3_w_ready),
		.io_internal_axi_mgmt_vcas_3_w_valid(_demux_m_axil_5_w_valid),
		.io_internal_axi_mgmt_vcas_3_w_bits_data(_demux_m_axil_5_w_bits_data),
		.io_internal_axi_mgmt_vcas_3_w_bits_strb(_demux_m_axil_5_w_bits_strb),
		.io_internal_axi_mgmt_vcas_3_b_ready(_demux_m_axil_5_b_ready),
		.io_internal_axi_mgmt_vcas_3_b_valid(_Allocator_io_internal_axi_mgmt_vcas_3_b_valid),
		.io_internal_axi_mgmt_vcas_3_b_bits_resp(_Allocator_io_internal_axi_mgmt_vcas_3_b_bits_resp)
	);
	ArgumentNotifier ArgumentNotifier(
		.clock(clock),
		.reset(reset),
		.io_export_argIn_0_TREADY(_ArgumentNotifier_io_export_argIn_0_TREADY),
		.io_export_argIn_0_TVALID(_peArray_0_argOut_TVALID),
		.io_export_argIn_0_TDATA(_peArray_0_argOut_TDATA[31:0]),
		.io_export_argIn_1_TREADY(_ArgumentNotifier_io_export_argIn_1_TREADY),
		.io_export_argIn_1_TVALID(_peArray_1_argOut_TVALID),
		.io_export_argIn_1_TDATA(_peArray_1_argOut_TDATA[31:0]),
		.io_export_argIn_2_TREADY(_ArgumentNotifier_io_export_argIn_2_TREADY),
		.io_export_argIn_2_TVALID(_peArray_2_argOut_TVALID),
		.io_export_argIn_2_TDATA(_peArray_2_argOut_TDATA[31:0]),
		.io_export_argIn_3_TREADY(_ArgumentNotifier_io_export_argIn_3_TREADY),
		.io_export_argIn_3_TVALID(_peArray_3_argOut_TVALID),
		.io_export_argIn_3_TDATA(_peArray_3_argOut_TDATA[31:0]),
		.io_export_argIn_4_TREADY(_ArgumentNotifier_io_export_argIn_4_TREADY),
		.io_export_argIn_4_TVALID(_peArray_4_argOut_TVALID),
		.io_export_argIn_4_TDATA(_peArray_4_argOut_TDATA[31:0]),
		.io_export_argIn_5_TREADY(_ArgumentNotifier_io_export_argIn_5_TREADY),
		.io_export_argIn_5_TVALID(_peArray_5_argOut_TVALID),
		.io_export_argIn_5_TDATA(_peArray_5_argOut_TDATA[31:0]),
		.io_export_argIn_6_TREADY(_ArgumentNotifier_io_export_argIn_6_TREADY),
		.io_export_argIn_6_TVALID(_peArray_6_argOut_TVALID),
		.io_export_argIn_6_TDATA(_peArray_6_argOut_TDATA[31:0]),
		.io_export_argIn_7_TREADY(_ArgumentNotifier_io_export_argIn_7_TREADY),
		.io_export_argIn_7_TVALID(_peArray_7_argOut_TVALID),
		.io_export_argIn_7_TDATA(_peArray_7_argOut_TDATA[31:0]),
		.io_export_argIn_8_TREADY(_ArgumentNotifier_io_export_argIn_8_TREADY),
		.io_export_argIn_8_TVALID(_peArray_8_argOut_TVALID),
		.io_export_argIn_8_TDATA(_peArray_8_argOut_TDATA[31:0]),
		.io_export_argIn_9_TREADY(_ArgumentNotifier_io_export_argIn_9_TREADY),
		.io_export_argIn_9_TVALID(_peArray_9_argOut_TVALID),
		.io_export_argIn_9_TDATA(_peArray_9_argOut_TDATA[31:0]),
		.io_export_argIn_10_TREADY(_ArgumentNotifier_io_export_argIn_10_TREADY),
		.io_export_argIn_10_TVALID(_peArray_10_argOut_TVALID),
		.io_export_argIn_10_TDATA(_peArray_10_argOut_TDATA[31:0]),
		.io_export_argIn_11_TREADY(_ArgumentNotifier_io_export_argIn_11_TREADY),
		.io_export_argIn_11_TVALID(_peArray_11_argOut_TVALID),
		.io_export_argIn_11_TDATA(_peArray_11_argOut_TDATA[31:0]),
		.io_export_argIn_12_TREADY(_ArgumentNotifier_io_export_argIn_12_TREADY),
		.io_export_argIn_12_TVALID(_peArray_12_argOut_TVALID),
		.io_export_argIn_12_TDATA(_peArray_12_argOut_TDATA[31:0]),
		.io_export_argIn_13_TREADY(_ArgumentNotifier_io_export_argIn_13_TREADY),
		.io_export_argIn_13_TVALID(_peArray_13_argOut_TVALID),
		.io_export_argIn_13_TDATA(_peArray_13_argOut_TDATA[31:0]),
		.io_export_argIn_14_TREADY(_ArgumentNotifier_io_export_argIn_14_TREADY),
		.io_export_argIn_14_TVALID(_peArray_14_argOut_TVALID),
		.io_export_argIn_14_TDATA(_peArray_14_argOut_TDATA[31:0]),
		.io_export_argIn_15_TREADY(_ArgumentNotifier_io_export_argIn_15_TREADY),
		.io_export_argIn_15_TVALID(_peArray_15_argOut_TVALID),
		.io_export_argIn_15_TDATA(_peArray_15_argOut_TDATA[31:0]),
		.io_export_argIn_16_TREADY(_ArgumentNotifier_io_export_argIn_16_TREADY),
		.io_export_argIn_16_TVALID(_peArray_16_argOut_TVALID),
		.io_export_argIn_16_TDATA(_peArray_16_argOut_TDATA[31:0]),
		.io_export_argIn_17_TREADY(_ArgumentNotifier_io_export_argIn_17_TREADY),
		.io_export_argIn_17_TVALID(_peArray_17_argOut_TVALID),
		.io_export_argIn_17_TDATA(_peArray_17_argOut_TDATA[31:0]),
		.io_export_argIn_18_TREADY(_ArgumentNotifier_io_export_argIn_18_TREADY),
		.io_export_argIn_18_TVALID(_peArray_18_argOut_TVALID),
		.io_export_argIn_18_TDATA(_peArray_18_argOut_TDATA[31:0]),
		.io_export_argIn_19_TREADY(_ArgumentNotifier_io_export_argIn_19_TREADY),
		.io_export_argIn_19_TVALID(_peArray_19_argOut_TVALID),
		.io_export_argIn_19_TDATA(_peArray_19_argOut_TDATA[31:0]),
		.io_export_argIn_20_TREADY(_ArgumentNotifier_io_export_argIn_20_TREADY),
		.io_export_argIn_20_TVALID(_peArray_20_argOut_TVALID),
		.io_export_argIn_20_TDATA(_peArray_20_argOut_TDATA[31:0]),
		.io_export_argIn_21_TREADY(_ArgumentNotifier_io_export_argIn_21_TREADY),
		.io_export_argIn_21_TVALID(_peArray_21_argOut_TVALID),
		.io_export_argIn_21_TDATA(_peArray_21_argOut_TDATA[31:0]),
		.io_export_argIn_22_TREADY(_ArgumentNotifier_io_export_argIn_22_TREADY),
		.io_export_argIn_22_TVALID(_peArray_22_argOut_TVALID),
		.io_export_argIn_22_TDATA(_peArray_22_argOut_TDATA[31:0]),
		.io_export_argIn_23_TREADY(_ArgumentNotifier_io_export_argIn_23_TREADY),
		.io_export_argIn_23_TVALID(_peArray_23_argOut_TVALID),
		.io_export_argIn_23_TDATA(_peArray_23_argOut_TDATA[31:0]),
		.io_export_argIn_24_TREADY(_ArgumentNotifier_io_export_argIn_24_TREADY),
		.io_export_argIn_24_TVALID(_peArray_24_argOut_TVALID),
		.io_export_argIn_24_TDATA(_peArray_24_argOut_TDATA[31:0]),
		.io_export_argIn_25_TREADY(_ArgumentNotifier_io_export_argIn_25_TREADY),
		.io_export_argIn_25_TVALID(_peArray_25_argOut_TVALID),
		.io_export_argIn_25_TDATA(_peArray_25_argOut_TDATA[31:0]),
		.io_export_argIn_26_TREADY(_ArgumentNotifier_io_export_argIn_26_TREADY),
		.io_export_argIn_26_TVALID(_peArray_26_argOut_TVALID),
		.io_export_argIn_26_TDATA(_peArray_26_argOut_TDATA[31:0]),
		.io_export_argIn_27_TREADY(_ArgumentNotifier_io_export_argIn_27_TREADY),
		.io_export_argIn_27_TVALID(_peArray_27_argOut_TVALID),
		.io_export_argIn_27_TDATA(_peArray_27_argOut_TDATA[31:0]),
		.io_export_argIn_28_TREADY(_ArgumentNotifier_io_export_argIn_28_TREADY),
		.io_export_argIn_28_TVALID(_peArray_28_argOut_TVALID),
		.io_export_argIn_28_TDATA(_peArray_28_argOut_TDATA[31:0]),
		.io_export_argIn_29_TREADY(_ArgumentNotifier_io_export_argIn_29_TREADY),
		.io_export_argIn_29_TVALID(_peArray_29_argOut_TVALID),
		.io_export_argIn_29_TDATA(_peArray_29_argOut_TDATA[31:0]),
		.io_export_argIn_30_TREADY(_ArgumentNotifier_io_export_argIn_30_TREADY),
		.io_export_argIn_30_TVALID(_peArray_30_argOut_TVALID),
		.io_export_argIn_30_TDATA(_peArray_30_argOut_TDATA[31:0]),
		.io_export_argIn_31_TREADY(_ArgumentNotifier_io_export_argIn_31_TREADY),
		.io_export_argIn_31_TVALID(_peArray_31_argOut_TVALID),
		.io_export_argIn_31_TDATA(_peArray_31_argOut_TDATA[31:0]),
		.io_export_argIn_32_TREADY(_ArgumentNotifier_io_export_argIn_32_TREADY),
		.io_export_argIn_32_TVALID(_peArray_32_argOut_TVALID),
		.io_export_argIn_32_TDATA(_peArray_32_argOut_TDATA[31:0]),
		.io_export_argIn_33_TREADY(_ArgumentNotifier_io_export_argIn_33_TREADY),
		.io_export_argIn_33_TVALID(_peArray_33_argOut_TVALID),
		.io_export_argIn_33_TDATA(_peArray_33_argOut_TDATA[31:0]),
		.io_export_argIn_34_TREADY(_ArgumentNotifier_io_export_argIn_34_TREADY),
		.io_export_argIn_34_TVALID(_peArray_34_argOut_TVALID),
		.io_export_argIn_34_TDATA(_peArray_34_argOut_TDATA[31:0]),
		.io_export_argIn_35_TREADY(_ArgumentNotifier_io_export_argIn_35_TREADY),
		.io_export_argIn_35_TVALID(_peArray_35_argOut_TVALID),
		.io_export_argIn_35_TDATA(_peArray_35_argOut_TDATA[31:0]),
		.io_export_argIn_36_TREADY(_ArgumentNotifier_io_export_argIn_36_TREADY),
		.io_export_argIn_36_TVALID(_peArray_36_argOut_TVALID),
		.io_export_argIn_36_TDATA(_peArray_36_argOut_TDATA[31:0]),
		.io_export_argIn_37_TREADY(_ArgumentNotifier_io_export_argIn_37_TREADY),
		.io_export_argIn_37_TVALID(_peArray_37_argOut_TVALID),
		.io_export_argIn_37_TDATA(_peArray_37_argOut_TDATA[31:0]),
		.io_export_argIn_38_TREADY(_ArgumentNotifier_io_export_argIn_38_TREADY),
		.io_export_argIn_38_TVALID(_peArray_38_argOut_TVALID),
		.io_export_argIn_38_TDATA(_peArray_38_argOut_TDATA[31:0]),
		.io_export_argIn_39_TREADY(_ArgumentNotifier_io_export_argIn_39_TREADY),
		.io_export_argIn_39_TVALID(_peArray_39_argOut_TVALID),
		.io_export_argIn_39_TDATA(_peArray_39_argOut_TDATA[31:0]),
		.io_export_argIn_40_TREADY(_ArgumentNotifier_io_export_argIn_40_TREADY),
		.io_export_argIn_40_TVALID(_peArray_40_argOut_TVALID),
		.io_export_argIn_40_TDATA(_peArray_40_argOut_TDATA[31:0]),
		.io_export_argIn_41_TREADY(_ArgumentNotifier_io_export_argIn_41_TREADY),
		.io_export_argIn_41_TVALID(_peArray_41_argOut_TVALID),
		.io_export_argIn_41_TDATA(_peArray_41_argOut_TDATA[31:0]),
		.io_export_argIn_42_TREADY(_ArgumentNotifier_io_export_argIn_42_TREADY),
		.io_export_argIn_42_TVALID(_peArray_42_argOut_TVALID),
		.io_export_argIn_42_TDATA(_peArray_42_argOut_TDATA[31:0]),
		.io_export_argIn_43_TREADY(_ArgumentNotifier_io_export_argIn_43_TREADY),
		.io_export_argIn_43_TVALID(_peArray_43_argOut_TVALID),
		.io_export_argIn_43_TDATA(_peArray_43_argOut_TDATA[31:0]),
		.io_export_argIn_44_TREADY(_ArgumentNotifier_io_export_argIn_44_TREADY),
		.io_export_argIn_44_TVALID(_peArray_44_argOut_TVALID),
		.io_export_argIn_44_TDATA(_peArray_44_argOut_TDATA[31:0]),
		.io_export_argIn_45_TREADY(_ArgumentNotifier_io_export_argIn_45_TREADY),
		.io_export_argIn_45_TVALID(_peArray_45_argOut_TVALID),
		.io_export_argIn_45_TDATA(_peArray_45_argOut_TDATA[31:0]),
		.io_export_argIn_46_TREADY(_ArgumentNotifier_io_export_argIn_46_TREADY),
		.io_export_argIn_46_TVALID(_peArray_46_argOut_TVALID),
		.io_export_argIn_46_TDATA(_peArray_46_argOut_TDATA[31:0]),
		.io_export_argIn_47_TREADY(_ArgumentNotifier_io_export_argIn_47_TREADY),
		.io_export_argIn_47_TVALID(_peArray_47_argOut_TVALID),
		.io_export_argIn_47_TDATA(_peArray_47_argOut_TDATA[31:0]),
		.io_export_argIn_48_TREADY(_ArgumentNotifier_io_export_argIn_48_TREADY),
		.io_export_argIn_48_TVALID(_peArray_48_argOut_TVALID),
		.io_export_argIn_48_TDATA(_peArray_48_argOut_TDATA[31:0]),
		.io_export_argIn_49_TREADY(_ArgumentNotifier_io_export_argIn_49_TREADY),
		.io_export_argIn_49_TVALID(_peArray_49_argOut_TVALID),
		.io_export_argIn_49_TDATA(_peArray_49_argOut_TDATA[31:0]),
		.io_export_argIn_50_TREADY(_ArgumentNotifier_io_export_argIn_50_TREADY),
		.io_export_argIn_50_TVALID(_peArray_50_argOut_TVALID),
		.io_export_argIn_50_TDATA(_peArray_50_argOut_TDATA[31:0]),
		.io_export_argIn_51_TREADY(_ArgumentNotifier_io_export_argIn_51_TREADY),
		.io_export_argIn_51_TVALID(_peArray_51_argOut_TVALID),
		.io_export_argIn_51_TDATA(_peArray_51_argOut_TDATA[31:0]),
		.io_export_argIn_52_TREADY(_ArgumentNotifier_io_export_argIn_52_TREADY),
		.io_export_argIn_52_TVALID(_peArray_52_argOut_TVALID),
		.io_export_argIn_52_TDATA(_peArray_52_argOut_TDATA[31:0]),
		.io_export_argIn_53_TREADY(_ArgumentNotifier_io_export_argIn_53_TREADY),
		.io_export_argIn_53_TVALID(_peArray_53_argOut_TVALID),
		.io_export_argIn_53_TDATA(_peArray_53_argOut_TDATA[31:0]),
		.io_export_argIn_54_TREADY(_ArgumentNotifier_io_export_argIn_54_TREADY),
		.io_export_argIn_54_TVALID(_peArray_54_argOut_TVALID),
		.io_export_argIn_54_TDATA(_peArray_54_argOut_TDATA[31:0]),
		.io_export_argIn_55_TREADY(_ArgumentNotifier_io_export_argIn_55_TREADY),
		.io_export_argIn_55_TVALID(_peArray_55_argOut_TVALID),
		.io_export_argIn_55_TDATA(_peArray_55_argOut_TDATA[31:0]),
		.io_export_argIn_56_TREADY(_ArgumentNotifier_io_export_argIn_56_TREADY),
		.io_export_argIn_56_TVALID(_peArray_56_argOut_TVALID),
		.io_export_argIn_56_TDATA(_peArray_56_argOut_TDATA[31:0]),
		.io_export_argIn_57_TREADY(_ArgumentNotifier_io_export_argIn_57_TREADY),
		.io_export_argIn_57_TVALID(_peArray_57_argOut_TVALID),
		.io_export_argIn_57_TDATA(_peArray_57_argOut_TDATA[31:0]),
		.io_export_argIn_58_TREADY(_ArgumentNotifier_io_export_argIn_58_TREADY),
		.io_export_argIn_58_TVALID(_peArray_58_argOut_TVALID),
		.io_export_argIn_58_TDATA(_peArray_58_argOut_TDATA[31:0]),
		.io_export_argIn_59_TREADY(_ArgumentNotifier_io_export_argIn_59_TREADY),
		.io_export_argIn_59_TVALID(_peArray_59_argOut_TVALID),
		.io_export_argIn_59_TDATA(_peArray_59_argOut_TDATA[31:0]),
		.io_export_argIn_60_TREADY(_ArgumentNotifier_io_export_argIn_60_TREADY),
		.io_export_argIn_60_TVALID(_peArray_60_argOut_TVALID),
		.io_export_argIn_60_TDATA(_peArray_60_argOut_TDATA[31:0]),
		.io_export_argIn_61_TREADY(_ArgumentNotifier_io_export_argIn_61_TREADY),
		.io_export_argIn_61_TVALID(_peArray_61_argOut_TVALID),
		.io_export_argIn_61_TDATA(_peArray_61_argOut_TDATA[31:0]),
		.io_export_argIn_62_TREADY(_ArgumentNotifier_io_export_argIn_62_TREADY),
		.io_export_argIn_62_TVALID(_peArray_62_argOut_TVALID),
		.io_export_argIn_62_TDATA(_peArray_62_argOut_TDATA[31:0]),
		.io_export_argIn_63_TREADY(_ArgumentNotifier_io_export_argIn_63_TREADY),
		.io_export_argIn_63_TVALID(_peArray_63_argOut_TVALID),
		.io_export_argIn_63_TDATA(_peArray_63_argOut_TDATA[31:0]),
		.io_export_argIn_64_TREADY(_ArgumentNotifier_io_export_argIn_64_TREADY),
		.io_export_argIn_64_TVALID(_peArray_0_1_argOut_TVALID),
		.io_export_argIn_64_TDATA(_peArray_0_1_argOut_TDATA[31:0]),
		.io_export_argIn_65_TREADY(_ArgumentNotifier_io_export_argIn_65_TREADY),
		.io_export_argIn_65_TVALID(_peArray_1_1_argOut_TVALID),
		.io_export_argIn_65_TDATA(_peArray_1_1_argOut_TDATA[31:0]),
		.io_export_argIn_66_TREADY(_ArgumentNotifier_io_export_argIn_66_TREADY),
		.io_export_argIn_66_TVALID(_peArray_2_1_argOut_TVALID),
		.io_export_argIn_66_TDATA(_peArray_2_1_argOut_TDATA[31:0]),
		.io_export_argIn_67_TREADY(_ArgumentNotifier_io_export_argIn_67_TREADY),
		.io_export_argIn_67_TVALID(_peArray_3_1_argOut_TVALID),
		.io_export_argIn_67_TDATA(_peArray_3_1_argOut_TDATA[31:0]),
		.io_export_argIn_68_TREADY(_ArgumentNotifier_io_export_argIn_68_TREADY),
		.io_export_argIn_68_TVALID(_peArray_4_1_argOut_TVALID),
		.io_export_argIn_68_TDATA(_peArray_4_1_argOut_TDATA[31:0]),
		.io_export_argIn_69_TREADY(_ArgumentNotifier_io_export_argIn_69_TREADY),
		.io_export_argIn_69_TVALID(_peArray_5_1_argOut_TVALID),
		.io_export_argIn_69_TDATA(_peArray_5_1_argOut_TDATA[31:0]),
		.io_export_argIn_70_TREADY(_ArgumentNotifier_io_export_argIn_70_TREADY),
		.io_export_argIn_70_TVALID(_peArray_6_1_argOut_TVALID),
		.io_export_argIn_70_TDATA(_peArray_6_1_argOut_TDATA[31:0]),
		.io_export_argIn_71_TREADY(_ArgumentNotifier_io_export_argIn_71_TREADY),
		.io_export_argIn_71_TVALID(_peArray_7_1_argOut_TVALID),
		.io_export_argIn_71_TDATA(_peArray_7_1_argOut_TDATA[31:0]),
		.io_export_argIn_72_TREADY(_ArgumentNotifier_io_export_argIn_72_TREADY),
		.io_export_argIn_72_TVALID(_peArray_8_1_argOut_TVALID),
		.io_export_argIn_72_TDATA(_peArray_8_1_argOut_TDATA[31:0]),
		.io_export_argIn_73_TREADY(_ArgumentNotifier_io_export_argIn_73_TREADY),
		.io_export_argIn_73_TVALID(_peArray_9_1_argOut_TVALID),
		.io_export_argIn_73_TDATA(_peArray_9_1_argOut_TDATA[31:0]),
		.io_export_argIn_74_TREADY(_ArgumentNotifier_io_export_argIn_74_TREADY),
		.io_export_argIn_74_TVALID(_peArray_10_1_argOut_TVALID),
		.io_export_argIn_74_TDATA(_peArray_10_1_argOut_TDATA[31:0]),
		.io_export_argIn_75_TREADY(_ArgumentNotifier_io_export_argIn_75_TREADY),
		.io_export_argIn_75_TVALID(_peArray_11_1_argOut_TVALID),
		.io_export_argIn_75_TDATA(_peArray_11_1_argOut_TDATA[31:0]),
		.io_export_argIn_76_TREADY(_ArgumentNotifier_io_export_argIn_76_TREADY),
		.io_export_argIn_76_TVALID(_peArray_12_1_argOut_TVALID),
		.io_export_argIn_76_TDATA(_peArray_12_1_argOut_TDATA[31:0]),
		.io_export_argIn_77_TREADY(_ArgumentNotifier_io_export_argIn_77_TREADY),
		.io_export_argIn_77_TVALID(_peArray_13_1_argOut_TVALID),
		.io_export_argIn_77_TDATA(_peArray_13_1_argOut_TDATA[31:0]),
		.io_export_argIn_78_TREADY(_ArgumentNotifier_io_export_argIn_78_TREADY),
		.io_export_argIn_78_TVALID(_peArray_14_1_argOut_TVALID),
		.io_export_argIn_78_TDATA(_peArray_14_1_argOut_TDATA[31:0]),
		.io_export_argIn_79_TREADY(_ArgumentNotifier_io_export_argIn_79_TREADY),
		.io_export_argIn_79_TVALID(_peArray_15_1_argOut_TVALID),
		.io_export_argIn_79_TDATA(_peArray_15_1_argOut_TDATA[31:0]),
		.connStealNtw_0_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_0_ctrl_serveStealReq_valid),
		.connStealNtw_0_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_0_ctrl_serveStealReq_ready),
		.connStealNtw_0_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_0_data_qOutTask_ready),
		.connStealNtw_0_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_0_data_qOutTask_valid),
		.connStealNtw_0_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_0_data_qOutTask_bits),
		.connStealNtw_1_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_1_ctrl_serveStealReq_valid),
		.connStealNtw_1_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_1_ctrl_serveStealReq_ready),
		.connStealNtw_1_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_1_data_qOutTask_ready),
		.connStealNtw_1_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_1_data_qOutTask_valid),
		.connStealNtw_1_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_1_data_qOutTask_bits),
		.connStealNtw_2_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_2_ctrl_serveStealReq_valid),
		.connStealNtw_2_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_2_ctrl_serveStealReq_ready),
		.connStealNtw_2_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_2_data_qOutTask_ready),
		.connStealNtw_2_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_2_data_qOutTask_valid),
		.connStealNtw_2_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_2_data_qOutTask_bits),
		.connStealNtw_3_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_3_ctrl_serveStealReq_valid),
		.connStealNtw_3_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_3_ctrl_serveStealReq_ready),
		.connStealNtw_3_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_3_data_qOutTask_ready),
		.connStealNtw_3_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_3_data_qOutTask_valid),
		.connStealNtw_3_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_3_data_qOutTask_bits),
		.connStealNtw_4_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_4_ctrl_serveStealReq_valid),
		.connStealNtw_4_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_4_ctrl_serveStealReq_ready),
		.connStealNtw_4_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_4_data_qOutTask_ready),
		.connStealNtw_4_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_4_data_qOutTask_valid),
		.connStealNtw_4_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_4_data_qOutTask_bits),
		.connStealNtw_5_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_5_ctrl_serveStealReq_valid),
		.connStealNtw_5_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_5_ctrl_serveStealReq_ready),
		.connStealNtw_5_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_5_data_qOutTask_ready),
		.connStealNtw_5_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_5_data_qOutTask_valid),
		.connStealNtw_5_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_5_data_qOutTask_bits),
		.connStealNtw_6_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_6_ctrl_serveStealReq_valid),
		.connStealNtw_6_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_6_ctrl_serveStealReq_ready),
		.connStealNtw_6_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_6_data_qOutTask_ready),
		.connStealNtw_6_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_6_data_qOutTask_valid),
		.connStealNtw_6_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_6_data_qOutTask_bits),
		.connStealNtw_7_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_7_ctrl_serveStealReq_valid),
		.connStealNtw_7_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_7_ctrl_serveStealReq_ready),
		.connStealNtw_7_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_7_data_qOutTask_ready),
		.connStealNtw_7_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_7_data_qOutTask_valid),
		.connStealNtw_7_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_7_data_qOutTask_bits),
		.connStealNtw_8_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_8_ctrl_serveStealReq_valid),
		.connStealNtw_8_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_8_ctrl_serveStealReq_ready),
		.connStealNtw_8_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_8_data_qOutTask_ready),
		.connStealNtw_8_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_8_data_qOutTask_valid),
		.connStealNtw_8_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_8_data_qOutTask_bits),
		.connStealNtw_9_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_9_ctrl_serveStealReq_valid),
		.connStealNtw_9_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_9_ctrl_serveStealReq_ready),
		.connStealNtw_9_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_9_data_qOutTask_ready),
		.connStealNtw_9_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_9_data_qOutTask_valid),
		.connStealNtw_9_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_9_data_qOutTask_bits),
		.connStealNtw_10_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_10_ctrl_serveStealReq_valid),
		.connStealNtw_10_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_10_ctrl_serveStealReq_ready),
		.connStealNtw_10_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_10_data_qOutTask_ready),
		.connStealNtw_10_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_10_data_qOutTask_valid),
		.connStealNtw_10_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_10_data_qOutTask_bits),
		.connStealNtw_11_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_11_ctrl_serveStealReq_valid),
		.connStealNtw_11_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_11_ctrl_serveStealReq_ready),
		.connStealNtw_11_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_11_data_qOutTask_ready),
		.connStealNtw_11_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_11_data_qOutTask_valid),
		.connStealNtw_11_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_11_data_qOutTask_bits),
		.connStealNtw_12_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_12_ctrl_serveStealReq_valid),
		.connStealNtw_12_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_12_ctrl_serveStealReq_ready),
		.connStealNtw_12_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_12_data_qOutTask_ready),
		.connStealNtw_12_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_12_data_qOutTask_valid),
		.connStealNtw_12_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_12_data_qOutTask_bits),
		.connStealNtw_13_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_13_ctrl_serveStealReq_valid),
		.connStealNtw_13_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_13_ctrl_serveStealReq_ready),
		.connStealNtw_13_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_13_data_qOutTask_ready),
		.connStealNtw_13_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_13_data_qOutTask_valid),
		.connStealNtw_13_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_13_data_qOutTask_bits),
		.connStealNtw_14_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_14_ctrl_serveStealReq_valid),
		.connStealNtw_14_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_14_ctrl_serveStealReq_ready),
		.connStealNtw_14_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_14_data_qOutTask_ready),
		.connStealNtw_14_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_14_data_qOutTask_valid),
		.connStealNtw_14_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_14_data_qOutTask_bits),
		.connStealNtw_15_ctrl_serveStealReq_valid(_ArgumentNotifier_connStealNtw_15_ctrl_serveStealReq_valid),
		.connStealNtw_15_ctrl_serveStealReq_ready(_Scheduler_1_connArgumentNotifier_15_ctrl_serveStealReq_ready),
		.connStealNtw_15_data_qOutTask_ready(_Scheduler_1_connArgumentNotifier_15_data_qOutTask_ready),
		.connStealNtw_15_data_qOutTask_valid(_ArgumentNotifier_connStealNtw_15_data_qOutTask_valid),
		.connStealNtw_15_data_qOutTask_bits(_ArgumentNotifier_connStealNtw_15_data_qOutTask_bits),
		.axi_full_argRoute_0_ar_ready(sync_argumentNotifierAXI_0_ARREADY),
		.axi_full_argRoute_0_ar_valid(sync_argumentNotifierAXI_0_ARVALID),
		.axi_full_argRoute_0_ar_bits_addr(sync_argumentNotifierAXI_0_ARADDR),
		.axi_full_argRoute_0_r_ready(sync_argumentNotifierAXI_0_RREADY),
		.axi_full_argRoute_0_r_valid(sync_argumentNotifierAXI_0_RVALID),
		.axi_full_argRoute_0_r_bits_data(sync_argumentNotifierAXI_0_RDATA),
		.axi_full_argRoute_0_aw_ready(sync_argumentNotifierAXI_0_AWREADY),
		.axi_full_argRoute_0_aw_valid(sync_argumentNotifierAXI_0_AWVALID),
		.axi_full_argRoute_0_aw_bits_addr(sync_argumentNotifierAXI_0_AWADDR),
		.axi_full_argRoute_0_w_ready(sync_argumentNotifierAXI_0_WREADY),
		.axi_full_argRoute_0_w_valid(sync_argumentNotifierAXI_0_WVALID),
		.axi_full_argRoute_0_w_bits_data(sync_argumentNotifierAXI_0_WDATA),
		.axi_full_argRoute_0_b_valid(sync_argumentNotifierAXI_0_BVALID),
		.axi_full_argRoute_1_ar_ready(sync_argumentNotifierAXI_1_ARREADY),
		.axi_full_argRoute_1_ar_valid(sync_argumentNotifierAXI_1_ARVALID),
		.axi_full_argRoute_1_ar_bits_addr(sync_argumentNotifierAXI_1_ARADDR),
		.axi_full_argRoute_1_r_ready(sync_argumentNotifierAXI_1_RREADY),
		.axi_full_argRoute_1_r_valid(sync_argumentNotifierAXI_1_RVALID),
		.axi_full_argRoute_1_r_bits_data(sync_argumentNotifierAXI_1_RDATA),
		.axi_full_argRoute_1_aw_ready(sync_argumentNotifierAXI_1_AWREADY),
		.axi_full_argRoute_1_aw_valid(sync_argumentNotifierAXI_1_AWVALID),
		.axi_full_argRoute_1_aw_bits_addr(sync_argumentNotifierAXI_1_AWADDR),
		.axi_full_argRoute_1_w_ready(sync_argumentNotifierAXI_1_WREADY),
		.axi_full_argRoute_1_w_valid(sync_argumentNotifierAXI_1_WVALID),
		.axi_full_argRoute_1_w_bits_data(sync_argumentNotifierAXI_1_WDATA),
		.axi_full_argRoute_1_b_valid(sync_argumentNotifierAXI_1_BVALID),
		.axi_full_argRoute_2_ar_ready(sync_argumentNotifierAXI_2_ARREADY),
		.axi_full_argRoute_2_ar_valid(sync_argumentNotifierAXI_2_ARVALID),
		.axi_full_argRoute_2_ar_bits_addr(sync_argumentNotifierAXI_2_ARADDR),
		.axi_full_argRoute_2_r_ready(sync_argumentNotifierAXI_2_RREADY),
		.axi_full_argRoute_2_r_valid(sync_argumentNotifierAXI_2_RVALID),
		.axi_full_argRoute_2_r_bits_data(sync_argumentNotifierAXI_2_RDATA),
		.axi_full_argRoute_2_aw_ready(sync_argumentNotifierAXI_2_AWREADY),
		.axi_full_argRoute_2_aw_valid(sync_argumentNotifierAXI_2_AWVALID),
		.axi_full_argRoute_2_aw_bits_addr(sync_argumentNotifierAXI_2_AWADDR),
		.axi_full_argRoute_2_w_ready(sync_argumentNotifierAXI_2_WREADY),
		.axi_full_argRoute_2_w_valid(sync_argumentNotifierAXI_2_WVALID),
		.axi_full_argRoute_2_w_bits_data(sync_argumentNotifierAXI_2_WDATA),
		.axi_full_argRoute_2_b_valid(sync_argumentNotifierAXI_2_BVALID),
		.axi_full_argRoute_3_ar_ready(sync_argumentNotifierAXI_3_ARREADY),
		.axi_full_argRoute_3_ar_valid(sync_argumentNotifierAXI_3_ARVALID),
		.axi_full_argRoute_3_ar_bits_addr(sync_argumentNotifierAXI_3_ARADDR),
		.axi_full_argRoute_3_r_ready(sync_argumentNotifierAXI_3_RREADY),
		.axi_full_argRoute_3_r_valid(sync_argumentNotifierAXI_3_RVALID),
		.axi_full_argRoute_3_r_bits_data(sync_argumentNotifierAXI_3_RDATA),
		.axi_full_argRoute_3_aw_ready(sync_argumentNotifierAXI_3_AWREADY),
		.axi_full_argRoute_3_aw_valid(sync_argumentNotifierAXI_3_AWVALID),
		.axi_full_argRoute_3_aw_bits_addr(sync_argumentNotifierAXI_3_AWADDR),
		.axi_full_argRoute_3_w_ready(sync_argumentNotifierAXI_3_WREADY),
		.axi_full_argRoute_3_w_valid(sync_argumentNotifierAXI_3_WVALID),
		.axi_full_argRoute_3_w_bits_data(sync_argumentNotifierAXI_3_WDATA),
		.axi_full_argRoute_3_b_valid(sync_argumentNotifierAXI_3_BVALID),
		.axi_full_argRoute_4_ar_ready(sync_argumentNotifierAXI_4_ARREADY),
		.axi_full_argRoute_4_ar_valid(sync_argumentNotifierAXI_4_ARVALID),
		.axi_full_argRoute_4_ar_bits_addr(sync_argumentNotifierAXI_4_ARADDR),
		.axi_full_argRoute_4_r_ready(sync_argumentNotifierAXI_4_RREADY),
		.axi_full_argRoute_4_r_valid(sync_argumentNotifierAXI_4_RVALID),
		.axi_full_argRoute_4_r_bits_data(sync_argumentNotifierAXI_4_RDATA),
		.axi_full_argRoute_4_aw_ready(sync_argumentNotifierAXI_4_AWREADY),
		.axi_full_argRoute_4_aw_valid(sync_argumentNotifierAXI_4_AWVALID),
		.axi_full_argRoute_4_aw_bits_addr(sync_argumentNotifierAXI_4_AWADDR),
		.axi_full_argRoute_4_w_ready(sync_argumentNotifierAXI_4_WREADY),
		.axi_full_argRoute_4_w_valid(sync_argumentNotifierAXI_4_WVALID),
		.axi_full_argRoute_4_w_bits_data(sync_argumentNotifierAXI_4_WDATA),
		.axi_full_argRoute_4_b_valid(sync_argumentNotifierAXI_4_BVALID),
		.axi_full_argRoute_5_ar_ready(sync_argumentNotifierAXI_5_ARREADY),
		.axi_full_argRoute_5_ar_valid(sync_argumentNotifierAXI_5_ARVALID),
		.axi_full_argRoute_5_ar_bits_addr(sync_argumentNotifierAXI_5_ARADDR),
		.axi_full_argRoute_5_r_ready(sync_argumentNotifierAXI_5_RREADY),
		.axi_full_argRoute_5_r_valid(sync_argumentNotifierAXI_5_RVALID),
		.axi_full_argRoute_5_r_bits_data(sync_argumentNotifierAXI_5_RDATA),
		.axi_full_argRoute_5_aw_ready(sync_argumentNotifierAXI_5_AWREADY),
		.axi_full_argRoute_5_aw_valid(sync_argumentNotifierAXI_5_AWVALID),
		.axi_full_argRoute_5_aw_bits_addr(sync_argumentNotifierAXI_5_AWADDR),
		.axi_full_argRoute_5_w_ready(sync_argumentNotifierAXI_5_WREADY),
		.axi_full_argRoute_5_w_valid(sync_argumentNotifierAXI_5_WVALID),
		.axi_full_argRoute_5_w_bits_data(sync_argumentNotifierAXI_5_WDATA),
		.axi_full_argRoute_5_b_valid(sync_argumentNotifierAXI_5_BVALID),
		.axi_full_argRoute_6_ar_ready(sync_argumentNotifierAXI_6_ARREADY),
		.axi_full_argRoute_6_ar_valid(sync_argumentNotifierAXI_6_ARVALID),
		.axi_full_argRoute_6_ar_bits_addr(sync_argumentNotifierAXI_6_ARADDR),
		.axi_full_argRoute_6_r_ready(sync_argumentNotifierAXI_6_RREADY),
		.axi_full_argRoute_6_r_valid(sync_argumentNotifierAXI_6_RVALID),
		.axi_full_argRoute_6_r_bits_data(sync_argumentNotifierAXI_6_RDATA),
		.axi_full_argRoute_6_aw_ready(sync_argumentNotifierAXI_6_AWREADY),
		.axi_full_argRoute_6_aw_valid(sync_argumentNotifierAXI_6_AWVALID),
		.axi_full_argRoute_6_aw_bits_addr(sync_argumentNotifierAXI_6_AWADDR),
		.axi_full_argRoute_6_w_ready(sync_argumentNotifierAXI_6_WREADY),
		.axi_full_argRoute_6_w_valid(sync_argumentNotifierAXI_6_WVALID),
		.axi_full_argRoute_6_w_bits_data(sync_argumentNotifierAXI_6_WDATA),
		.axi_full_argRoute_6_b_valid(sync_argumentNotifierAXI_6_BVALID),
		.axi_full_argRoute_7_ar_ready(sync_argumentNotifierAXI_7_ARREADY),
		.axi_full_argRoute_7_ar_valid(sync_argumentNotifierAXI_7_ARVALID),
		.axi_full_argRoute_7_ar_bits_addr(sync_argumentNotifierAXI_7_ARADDR),
		.axi_full_argRoute_7_r_ready(sync_argumentNotifierAXI_7_RREADY),
		.axi_full_argRoute_7_r_valid(sync_argumentNotifierAXI_7_RVALID),
		.axi_full_argRoute_7_r_bits_data(sync_argumentNotifierAXI_7_RDATA),
		.axi_full_argRoute_7_aw_ready(sync_argumentNotifierAXI_7_AWREADY),
		.axi_full_argRoute_7_aw_valid(sync_argumentNotifierAXI_7_AWVALID),
		.axi_full_argRoute_7_aw_bits_addr(sync_argumentNotifierAXI_7_AWADDR),
		.axi_full_argRoute_7_w_ready(sync_argumentNotifierAXI_7_WREADY),
		.axi_full_argRoute_7_w_valid(sync_argumentNotifierAXI_7_WVALID),
		.axi_full_argRoute_7_w_bits_data(sync_argumentNotifierAXI_7_WDATA),
		.axi_full_argRoute_7_b_valid(sync_argumentNotifierAXI_7_BVALID),
		.axi_full_argRoute_8_ar_ready(sync_argumentNotifierAXI_8_ARREADY),
		.axi_full_argRoute_8_ar_valid(sync_argumentNotifierAXI_8_ARVALID),
		.axi_full_argRoute_8_ar_bits_addr(sync_argumentNotifierAXI_8_ARADDR),
		.axi_full_argRoute_8_r_ready(sync_argumentNotifierAXI_8_RREADY),
		.axi_full_argRoute_8_r_valid(sync_argumentNotifierAXI_8_RVALID),
		.axi_full_argRoute_8_r_bits_data(sync_argumentNotifierAXI_8_RDATA),
		.axi_full_argRoute_8_aw_ready(sync_argumentNotifierAXI_8_AWREADY),
		.axi_full_argRoute_8_aw_valid(sync_argumentNotifierAXI_8_AWVALID),
		.axi_full_argRoute_8_aw_bits_addr(sync_argumentNotifierAXI_8_AWADDR),
		.axi_full_argRoute_8_w_ready(sync_argumentNotifierAXI_8_WREADY),
		.axi_full_argRoute_8_w_valid(sync_argumentNotifierAXI_8_WVALID),
		.axi_full_argRoute_8_w_bits_data(sync_argumentNotifierAXI_8_WDATA),
		.axi_full_argRoute_8_b_valid(sync_argumentNotifierAXI_8_BVALID),
		.axi_full_argRoute_9_ar_ready(sync_argumentNotifierAXI_9_ARREADY),
		.axi_full_argRoute_9_ar_valid(sync_argumentNotifierAXI_9_ARVALID),
		.axi_full_argRoute_9_ar_bits_addr(sync_argumentNotifierAXI_9_ARADDR),
		.axi_full_argRoute_9_r_ready(sync_argumentNotifierAXI_9_RREADY),
		.axi_full_argRoute_9_r_valid(sync_argumentNotifierAXI_9_RVALID),
		.axi_full_argRoute_9_r_bits_data(sync_argumentNotifierAXI_9_RDATA),
		.axi_full_argRoute_9_aw_ready(sync_argumentNotifierAXI_9_AWREADY),
		.axi_full_argRoute_9_aw_valid(sync_argumentNotifierAXI_9_AWVALID),
		.axi_full_argRoute_9_aw_bits_addr(sync_argumentNotifierAXI_9_AWADDR),
		.axi_full_argRoute_9_w_ready(sync_argumentNotifierAXI_9_WREADY),
		.axi_full_argRoute_9_w_valid(sync_argumentNotifierAXI_9_WVALID),
		.axi_full_argRoute_9_w_bits_data(sync_argumentNotifierAXI_9_WDATA),
		.axi_full_argRoute_9_b_valid(sync_argumentNotifierAXI_9_BVALID),
		.axi_full_argRoute_10_ar_ready(sync_argumentNotifierAXI_10_ARREADY),
		.axi_full_argRoute_10_ar_valid(sync_argumentNotifierAXI_10_ARVALID),
		.axi_full_argRoute_10_ar_bits_addr(sync_argumentNotifierAXI_10_ARADDR),
		.axi_full_argRoute_10_r_ready(sync_argumentNotifierAXI_10_RREADY),
		.axi_full_argRoute_10_r_valid(sync_argumentNotifierAXI_10_RVALID),
		.axi_full_argRoute_10_r_bits_data(sync_argumentNotifierAXI_10_RDATA),
		.axi_full_argRoute_10_aw_ready(sync_argumentNotifierAXI_10_AWREADY),
		.axi_full_argRoute_10_aw_valid(sync_argumentNotifierAXI_10_AWVALID),
		.axi_full_argRoute_10_aw_bits_addr(sync_argumentNotifierAXI_10_AWADDR),
		.axi_full_argRoute_10_w_ready(sync_argumentNotifierAXI_10_WREADY),
		.axi_full_argRoute_10_w_valid(sync_argumentNotifierAXI_10_WVALID),
		.axi_full_argRoute_10_w_bits_data(sync_argumentNotifierAXI_10_WDATA),
		.axi_full_argRoute_10_b_valid(sync_argumentNotifierAXI_10_BVALID),
		.axi_full_argRoute_11_ar_ready(sync_argumentNotifierAXI_11_ARREADY),
		.axi_full_argRoute_11_ar_valid(sync_argumentNotifierAXI_11_ARVALID),
		.axi_full_argRoute_11_ar_bits_addr(sync_argumentNotifierAXI_11_ARADDR),
		.axi_full_argRoute_11_r_ready(sync_argumentNotifierAXI_11_RREADY),
		.axi_full_argRoute_11_r_valid(sync_argumentNotifierAXI_11_RVALID),
		.axi_full_argRoute_11_r_bits_data(sync_argumentNotifierAXI_11_RDATA),
		.axi_full_argRoute_11_aw_ready(sync_argumentNotifierAXI_11_AWREADY),
		.axi_full_argRoute_11_aw_valid(sync_argumentNotifierAXI_11_AWVALID),
		.axi_full_argRoute_11_aw_bits_addr(sync_argumentNotifierAXI_11_AWADDR),
		.axi_full_argRoute_11_w_ready(sync_argumentNotifierAXI_11_WREADY),
		.axi_full_argRoute_11_w_valid(sync_argumentNotifierAXI_11_WVALID),
		.axi_full_argRoute_11_w_bits_data(sync_argumentNotifierAXI_11_WDATA),
		.axi_full_argRoute_11_b_valid(sync_argumentNotifierAXI_11_BVALID),
		.axi_full_argRoute_12_ar_ready(sync_argumentNotifierAXI_12_ARREADY),
		.axi_full_argRoute_12_ar_valid(sync_argumentNotifierAXI_12_ARVALID),
		.axi_full_argRoute_12_ar_bits_addr(sync_argumentNotifierAXI_12_ARADDR),
		.axi_full_argRoute_12_r_ready(sync_argumentNotifierAXI_12_RREADY),
		.axi_full_argRoute_12_r_valid(sync_argumentNotifierAXI_12_RVALID),
		.axi_full_argRoute_12_r_bits_data(sync_argumentNotifierAXI_12_RDATA),
		.axi_full_argRoute_12_aw_ready(sync_argumentNotifierAXI_12_AWREADY),
		.axi_full_argRoute_12_aw_valid(sync_argumentNotifierAXI_12_AWVALID),
		.axi_full_argRoute_12_aw_bits_addr(sync_argumentNotifierAXI_12_AWADDR),
		.axi_full_argRoute_12_w_ready(sync_argumentNotifierAXI_12_WREADY),
		.axi_full_argRoute_12_w_valid(sync_argumentNotifierAXI_12_WVALID),
		.axi_full_argRoute_12_w_bits_data(sync_argumentNotifierAXI_12_WDATA),
		.axi_full_argRoute_12_b_valid(sync_argumentNotifierAXI_12_BVALID),
		.axi_full_argRoute_13_ar_ready(sync_argumentNotifierAXI_13_ARREADY),
		.axi_full_argRoute_13_ar_valid(sync_argumentNotifierAXI_13_ARVALID),
		.axi_full_argRoute_13_ar_bits_addr(sync_argumentNotifierAXI_13_ARADDR),
		.axi_full_argRoute_13_r_ready(sync_argumentNotifierAXI_13_RREADY),
		.axi_full_argRoute_13_r_valid(sync_argumentNotifierAXI_13_RVALID),
		.axi_full_argRoute_13_r_bits_data(sync_argumentNotifierAXI_13_RDATA),
		.axi_full_argRoute_13_aw_ready(sync_argumentNotifierAXI_13_AWREADY),
		.axi_full_argRoute_13_aw_valid(sync_argumentNotifierAXI_13_AWVALID),
		.axi_full_argRoute_13_aw_bits_addr(sync_argumentNotifierAXI_13_AWADDR),
		.axi_full_argRoute_13_w_ready(sync_argumentNotifierAXI_13_WREADY),
		.axi_full_argRoute_13_w_valid(sync_argumentNotifierAXI_13_WVALID),
		.axi_full_argRoute_13_w_bits_data(sync_argumentNotifierAXI_13_WDATA),
		.axi_full_argRoute_13_b_valid(sync_argumentNotifierAXI_13_BVALID),
		.axi_full_argRoute_14_ar_ready(sync_argumentNotifierAXI_14_ARREADY),
		.axi_full_argRoute_14_ar_valid(sync_argumentNotifierAXI_14_ARVALID),
		.axi_full_argRoute_14_ar_bits_addr(sync_argumentNotifierAXI_14_ARADDR),
		.axi_full_argRoute_14_r_ready(sync_argumentNotifierAXI_14_RREADY),
		.axi_full_argRoute_14_r_valid(sync_argumentNotifierAXI_14_RVALID),
		.axi_full_argRoute_14_r_bits_data(sync_argumentNotifierAXI_14_RDATA),
		.axi_full_argRoute_14_aw_ready(sync_argumentNotifierAXI_14_AWREADY),
		.axi_full_argRoute_14_aw_valid(sync_argumentNotifierAXI_14_AWVALID),
		.axi_full_argRoute_14_aw_bits_addr(sync_argumentNotifierAXI_14_AWADDR),
		.axi_full_argRoute_14_w_ready(sync_argumentNotifierAXI_14_WREADY),
		.axi_full_argRoute_14_w_valid(sync_argumentNotifierAXI_14_WVALID),
		.axi_full_argRoute_14_w_bits_data(sync_argumentNotifierAXI_14_WDATA),
		.axi_full_argRoute_14_b_valid(sync_argumentNotifierAXI_14_BVALID),
		.axi_full_argRoute_15_ar_ready(sync_argumentNotifierAXI_15_ARREADY),
		.axi_full_argRoute_15_ar_valid(sync_argumentNotifierAXI_15_ARVALID),
		.axi_full_argRoute_15_ar_bits_addr(sync_argumentNotifierAXI_15_ARADDR),
		.axi_full_argRoute_15_r_ready(sync_argumentNotifierAXI_15_RREADY),
		.axi_full_argRoute_15_r_valid(sync_argumentNotifierAXI_15_RVALID),
		.axi_full_argRoute_15_r_bits_data(sync_argumentNotifierAXI_15_RDATA),
		.axi_full_argRoute_15_aw_ready(sync_argumentNotifierAXI_15_AWREADY),
		.axi_full_argRoute_15_aw_valid(sync_argumentNotifierAXI_15_AWVALID),
		.axi_full_argRoute_15_aw_bits_addr(sync_argumentNotifierAXI_15_AWADDR),
		.axi_full_argRoute_15_w_ready(sync_argumentNotifierAXI_15_WREADY),
		.axi_full_argRoute_15_w_valid(sync_argumentNotifierAXI_15_WVALID),
		.axi_full_argRoute_15_w_bits_data(sync_argumentNotifierAXI_15_WDATA),
		.axi_full_argRoute_15_b_valid(sync_argumentNotifierAXI_15_BVALID),
		.axi_full_argRoute_16_ar_ready(sync_argumentNotifierAXI_16_ARREADY),
		.axi_full_argRoute_16_ar_valid(sync_argumentNotifierAXI_16_ARVALID),
		.axi_full_argRoute_16_ar_bits_addr(sync_argumentNotifierAXI_16_ARADDR),
		.axi_full_argRoute_16_r_ready(sync_argumentNotifierAXI_16_RREADY),
		.axi_full_argRoute_16_r_valid(sync_argumentNotifierAXI_16_RVALID),
		.axi_full_argRoute_16_r_bits_data(sync_argumentNotifierAXI_16_RDATA),
		.axi_full_argRoute_17_ar_ready(sync_argumentNotifierAXI_17_ARREADY),
		.axi_full_argRoute_17_ar_valid(sync_argumentNotifierAXI_17_ARVALID),
		.axi_full_argRoute_17_ar_bits_addr(sync_argumentNotifierAXI_17_ARADDR),
		.axi_full_argRoute_17_r_ready(sync_argumentNotifierAXI_17_RREADY),
		.axi_full_argRoute_17_r_valid(sync_argumentNotifierAXI_17_RVALID),
		.axi_full_argRoute_17_r_bits_data(sync_argumentNotifierAXI_17_RDATA),
		.axi_full_argRoute_18_ar_ready(sync_argumentNotifierAXI_18_ARREADY),
		.axi_full_argRoute_18_ar_valid(sync_argumentNotifierAXI_18_ARVALID),
		.axi_full_argRoute_18_ar_bits_addr(sync_argumentNotifierAXI_18_ARADDR),
		.axi_full_argRoute_18_r_ready(sync_argumentNotifierAXI_18_RREADY),
		.axi_full_argRoute_18_r_valid(sync_argumentNotifierAXI_18_RVALID),
		.axi_full_argRoute_18_r_bits_data(sync_argumentNotifierAXI_18_RDATA),
		.axi_full_argRoute_19_ar_ready(sync_argumentNotifierAXI_19_ARREADY),
		.axi_full_argRoute_19_ar_valid(sync_argumentNotifierAXI_19_ARVALID),
		.axi_full_argRoute_19_ar_bits_addr(sync_argumentNotifierAXI_19_ARADDR),
		.axi_full_argRoute_19_r_ready(sync_argumentNotifierAXI_19_RREADY),
		.axi_full_argRoute_19_r_valid(sync_argumentNotifierAXI_19_RVALID),
		.axi_full_argRoute_19_r_bits_data(sync_argumentNotifierAXI_19_RDATA),
		.axi_full_argRoute_20_ar_ready(sync_argumentNotifierAXI_20_ARREADY),
		.axi_full_argRoute_20_ar_valid(sync_argumentNotifierAXI_20_ARVALID),
		.axi_full_argRoute_20_ar_bits_addr(sync_argumentNotifierAXI_20_ARADDR),
		.axi_full_argRoute_20_r_ready(sync_argumentNotifierAXI_20_RREADY),
		.axi_full_argRoute_20_r_valid(sync_argumentNotifierAXI_20_RVALID),
		.axi_full_argRoute_20_r_bits_data(sync_argumentNotifierAXI_20_RDATA),
		.axi_full_argRoute_21_ar_ready(sync_argumentNotifierAXI_21_ARREADY),
		.axi_full_argRoute_21_ar_valid(sync_argumentNotifierAXI_21_ARVALID),
		.axi_full_argRoute_21_ar_bits_addr(sync_argumentNotifierAXI_21_ARADDR),
		.axi_full_argRoute_21_r_ready(sync_argumentNotifierAXI_21_RREADY),
		.axi_full_argRoute_21_r_valid(sync_argumentNotifierAXI_21_RVALID),
		.axi_full_argRoute_21_r_bits_data(sync_argumentNotifierAXI_21_RDATA),
		.axi_full_argRoute_22_ar_ready(sync_argumentNotifierAXI_22_ARREADY),
		.axi_full_argRoute_22_ar_valid(sync_argumentNotifierAXI_22_ARVALID),
		.axi_full_argRoute_22_ar_bits_addr(sync_argumentNotifierAXI_22_ARADDR),
		.axi_full_argRoute_22_r_ready(sync_argumentNotifierAXI_22_RREADY),
		.axi_full_argRoute_22_r_valid(sync_argumentNotifierAXI_22_RVALID),
		.axi_full_argRoute_22_r_bits_data(sync_argumentNotifierAXI_22_RDATA),
		.axi_full_argRoute_23_ar_ready(sync_argumentNotifierAXI_23_ARREADY),
		.axi_full_argRoute_23_ar_valid(sync_argumentNotifierAXI_23_ARVALID),
		.axi_full_argRoute_23_ar_bits_addr(sync_argumentNotifierAXI_23_ARADDR),
		.axi_full_argRoute_23_r_ready(sync_argumentNotifierAXI_23_RREADY),
		.axi_full_argRoute_23_r_valid(sync_argumentNotifierAXI_23_RVALID),
		.axi_full_argRoute_23_r_bits_data(sync_argumentNotifierAXI_23_RDATA),
		.axi_full_argRoute_24_ar_ready(sync_argumentNotifierAXI_24_ARREADY),
		.axi_full_argRoute_24_ar_valid(sync_argumentNotifierAXI_24_ARVALID),
		.axi_full_argRoute_24_ar_bits_addr(sync_argumentNotifierAXI_24_ARADDR),
		.axi_full_argRoute_24_r_ready(sync_argumentNotifierAXI_24_RREADY),
		.axi_full_argRoute_24_r_valid(sync_argumentNotifierAXI_24_RVALID),
		.axi_full_argRoute_24_r_bits_data(sync_argumentNotifierAXI_24_RDATA),
		.axi_full_argRoute_25_ar_ready(sync_argumentNotifierAXI_25_ARREADY),
		.axi_full_argRoute_25_ar_valid(sync_argumentNotifierAXI_25_ARVALID),
		.axi_full_argRoute_25_ar_bits_addr(sync_argumentNotifierAXI_25_ARADDR),
		.axi_full_argRoute_25_r_ready(sync_argumentNotifierAXI_25_RREADY),
		.axi_full_argRoute_25_r_valid(sync_argumentNotifierAXI_25_RVALID),
		.axi_full_argRoute_25_r_bits_data(sync_argumentNotifierAXI_25_RDATA),
		.axi_full_argRoute_26_ar_ready(sync_argumentNotifierAXI_26_ARREADY),
		.axi_full_argRoute_26_ar_valid(sync_argumentNotifierAXI_26_ARVALID),
		.axi_full_argRoute_26_ar_bits_addr(sync_argumentNotifierAXI_26_ARADDR),
		.axi_full_argRoute_26_r_ready(sync_argumentNotifierAXI_26_RREADY),
		.axi_full_argRoute_26_r_valid(sync_argumentNotifierAXI_26_RVALID),
		.axi_full_argRoute_26_r_bits_data(sync_argumentNotifierAXI_26_RDATA),
		.axi_full_argRoute_27_ar_ready(sync_argumentNotifierAXI_27_ARREADY),
		.axi_full_argRoute_27_ar_valid(sync_argumentNotifierAXI_27_ARVALID),
		.axi_full_argRoute_27_ar_bits_addr(sync_argumentNotifierAXI_27_ARADDR),
		.axi_full_argRoute_27_r_ready(sync_argumentNotifierAXI_27_RREADY),
		.axi_full_argRoute_27_r_valid(sync_argumentNotifierAXI_27_RVALID),
		.axi_full_argRoute_27_r_bits_data(sync_argumentNotifierAXI_27_RDATA),
		.axi_full_argRoute_28_ar_ready(sync_argumentNotifierAXI_28_ARREADY),
		.axi_full_argRoute_28_ar_valid(sync_argumentNotifierAXI_28_ARVALID),
		.axi_full_argRoute_28_ar_bits_addr(sync_argumentNotifierAXI_28_ARADDR),
		.axi_full_argRoute_28_r_ready(sync_argumentNotifierAXI_28_RREADY),
		.axi_full_argRoute_28_r_valid(sync_argumentNotifierAXI_28_RVALID),
		.axi_full_argRoute_28_r_bits_data(sync_argumentNotifierAXI_28_RDATA),
		.axi_full_argRoute_29_ar_ready(sync_argumentNotifierAXI_29_ARREADY),
		.axi_full_argRoute_29_ar_valid(sync_argumentNotifierAXI_29_ARVALID),
		.axi_full_argRoute_29_ar_bits_addr(sync_argumentNotifierAXI_29_ARADDR),
		.axi_full_argRoute_29_r_ready(sync_argumentNotifierAXI_29_RREADY),
		.axi_full_argRoute_29_r_valid(sync_argumentNotifierAXI_29_RVALID),
		.axi_full_argRoute_29_r_bits_data(sync_argumentNotifierAXI_29_RDATA),
		.axi_full_argRoute_30_ar_ready(sync_argumentNotifierAXI_30_ARREADY),
		.axi_full_argRoute_30_ar_valid(sync_argumentNotifierAXI_30_ARVALID),
		.axi_full_argRoute_30_ar_bits_addr(sync_argumentNotifierAXI_30_ARADDR),
		.axi_full_argRoute_30_r_ready(sync_argumentNotifierAXI_30_RREADY),
		.axi_full_argRoute_30_r_valid(sync_argumentNotifierAXI_30_RVALID),
		.axi_full_argRoute_30_r_bits_data(sync_argumentNotifierAXI_30_RDATA),
		.axi_full_argRoute_31_ar_ready(sync_argumentNotifierAXI_31_ARREADY),
		.axi_full_argRoute_31_ar_valid(sync_argumentNotifierAXI_31_ARVALID),
		.axi_full_argRoute_31_ar_bits_addr(sync_argumentNotifierAXI_31_ARADDR),
		.axi_full_argRoute_31_r_ready(sync_argumentNotifierAXI_31_RREADY),
		.axi_full_argRoute_31_r_valid(sync_argumentNotifierAXI_31_RVALID),
		.axi_full_argRoute_31_r_bits_data(sync_argumentNotifierAXI_31_RDATA)
	);
	assign qsort_schedulerAXI_0_ARID = 1'h0;
	assign qsort_schedulerAXI_0_AWID = 1'h0;
	assign qsort_schedulerAXI_0_WSTRB = 32'hffffffff;
	assign qsort_schedulerAXI_0_BREADY = 1'h1;
	assign sync_schedulerAXI_0_ARID = 1'h0;
	assign sync_schedulerAXI_0_AWID = 1'h0;
	assign sync_schedulerAXI_0_WSTRB = 16'hffff;
	assign sync_schedulerAXI_0_BREADY = 1'h1;
	assign sync_closureAllocatorAXI_0_ARID = 5'h00;
	assign sync_closureAllocatorAXI_0_ARLEN = 8'h0f;
	assign sync_closureAllocatorAXI_0_ARSIZE = 3'h3;
	assign sync_closureAllocatorAXI_0_ARBURST = 2'h1;
	assign sync_closureAllocatorAXI_0_ARLOCK = 1'h0;
	assign sync_closureAllocatorAXI_0_ARCACHE = 4'h0;
	assign sync_closureAllocatorAXI_0_ARPROT = 3'h0;
	assign sync_closureAllocatorAXI_0_ARQOS = 4'h0;
	assign sync_closureAllocatorAXI_0_ARREGION = 4'h0;
	assign sync_closureAllocatorAXI_0_AWVALID = 1'h0;
	assign sync_closureAllocatorAXI_0_AWID = 5'h00;
	assign sync_closureAllocatorAXI_0_AWADDR = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_0_AWLEN = 8'h00;
	assign sync_closureAllocatorAXI_0_AWSIZE = 3'h0;
	assign sync_closureAllocatorAXI_0_AWBURST = 2'h0;
	assign sync_closureAllocatorAXI_0_AWLOCK = 1'h0;
	assign sync_closureAllocatorAXI_0_AWCACHE = 4'h0;
	assign sync_closureAllocatorAXI_0_AWPROT = 3'h0;
	assign sync_closureAllocatorAXI_0_AWQOS = 4'h0;
	assign sync_closureAllocatorAXI_0_AWREGION = 4'h0;
	assign sync_closureAllocatorAXI_0_WVALID = 1'h0;
	assign sync_closureAllocatorAXI_0_WDATA = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_0_WSTRB = 8'h00;
	assign sync_closureAllocatorAXI_0_WLAST = 1'h0;
	assign sync_closureAllocatorAXI_0_BREADY = 1'h0;
	assign sync_closureAllocatorAXI_1_ARID = 5'h00;
	assign sync_closureAllocatorAXI_1_ARLEN = 8'h0f;
	assign sync_closureAllocatorAXI_1_ARSIZE = 3'h3;
	assign sync_closureAllocatorAXI_1_ARBURST = 2'h1;
	assign sync_closureAllocatorAXI_1_ARLOCK = 1'h0;
	assign sync_closureAllocatorAXI_1_ARCACHE = 4'h0;
	assign sync_closureAllocatorAXI_1_ARPROT = 3'h0;
	assign sync_closureAllocatorAXI_1_ARQOS = 4'h0;
	assign sync_closureAllocatorAXI_1_ARREGION = 4'h0;
	assign sync_closureAllocatorAXI_1_AWVALID = 1'h0;
	assign sync_closureAllocatorAXI_1_AWID = 5'h00;
	assign sync_closureAllocatorAXI_1_AWADDR = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_1_AWLEN = 8'h00;
	assign sync_closureAllocatorAXI_1_AWSIZE = 3'h0;
	assign sync_closureAllocatorAXI_1_AWBURST = 2'h0;
	assign sync_closureAllocatorAXI_1_AWLOCK = 1'h0;
	assign sync_closureAllocatorAXI_1_AWCACHE = 4'h0;
	assign sync_closureAllocatorAXI_1_AWPROT = 3'h0;
	assign sync_closureAllocatorAXI_1_AWQOS = 4'h0;
	assign sync_closureAllocatorAXI_1_AWREGION = 4'h0;
	assign sync_closureAllocatorAXI_1_WVALID = 1'h0;
	assign sync_closureAllocatorAXI_1_WDATA = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_1_WSTRB = 8'h00;
	assign sync_closureAllocatorAXI_1_WLAST = 1'h0;
	assign sync_closureAllocatorAXI_1_BREADY = 1'h0;
	assign sync_closureAllocatorAXI_2_ARID = 5'h00;
	assign sync_closureAllocatorAXI_2_ARLEN = 8'h0f;
	assign sync_closureAllocatorAXI_2_ARSIZE = 3'h3;
	assign sync_closureAllocatorAXI_2_ARBURST = 2'h1;
	assign sync_closureAllocatorAXI_2_ARLOCK = 1'h0;
	assign sync_closureAllocatorAXI_2_ARCACHE = 4'h0;
	assign sync_closureAllocatorAXI_2_ARPROT = 3'h0;
	assign sync_closureAllocatorAXI_2_ARQOS = 4'h0;
	assign sync_closureAllocatorAXI_2_ARREGION = 4'h0;
	assign sync_closureAllocatorAXI_2_AWVALID = 1'h0;
	assign sync_closureAllocatorAXI_2_AWID = 5'h00;
	assign sync_closureAllocatorAXI_2_AWADDR = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_2_AWLEN = 8'h00;
	assign sync_closureAllocatorAXI_2_AWSIZE = 3'h0;
	assign sync_closureAllocatorAXI_2_AWBURST = 2'h0;
	assign sync_closureAllocatorAXI_2_AWLOCK = 1'h0;
	assign sync_closureAllocatorAXI_2_AWCACHE = 4'h0;
	assign sync_closureAllocatorAXI_2_AWPROT = 3'h0;
	assign sync_closureAllocatorAXI_2_AWQOS = 4'h0;
	assign sync_closureAllocatorAXI_2_AWREGION = 4'h0;
	assign sync_closureAllocatorAXI_2_WVALID = 1'h0;
	assign sync_closureAllocatorAXI_2_WDATA = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_2_WSTRB = 8'h00;
	assign sync_closureAllocatorAXI_2_WLAST = 1'h0;
	assign sync_closureAllocatorAXI_2_BREADY = 1'h0;
	assign sync_closureAllocatorAXI_3_ARID = 5'h00;
	assign sync_closureAllocatorAXI_3_ARLEN = 8'h0f;
	assign sync_closureAllocatorAXI_3_ARSIZE = 3'h3;
	assign sync_closureAllocatorAXI_3_ARBURST = 2'h1;
	assign sync_closureAllocatorAXI_3_ARLOCK = 1'h0;
	assign sync_closureAllocatorAXI_3_ARCACHE = 4'h0;
	assign sync_closureAllocatorAXI_3_ARPROT = 3'h0;
	assign sync_closureAllocatorAXI_3_ARQOS = 4'h0;
	assign sync_closureAllocatorAXI_3_ARREGION = 4'h0;
	assign sync_closureAllocatorAXI_3_AWVALID = 1'h0;
	assign sync_closureAllocatorAXI_3_AWID = 5'h00;
	assign sync_closureAllocatorAXI_3_AWADDR = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_3_AWLEN = 8'h00;
	assign sync_closureAllocatorAXI_3_AWSIZE = 3'h0;
	assign sync_closureAllocatorAXI_3_AWBURST = 2'h0;
	assign sync_closureAllocatorAXI_3_AWLOCK = 1'h0;
	assign sync_closureAllocatorAXI_3_AWCACHE = 4'h0;
	assign sync_closureAllocatorAXI_3_AWPROT = 3'h0;
	assign sync_closureAllocatorAXI_3_AWQOS = 4'h0;
	assign sync_closureAllocatorAXI_3_AWREGION = 4'h0;
	assign sync_closureAllocatorAXI_3_WVALID = 1'h0;
	assign sync_closureAllocatorAXI_3_WDATA = 64'h0000000000000000;
	assign sync_closureAllocatorAXI_3_WSTRB = 8'h00;
	assign sync_closureAllocatorAXI_3_WLAST = 1'h0;
	assign sync_closureAllocatorAXI_3_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_0_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_0_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_0_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_0_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_0_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_0_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_0_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_0_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_0_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_0_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_0_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_0_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_0_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_0_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_0_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_0_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_0_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_0_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_0_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_1_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_1_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_1_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_1_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_1_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_1_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_1_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_1_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_1_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_1_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_1_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_1_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_1_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_1_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_1_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_1_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_1_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_1_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_1_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_2_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_2_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_2_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_2_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_2_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_2_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_2_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_2_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_2_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_2_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_2_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_2_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_2_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_2_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_2_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_2_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_2_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_2_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_2_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_3_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_3_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_3_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_3_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_3_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_3_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_3_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_3_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_3_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_3_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_3_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_3_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_3_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_3_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_3_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_3_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_3_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_3_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_3_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_4_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_4_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_4_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_4_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_4_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_4_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_4_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_4_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_4_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_4_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_4_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_4_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_4_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_4_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_4_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_4_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_4_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_4_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_4_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_5_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_5_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_5_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_5_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_5_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_5_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_5_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_5_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_5_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_5_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_5_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_5_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_5_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_5_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_5_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_5_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_5_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_5_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_5_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_6_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_6_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_6_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_6_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_6_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_6_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_6_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_6_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_6_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_6_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_6_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_6_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_6_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_6_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_6_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_6_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_6_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_6_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_6_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_7_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_7_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_7_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_7_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_7_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_7_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_7_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_7_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_7_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_7_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_7_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_7_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_7_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_7_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_7_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_7_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_7_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_7_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_7_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_8_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_8_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_8_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_8_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_8_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_8_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_8_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_8_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_8_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_8_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_8_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_8_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_8_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_8_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_8_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_8_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_8_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_8_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_8_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_9_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_9_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_9_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_9_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_9_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_9_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_9_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_9_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_9_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_9_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_9_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_9_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_9_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_9_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_9_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_9_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_9_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_9_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_9_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_10_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_10_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_10_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_10_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_10_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_10_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_10_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_10_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_10_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_10_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_10_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_10_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_10_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_10_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_10_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_10_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_10_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_10_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_10_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_11_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_11_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_11_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_11_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_11_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_11_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_11_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_11_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_11_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_11_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_11_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_11_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_11_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_11_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_11_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_11_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_11_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_11_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_11_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_12_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_12_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_12_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_12_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_12_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_12_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_12_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_12_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_12_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_12_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_12_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_12_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_12_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_12_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_12_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_12_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_12_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_12_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_12_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_13_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_13_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_13_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_13_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_13_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_13_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_13_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_13_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_13_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_13_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_13_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_13_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_13_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_13_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_13_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_13_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_13_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_13_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_13_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_14_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_14_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_14_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_14_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_14_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_14_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_14_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_14_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_14_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_14_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_14_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_14_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_14_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_14_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_14_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_14_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_14_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_14_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_14_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_15_ARLEN = 8'h00;
	assign sync_argumentNotifierAXI_15_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_15_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_15_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_15_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_15_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_15_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_15_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_15_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_15_AWSIZE = 3'h2;
	assign sync_argumentNotifierAXI_15_AWBURST = 2'h1;
	assign sync_argumentNotifierAXI_15_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_15_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_15_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_15_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_15_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_15_WSTRB = 4'hf;
	assign sync_argumentNotifierAXI_15_WLAST = 1'h1;
	assign sync_argumentNotifierAXI_15_BREADY = 1'h1;
	assign sync_argumentNotifierAXI_16_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_16_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_16_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_16_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_16_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_16_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_16_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_16_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_16_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_16_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_16_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_16_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_16_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_16_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_16_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_16_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_16_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_16_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_16_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_16_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_16_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_16_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_16_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_17_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_17_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_17_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_17_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_17_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_17_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_17_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_17_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_17_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_17_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_17_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_17_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_17_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_17_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_17_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_17_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_17_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_17_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_17_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_17_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_17_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_17_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_17_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_18_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_18_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_18_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_18_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_18_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_18_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_18_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_18_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_18_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_18_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_18_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_18_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_18_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_18_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_18_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_18_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_18_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_18_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_18_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_18_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_18_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_18_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_18_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_19_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_19_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_19_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_19_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_19_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_19_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_19_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_19_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_19_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_19_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_19_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_19_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_19_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_19_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_19_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_19_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_19_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_19_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_19_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_19_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_19_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_19_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_19_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_20_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_20_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_20_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_20_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_20_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_20_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_20_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_20_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_20_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_20_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_20_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_20_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_20_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_20_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_20_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_20_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_20_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_20_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_20_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_20_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_20_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_20_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_20_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_21_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_21_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_21_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_21_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_21_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_21_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_21_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_21_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_21_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_21_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_21_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_21_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_21_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_21_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_21_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_21_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_21_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_21_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_21_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_21_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_21_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_21_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_21_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_22_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_22_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_22_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_22_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_22_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_22_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_22_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_22_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_22_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_22_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_22_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_22_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_22_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_22_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_22_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_22_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_22_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_22_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_22_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_22_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_22_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_22_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_22_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_23_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_23_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_23_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_23_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_23_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_23_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_23_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_23_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_23_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_23_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_23_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_23_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_23_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_23_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_23_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_23_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_23_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_23_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_23_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_23_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_23_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_23_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_23_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_24_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_24_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_24_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_24_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_24_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_24_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_24_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_24_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_24_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_24_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_24_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_24_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_24_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_24_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_24_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_24_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_24_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_24_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_24_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_24_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_24_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_24_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_24_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_25_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_25_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_25_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_25_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_25_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_25_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_25_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_25_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_25_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_25_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_25_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_25_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_25_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_25_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_25_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_25_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_25_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_25_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_25_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_25_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_25_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_25_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_25_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_26_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_26_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_26_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_26_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_26_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_26_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_26_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_26_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_26_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_26_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_26_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_26_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_26_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_26_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_26_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_26_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_26_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_26_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_26_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_26_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_26_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_26_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_26_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_27_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_27_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_27_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_27_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_27_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_27_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_27_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_27_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_27_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_27_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_27_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_27_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_27_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_27_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_27_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_27_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_27_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_27_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_27_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_27_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_27_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_27_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_27_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_28_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_28_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_28_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_28_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_28_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_28_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_28_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_28_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_28_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_28_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_28_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_28_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_28_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_28_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_28_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_28_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_28_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_28_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_28_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_28_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_28_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_28_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_28_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_29_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_29_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_29_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_29_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_29_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_29_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_29_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_29_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_29_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_29_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_29_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_29_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_29_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_29_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_29_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_29_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_29_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_29_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_29_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_29_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_29_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_29_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_29_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_30_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_30_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_30_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_30_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_30_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_30_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_30_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_30_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_30_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_30_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_30_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_30_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_30_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_30_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_30_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_30_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_30_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_30_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_30_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_30_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_30_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_30_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_30_BREADY = 1'h0;
	assign sync_argumentNotifierAXI_31_ARLEN = 8'h02;
	assign sync_argumentNotifierAXI_31_ARSIZE = 3'h2;
	assign sync_argumentNotifierAXI_31_ARBURST = 2'h1;
	assign sync_argumentNotifierAXI_31_ARLOCK = 1'h0;
	assign sync_argumentNotifierAXI_31_ARCACHE = 4'h0;
	assign sync_argumentNotifierAXI_31_ARPROT = 3'h0;
	assign sync_argumentNotifierAXI_31_ARQOS = 4'h0;
	assign sync_argumentNotifierAXI_31_ARREGION = 4'h0;
	assign sync_argumentNotifierAXI_31_AWVALID = 1'h0;
	assign sync_argumentNotifierAXI_31_AWADDR = 64'h0000000000000000;
	assign sync_argumentNotifierAXI_31_AWLEN = 8'h00;
	assign sync_argumentNotifierAXI_31_AWSIZE = 3'h0;
	assign sync_argumentNotifierAXI_31_AWBURST = 2'h0;
	assign sync_argumentNotifierAXI_31_AWLOCK = 1'h0;
	assign sync_argumentNotifierAXI_31_AWCACHE = 4'h0;
	assign sync_argumentNotifierAXI_31_AWPROT = 3'h0;
	assign sync_argumentNotifierAXI_31_AWQOS = 4'h0;
	assign sync_argumentNotifierAXI_31_AWREGION = 4'h0;
	assign sync_argumentNotifierAXI_31_WVALID = 1'h0;
	assign sync_argumentNotifierAXI_31_WDATA = 32'h00000000;
	assign sync_argumentNotifierAXI_31_WSTRB = 4'h0;
	assign sync_argumentNotifierAXI_31_WLAST = 1'h0;
	assign sync_argumentNotifierAXI_31_BREADY = 1'h0;
endmodule
